// Gate Level Verilog Code Generated!
// GateLvl:200 GateNum:200 GateInputNum:2
// ****** Basic Gate Module Defination ******
module or2(out, in1, in2);
  output out;
  input in1, in2;
  wire in1, in2, out;
  assign out = in1 || in2;
endmodule

module and2(out, in1, in2);
  output out;
  input in1, in2;
  wire in1, in2, out;
  assign out = in1 && in2;
endmodule

module not1(out, in);
  output out;
  input in;
  wire in,out;
  assign out = ~in;
endmodule

module nand2(out, in1, in2);
  output out;
  input in1, in2;
  wire in1, in2, out;
  assign out = ~(in1 && in2);
endmodule
// ****** Basic Gate Module Defination End ******

// ****** Combined Logic Module Defination ******
module combLogic( w_000_000, w_000_001, w_000_002, w_000_003, w_000_004, w_000_005, w_000_006, w_000_007, w_000_008, w_000_009, w_000_010, w_000_011, w_000_012, w_000_013, w_000_014, w_000_015, w_000_016, w_000_017, w_000_018, w_000_019, w_000_020, w_000_021, w_000_022, w_000_023, w_000_024, w_000_025, w_000_026, w_000_027, w_000_028, w_000_029, w_000_030, w_000_031, w_000_032, w_000_033, w_000_034, w_000_035, w_000_036, w_000_037, w_000_038, w_000_039, w_000_040, w_000_041, w_000_042, w_000_043, w_000_044, w_000_045, w_000_046, w_000_047, w_000_048, w_000_049, w_000_050, w_000_051, w_000_052, w_000_053, w_000_054, w_000_055, w_000_056, w_000_057, w_000_058, w_000_059, w_000_060, w_000_061, w_000_062, w_000_063, w_000_064, w_000_065, w_000_066, w_000_067, w_000_068, w_000_069, w_000_070, w_000_071, w_000_072, w_000_073, w_000_074, w_000_075, w_000_076, w_000_077, w_000_078, w_000_079, w_000_080, w_000_081, w_000_082, w_000_083, w_000_084, w_000_085, w_000_086, w_000_087, w_000_088, w_000_089, w_000_090, w_000_091, w_000_092, w_000_093, w_000_094, w_000_095, w_000_096, w_000_097, w_000_098, w_000_099, w_000_100, w_000_102, w_000_103, w_000_104, w_000_105, w_000_106, w_000_109, w_000_110, w_000_111, w_000_112, w_000_113, w_000_114, w_000_115, w_000_116, w_000_117, w_000_119, w_000_120, w_000_121, w_000_122, w_000_124, w_000_125, w_000_126, w_000_127, w_000_128, w_000_129, w_000_130, w_000_131, w_000_132, w_000_135, w_000_136, w_000_137, w_000_138, w_000_139, w_000_140, w_000_142, w_000_143, w_000_144, w_000_145, w_000_148, w_000_150, w_000_151, w_000_152, w_000_153, w_000_154, w_000_155, w_000_157, w_000_159, w_000_160, w_000_161, w_000_162, w_000_165, w_000_166, w_000_168, w_000_169, w_000_170, w_000_172, w_000_173, w_000_175, w_000_177, w_000_178, w_000_180, w_000_186, w_000_189, w_200_000, w_200_001, w_200_002, w_200_003, w_200_004, w_200_005, w_200_006, w_200_007, w_200_008, w_200_009, w_200_010, w_200_011, w_200_012, w_200_013, w_200_014, w_200_015, w_200_016, w_200_017, w_200_018, w_200_019, w_200_020, w_200_021, w_200_022, w_200_023, w_200_024, w_200_025, w_200_026, w_200_027, w_200_028, w_200_029, w_200_030, w_200_031, w_200_032, w_200_033, w_200_034, w_200_035, w_200_036, w_200_037, w_200_038, w_200_039, w_200_040, w_200_041, w_200_042, w_200_043, w_200_044, w_200_045, w_200_046, w_200_047, w_200_048, w_200_049, w_200_050, w_200_051, w_200_052, w_200_053, w_200_054, w_200_055, w_200_056, w_200_057, w_200_058, w_200_059, w_200_060, w_200_061, w_200_062, w_200_063, w_200_064, w_200_065, w_200_066, w_200_067, w_200_068, w_200_069, w_200_070, w_200_071, w_200_072, w_200_073, w_200_074, w_200_075, w_200_076, w_200_077, w_200_078, w_200_079, w_200_080, w_200_081, w_200_082, w_200_083, w_200_084, w_200_085, w_200_086, w_200_087 );
  inout w_000_000, w_000_001, w_000_002, w_000_003, w_000_004, w_000_005, w_000_006, w_000_007, w_000_008, w_000_009, w_000_010, w_000_011, w_000_012, w_000_013, w_000_014, w_000_015, w_000_016, w_000_017, w_000_018, w_000_019, w_000_020, w_000_021, w_000_022, w_000_023, w_000_024, w_000_025, w_000_026, w_000_027, w_000_028, w_000_029, w_000_030, w_000_031, w_000_032, w_000_033, w_000_034, w_000_035, w_000_036, w_000_037, w_000_038, w_000_039, w_000_040, w_000_041, w_000_042, w_000_043, w_000_044, w_000_045, w_000_046, w_000_047, w_000_048, w_000_049, w_000_050, w_000_051, w_000_052, w_000_053, w_000_054, w_000_055, w_000_056, w_000_057, w_000_058, w_000_059, w_000_060, w_000_061, w_000_062, w_000_063, w_000_064, w_000_065, w_000_066, w_000_067, w_000_068, w_000_069, w_000_070, w_000_071, w_000_072, w_000_073, w_000_074, w_000_075, w_000_076, w_000_077, w_000_078, w_000_079, w_000_080, w_000_081, w_000_082, w_000_083, w_000_084, w_000_085, w_000_086, w_000_087, w_000_088, w_000_089, w_000_090, w_000_091, w_000_092, w_000_093, w_000_094, w_000_095, w_000_096, w_000_097, w_000_098, w_000_099, w_000_100, w_000_102, w_000_103, w_000_104, w_000_105, w_000_106, w_000_109, w_000_110, w_000_111, w_000_112, w_000_113, w_000_114, w_000_115, w_000_116, w_000_117, w_000_119, w_000_120, w_000_121, w_000_122, w_000_124, w_000_125, w_000_126, w_000_127, w_000_128, w_000_129, w_000_130, w_000_131, w_000_132, w_000_135, w_000_136, w_000_137, w_000_138, w_000_139, w_000_140, w_000_142, w_000_143, w_000_144, w_000_145, w_000_148, w_000_150, w_000_151, w_000_152, w_000_153, w_000_154, w_000_155, w_000_157, w_000_159, w_000_160, w_000_161, w_000_162, w_000_165, w_000_166, w_000_168, w_000_169, w_000_170, w_000_172, w_000_173, w_000_175, w_000_177, w_000_178, w_000_180, w_000_186, w_000_189;
  output w_200_000, w_200_001, w_200_002, w_200_003, w_200_004, w_200_005, w_200_006, w_200_007, w_200_008, w_200_009, w_200_010, w_200_011, w_200_012, w_200_013, w_200_014, w_200_015, w_200_016, w_200_017, w_200_018, w_200_019, w_200_020, w_200_021, w_200_022, w_200_023, w_200_024, w_200_025, w_200_026, w_200_027, w_200_028, w_200_029, w_200_030, w_200_031, w_200_032, w_200_033, w_200_034, w_200_035, w_200_036, w_200_037, w_200_038, w_200_039, w_200_040, w_200_041, w_200_042, w_200_043, w_200_044, w_200_045, w_200_046, w_200_047, w_200_048, w_200_049, w_200_050, w_200_051, w_200_052, w_200_053, w_200_054, w_200_055, w_200_056, w_200_057, w_200_058, w_200_059, w_200_060, w_200_061, w_200_062, w_200_063, w_200_064, w_200_065, w_200_066, w_200_067, w_200_068, w_200_069, w_200_070, w_200_071, w_200_072, w_200_073, w_200_074, w_200_075, w_200_076, w_200_077, w_200_078, w_200_079, w_200_080, w_200_081, w_200_082, w_200_083, w_200_084, w_200_085, w_200_086, w_200_087;
  wire w_000_000, w_000_001, w_000_002, w_000_003, w_000_004, w_000_005, w_000_006, w_000_007, w_000_008, w_000_009, w_000_010, w_000_011, w_000_012, w_000_013, w_000_014, w_000_015, w_000_016, w_000_017, w_000_018, w_000_019, w_000_020, w_000_021, w_000_022, w_000_023, w_000_024, w_000_025, w_000_026, w_000_027, w_000_028, w_000_029, w_000_030, w_000_031, w_000_032, w_000_033, w_000_034, w_000_035, w_000_036, w_000_037, w_000_038, w_000_039, w_000_040, w_000_041, w_000_042, w_000_043, w_000_044, w_000_045, w_000_046, w_000_047, w_000_048, w_000_049, w_000_050, w_000_051, w_000_052, w_000_053, w_000_054, w_000_055, w_000_056, w_000_057, w_000_058, w_000_059, w_000_060, w_000_061, w_000_062, w_000_063, w_000_064, w_000_065, w_000_066, w_000_067, w_000_068, w_000_069, w_000_070, w_000_071, w_000_072, w_000_073, w_000_074, w_000_075, w_000_076, w_000_077, w_000_078, w_000_079, w_000_080, w_000_081, w_000_082, w_000_083, w_000_084, w_000_085, w_000_086, w_000_087, w_000_088, w_000_089, w_000_090, w_000_091, w_000_092, w_000_093, w_000_094, w_000_095, w_000_096, w_000_097, w_000_098, w_000_099, w_000_100, w_000_102, w_000_103, w_000_104, w_000_105, w_000_106, w_000_109, w_000_110, w_000_111, w_000_112, w_000_113, w_000_114, w_000_115, w_000_116, w_000_117, w_000_119, w_000_120, w_000_121, w_000_122, w_000_124, w_000_125, w_000_126, w_000_127, w_000_128, w_000_129, w_000_130, w_000_131, w_000_132, w_000_135, w_000_136, w_000_137, w_000_138, w_000_139, w_000_140, w_000_142, w_000_143, w_000_144, w_000_145, w_000_148, w_000_150, w_000_151, w_000_152, w_000_153, w_000_154, w_000_155, w_000_157, w_000_159, w_000_160, w_000_161, w_000_162, w_000_165, w_000_166, w_000_168, w_000_169, w_000_170, w_000_172, w_000_173, w_000_175, w_000_177, w_000_178, w_000_180, w_000_186, w_000_189;
  wire w_001_000, w_001_001, w_001_002, w_001_003, w_001_004, w_001_005, w_001_006, w_001_007, w_001_008, w_001_009, w_001_010, w_001_011, w_001_012, w_001_013, w_001_014, w_001_015, w_001_016, w_001_017, w_001_018;
  wire w_002_000, w_002_001, w_002_002, w_002_003, w_002_004, w_002_005, w_002_006, w_002_007, w_002_008, w_002_009, w_002_010, w_002_011, w_002_012, w_002_014, w_002_015, w_002_016, w_002_017, w_002_018, w_002_019, w_002_020, w_002_021, w_002_022, w_002_023, w_002_024, w_002_025, w_002_026, w_002_027, w_002_028, w_002_029, w_002_030, w_002_031, w_002_032, w_002_033, w_002_034, w_002_035, w_002_036, w_002_037, w_002_038, w_002_039, w_002_040, w_002_041, w_002_042, w_002_043, w_002_044, w_002_045, w_002_046, w_002_047, w_002_048, w_002_049, w_002_050, w_002_051, w_002_052, w_002_053, w_002_054, w_002_055, w_002_056, w_002_057, w_002_058, w_002_059, w_002_060, w_002_061, w_002_062, w_002_063, w_002_064;
  wire w_003_000, w_003_001, w_003_002, w_003_003, w_003_004, w_003_005, w_003_006, w_003_007, w_003_008, w_003_009, w_003_010, w_003_011, w_003_012, w_003_013, w_003_014, w_003_015, w_003_016, w_003_017, w_003_018, w_003_019, w_003_020, w_003_021, w_003_022, w_003_023, w_003_024, w_003_025, w_003_026, w_003_027, w_003_028, w_003_029, w_003_030, w_003_031, w_003_032;
  wire w_004_000, w_004_001, w_004_003, w_004_004, w_004_005, w_004_006, w_004_007, w_004_009, w_004_010, w_004_011, w_004_012, w_004_014, w_004_015, w_004_016, w_004_017, w_004_018, w_004_021, w_004_022, w_004_023, w_004_024, w_004_025, w_004_026, w_004_028, w_004_030, w_004_031, w_004_032, w_004_033, w_004_034, w_004_035, w_004_036, w_004_037, w_004_038, w_004_039, w_004_040, w_004_042, w_004_043, w_004_044, w_004_045, w_004_046, w_004_047, w_004_048, w_004_049, w_004_050, w_004_051, w_004_052, w_004_053, w_004_057, w_004_058, w_004_059, w_004_061, w_004_062, w_004_063, w_004_064, w_004_065, w_004_067, w_004_069, w_004_071, w_004_072, w_004_073, w_004_074, w_004_076, w_004_077, w_004_079, w_004_080, w_004_082, w_004_085, w_004_088, w_004_090, w_004_092, w_004_094, w_004_096, w_004_098, w_004_104, w_004_105, w_004_107, w_004_110, w_004_111, w_004_112, w_004_115;
  wire w_005_000, w_005_001, w_005_003, w_005_004, w_005_005, w_005_007, w_005_008, w_005_009, w_005_010, w_005_011, w_005_012, w_005_013, w_005_014, w_005_015, w_005_016, w_005_017, w_005_018, w_005_019, w_005_020, w_005_022, w_005_023, w_005_024, w_005_025, w_005_026, w_005_027, w_005_028, w_005_029, w_005_030, w_005_031, w_005_032, w_005_033, w_005_035, w_005_036, w_005_037, w_005_038, w_005_039, w_005_040, w_005_041, w_005_042, w_005_044, w_005_045, w_005_047, w_005_048, w_005_050, w_005_051, w_005_052, w_005_053, w_005_054, w_005_055, w_005_056, w_005_058, w_005_060, w_005_061, w_005_062, w_005_063, w_005_064, w_005_065, w_005_066, w_005_068, w_005_069, w_005_070, w_005_071;
  wire w_006_000, w_006_001, w_006_002, w_006_003, w_006_004, w_006_005, w_006_006, w_006_008, w_006_009, w_006_012, w_006_013, w_006_015, w_006_016, w_006_017, w_006_018, w_006_020, w_006_021, w_006_022, w_006_023, w_006_024, w_006_027, w_006_028, w_006_029, w_006_031, w_006_032, w_006_033, w_006_034, w_006_035, w_006_038, w_006_043, w_006_044, w_006_045, w_006_047, w_006_048, w_006_049, w_006_050, w_006_051, w_006_053, w_006_054, w_006_055, w_006_056, w_006_058, w_006_059, w_006_060, w_006_061, w_006_062, w_006_065, w_006_066, w_006_068, w_006_069, w_006_070, w_006_072, w_006_074, w_006_075, w_006_078, w_006_080, w_006_081, w_006_083, w_006_084, w_006_086, w_006_090, w_006_092, w_006_093, w_006_094, w_006_096, w_006_097, w_006_099, w_006_100, w_006_101, w_006_103, w_006_104, w_006_106, w_006_107, w_006_109, w_006_112, w_006_117, w_006_118, w_006_119, w_006_120, w_006_121, w_006_123;
  wire w_007_000, w_007_001, w_007_002, w_007_003, w_007_004, w_007_005, w_007_006, w_007_008, w_007_009, w_007_010, w_007_012, w_007_013, w_007_014, w_007_015, w_007_016, w_007_017, w_007_019, w_007_020, w_007_021, w_007_022, w_007_023, w_007_024, w_007_025, w_007_027, w_007_029, w_007_031, w_007_032, w_007_033, w_007_034, w_007_036, w_007_037, w_007_038, w_007_039, w_007_040, w_007_041, w_007_042, w_007_043, w_007_044, w_007_046, w_007_047, w_007_048, w_007_049, w_007_050, w_007_051, w_007_052, w_007_053, w_007_054;
  wire w_008_000, w_008_001, w_008_002, w_008_003, w_008_004, w_008_005, w_008_006, w_008_008, w_008_009, w_008_010, w_008_012, w_008_013, w_008_014, w_008_015, w_008_018, w_008_020, w_008_021, w_008_025, w_008_026, w_008_028, w_008_031, w_008_033, w_008_036, w_008_038, w_008_039, w_008_040, w_008_044, w_008_047, w_008_048, w_008_049, w_008_050, w_008_051, w_008_052, w_008_054, w_008_055, w_008_056, w_008_057, w_008_059, w_008_062, w_008_063, w_008_064, w_008_065, w_008_066, w_008_069, w_008_071, w_008_075, w_008_076, w_008_078, w_008_080, w_008_081, w_008_084, w_008_086, w_008_088, w_008_090, w_008_091, w_008_093, w_008_099, w_008_100, w_008_104, w_008_105, w_008_108, w_008_109, w_008_110, w_008_112, w_008_115, w_008_120;
  wire w_009_004, w_009_005, w_009_006, w_009_010, w_009_012, w_009_015, w_009_018, w_009_023, w_009_026, w_009_027, w_009_028, w_009_030, w_009_031, w_009_033, w_009_034, w_009_035, w_009_037, w_009_038, w_009_040, w_009_041, w_009_042, w_009_043, w_009_044, w_009_046, w_009_047, w_009_052, w_009_054, w_009_055, w_009_057, w_009_060, w_009_062, w_009_063, w_009_064, w_009_071, w_009_077, w_009_078, w_009_080, w_009_081, w_009_082, w_009_083, w_009_086, w_009_089, w_009_091, w_009_092, w_009_095, w_009_097, w_009_105, w_009_107, w_009_114, w_009_117, w_009_118, w_009_122, w_009_123, w_009_125, w_009_127, w_009_134, w_009_135, w_009_138, w_009_139;
  wire w_010_000, w_010_002, w_010_003, w_010_004, w_010_005, w_010_006, w_010_007, w_010_008, w_010_009, w_010_010, w_010_011, w_010_012, w_010_014, w_010_015, w_010_016, w_010_017, w_010_019, w_010_022, w_010_023, w_010_025, w_010_026, w_010_027, w_010_028, w_010_029, w_010_030, w_010_032, w_010_033, w_010_034, w_010_035, w_010_037, w_010_038, w_010_040, w_010_042, w_010_043, w_010_044, w_010_046, w_010_047, w_010_048, w_010_049;
  wire w_011_000, w_011_002, w_011_008, w_011_015, w_011_016, w_011_020, w_011_023, w_011_024, w_011_026, w_011_029, w_011_031, w_011_032, w_011_033, w_011_034, w_011_040, w_011_042, w_011_043, w_011_047, w_011_050, w_011_051, w_011_052, w_011_053, w_011_054, w_011_055, w_011_057, w_011_060, w_011_071, w_011_072, w_011_073, w_011_074, w_011_077, w_011_079, w_011_080, w_011_082, w_011_085, w_011_091, w_011_092, w_011_093, w_011_095, w_011_101, w_011_106, w_011_108, w_011_113, w_011_115, w_011_116, w_011_117, w_011_119, w_011_122, w_011_124, w_011_125, w_011_128, w_011_132, w_011_133, w_011_134, w_011_136, w_011_137, w_011_140;
  wire w_012_000, w_012_001, w_012_003, w_012_009, w_012_010, w_012_011, w_012_012, w_012_013, w_012_015, w_012_016, w_012_018, w_012_025, w_012_027, w_012_029, w_012_030, w_012_031, w_012_032, w_012_033, w_012_035, w_012_039, w_012_043, w_012_045, w_012_048, w_012_049, w_012_054, w_012_056, w_012_057, w_012_067, w_012_072, w_012_075, w_012_078, w_012_080, w_012_082, w_012_084, w_012_086, w_012_087, w_012_090, w_012_095, w_012_103, w_012_107, w_012_110, w_012_116, w_012_119, w_012_127, w_012_128;
  wire w_013_000, w_013_001, w_013_002, w_013_003, w_013_008, w_013_009, w_013_010, w_013_012, w_013_016, w_013_017, w_013_018, w_013_020, w_013_021, w_013_022, w_013_023, w_013_024, w_013_026, w_013_027, w_013_030, w_013_031, w_013_032, w_013_036, w_013_037, w_013_038, w_013_042, w_013_044, w_013_045, w_013_046, w_013_047, w_013_048, w_013_049, w_013_050, w_013_057, w_013_059, w_013_060, w_013_061, w_013_063, w_013_064, w_013_067, w_013_071;
  wire w_014_004, w_014_005, w_014_007, w_014_009, w_014_015, w_014_020, w_014_021, w_014_030, w_014_031, w_014_035, w_014_037, w_014_038, w_014_040, w_014_042, w_014_046, w_014_047, w_014_052, w_014_053, w_014_055, w_014_056, w_014_057, w_014_058, w_014_059, w_014_064, w_014_065, w_014_066, w_014_070, w_014_072, w_014_074, w_014_077, w_014_078, w_014_080, w_014_081, w_014_093, w_014_100, w_014_102, w_014_118, w_014_121, w_014_122, w_014_125, w_014_130, w_014_139;
  wire w_015_002, w_015_003, w_015_005, w_015_012, w_015_015, w_015_021, w_015_022, w_015_024, w_015_025, w_015_027, w_015_029, w_015_033, w_015_034, w_015_036, w_015_037, w_015_043, w_015_044, w_015_047, w_015_050, w_015_053, w_015_054, w_015_056, w_015_057, w_015_058, w_015_059, w_015_062, w_015_064, w_015_065, w_015_066, w_015_076, w_015_084, w_015_085, w_015_086, w_015_092, w_015_106, w_015_113, w_015_115, w_015_118, w_015_120, w_015_123, w_015_126;
  wire w_016_005, w_016_007, w_016_008, w_016_009, w_016_012, w_016_015, w_016_016, w_016_017, w_016_021, w_016_022, w_016_023, w_016_025, w_016_027, w_016_029, w_016_030, w_016_031, w_016_036, w_016_039, w_016_043, w_016_045, w_016_046, w_016_049, w_016_050, w_016_051, w_016_056, w_016_065, w_016_066, w_016_067, w_016_070, w_016_071, w_016_073, w_016_074, w_016_075, w_016_076, w_016_079;
  wire w_017_002, w_017_004, w_017_006, w_017_010, w_017_011, w_017_022, w_017_026, w_017_027, w_017_030, w_017_031, w_017_032, w_017_033, w_017_038, w_017_041, w_017_042, w_017_045, w_017_047, w_017_056, w_017_059, w_017_061, w_017_065, w_017_070, w_017_076, w_017_080, w_017_090, w_017_097, w_017_100, w_017_104, w_017_107, w_017_108, w_017_113, w_017_134;
  wire w_018_000, w_018_012, w_018_017, w_018_020, w_018_023, w_018_028, w_018_032, w_018_033, w_018_035, w_018_037, w_018_046, w_018_051, w_018_052, w_018_058, w_018_059, w_018_061, w_018_062, w_018_064, w_018_072, w_018_073, w_018_081, w_018_082, w_018_083, w_018_089, w_018_110, w_018_118, w_018_122;
  wire w_019_003, w_019_017, w_019_020, w_019_021, w_019_028, w_019_033, w_019_036, w_019_043, w_019_051, w_019_052, w_019_053, w_019_057, w_019_071, w_019_074, w_019_078, w_019_087, w_019_091, w_019_103, w_019_105, w_019_106, w_019_111, w_019_113, w_019_121, w_019_124, w_019_125, w_019_126, w_019_135, w_019_136;
  wire w_020_000, w_020_003, w_020_004, w_020_005, w_020_007, w_020_008, w_020_009, w_020_010, w_020_011, w_020_014, w_020_015;
  wire w_021_001, w_021_003, w_021_007, w_021_008, w_021_011, w_021_013, w_021_015, w_021_023, w_021_024, w_021_032, w_021_036, w_021_043, w_021_044, w_021_048, w_021_051, w_021_054, w_021_055, w_021_080, w_021_097, w_021_108, w_021_112, w_021_113, w_021_114, w_021_121, w_021_139, w_021_156, w_021_157, w_021_158, w_021_159, w_021_160, w_021_161, w_021_162, w_021_166, w_021_167, w_021_168, w_021_169, w_021_170, w_021_171, w_021_172, w_021_173, w_021_174, w_021_176, w_021_178, w_021_179, w_021_180, w_021_181, w_021_182, w_021_183;
  wire w_022_000, w_022_008, w_022_009, w_022_015, w_022_018, w_022_019, w_022_022, w_022_026, w_022_027, w_022_030, w_022_033, w_022_034, w_022_045, w_022_054, w_022_055, w_022_071, w_022_075, w_022_078, w_022_079, w_022_088, w_022_094, w_022_101;
  wire w_023_013, w_023_015, w_023_018, w_023_028, w_023_030, w_023_033, w_023_036, w_023_038, w_023_039, w_023_041, w_023_044, w_023_048, w_023_053, w_023_056, w_023_060, w_023_061, w_023_067, w_023_087, w_023_091, w_023_098, w_023_116, w_023_118;
  wire w_024_000, w_024_001, w_024_002, w_024_003, w_024_005, w_024_006, w_024_008, w_024_009, w_024_010;
  wire w_025_004, w_025_009, w_025_027, w_025_028, w_025_033, w_025_036, w_025_050, w_025_065, w_025_068, w_025_072, w_025_082, w_025_087, w_025_093, w_025_096, w_025_106, w_025_109, w_025_111, w_025_123, w_025_128, w_025_132;
  wire w_026_001, w_026_004, w_026_005, w_026_006, w_026_012, w_026_015, w_026_017, w_026_029, w_026_035, w_026_040, w_026_042, w_026_053, w_026_054, w_026_069, w_026_070, w_026_074, w_026_077, w_026_085, w_026_087, w_026_088, w_026_092, w_026_093, w_026_094, w_026_095;
  wire w_027_005, w_027_006, w_027_014, w_027_020, w_027_030, w_027_031, w_027_032, w_027_037, w_027_043, w_027_048, w_027_050, w_027_051, w_027_054, w_027_055, w_027_058, w_027_060, w_027_062, w_027_063;
  wire w_028_000, w_028_001, w_028_007, w_028_009, w_028_010, w_028_011, w_028_013, w_028_018, w_028_026, w_028_029, w_028_034, w_028_039, w_028_041, w_028_045, w_028_056, w_028_066, w_028_070, w_028_080, w_028_086, w_028_087, w_028_091, w_028_101, w_028_113, w_028_132, w_028_138, w_028_160, w_028_161, w_028_162, w_028_163, w_028_164, w_028_165, w_028_166, w_028_167, w_028_168, w_028_169, w_028_171, w_028_173, w_028_174, w_028_175, w_028_176, w_028_177;
  wire w_029_000, w_029_001, w_029_003, w_029_004, w_029_005, w_029_006, w_029_007, w_029_008, w_029_009, w_029_011, w_029_012, w_029_013, w_029_014, w_029_015, w_029_016, w_029_017, w_029_018, w_029_019, w_029_020;
  wire w_030_003, w_030_005, w_030_022, w_030_026, w_030_033, w_030_061, w_030_063;
  wire w_031_002, w_031_005, w_031_009, w_031_014, w_031_016, w_031_021, w_031_022, w_031_036, w_031_039, w_031_044, w_031_045, w_031_054, w_031_057, w_031_068, w_031_076, w_031_087, w_031_089, w_031_093, w_031_097, w_031_103, w_031_105, w_031_118, w_031_129, w_031_131, w_031_135;
  wire w_032_001, w_032_011, w_032_019, w_032_024, w_032_029, w_032_033, w_032_039, w_032_054, w_032_062, w_032_065, w_032_067, w_032_069, w_032_082, w_032_103, w_032_105, w_032_122;
  wire w_033_005, w_033_006, w_033_007, w_033_008, w_033_012, w_033_014, w_033_018, w_033_029, w_033_030, w_033_031, w_033_034, w_033_035, w_033_037, w_033_040, w_033_044, w_033_049;
  wire w_034_001, w_034_002, w_034_014, w_034_017, w_034_018, w_034_030, w_034_041, w_034_050, w_034_065, w_034_069, w_034_072, w_034_074, w_034_088, w_034_105, w_034_117, w_034_128, w_034_134, w_034_136;
  wire w_035_005, w_035_018, w_035_027, w_035_031, w_035_040, w_035_042, w_035_044, w_035_052, w_035_057, w_035_070, w_035_073, w_035_076, w_035_079, w_035_082, w_035_083;
  wire w_036_000, w_036_002, w_036_003, w_036_004, w_036_005, w_036_006, w_036_008, w_036_012;
  wire w_037_000, w_037_003, w_037_004, w_037_012, w_037_075, w_037_090, w_037_126, w_037_128, w_037_153;
  wire w_038_000, w_038_002, w_038_003, w_038_004, w_038_005, w_038_006, w_038_007, w_038_012, w_038_013, w_038_014, w_038_016, w_038_017, w_038_020, w_038_021, w_038_022, w_038_023, w_038_024;
  wire w_039_000, w_039_001, w_039_002, w_039_004, w_039_005, w_039_006, w_039_007, w_039_011, w_039_012, w_039_013, w_039_014, w_039_015, w_039_016, w_039_017, w_039_018, w_039_019, w_039_020, w_039_021, w_039_025, w_039_026, w_039_027, w_039_028, w_039_029, w_039_030, w_039_031, w_039_032, w_039_033, w_039_034, w_039_036;
  wire w_040_009, w_040_016, w_040_018, w_040_037, w_040_043, w_040_047, w_040_053, w_040_059, w_040_069, w_040_082, w_040_106, w_040_115;
  wire w_041_023, w_041_029, w_041_035, w_041_059, w_041_081, w_041_116;
  wire w_042_011, w_042_015, w_042_016, w_042_034, w_042_041, w_042_049, w_042_054;
  wire w_043_016, w_043_020, w_043_025, w_043_030, w_043_036, w_043_053, w_043_062;
  wire w_044_000, w_044_013, w_044_040, w_044_058, w_044_099, w_044_139, w_044_159, w_044_161, w_044_166, w_044_170, w_044_180;
  wire w_045_009, w_045_013, w_045_038, w_045_039, w_045_041, w_045_042, w_045_051;
  wire w_046_010, w_046_020, w_046_028, w_046_030, w_046_051, w_046_055, w_046_056, w_046_090, w_046_092, w_046_103, w_046_130;
  wire w_047_006, w_047_012, w_047_013, w_047_021, w_047_027, w_047_030, w_047_033, w_047_035, w_047_048;
  wire w_048_008, w_048_017, w_048_051, w_048_058, w_048_076, w_048_109, w_048_136, w_048_157;
  wire w_049_008, w_049_036, w_049_045, w_049_046, w_049_059, w_049_069, w_049_103, w_049_107, w_049_125, w_049_126, w_049_129;
  wire w_050_006, w_050_020, w_050_025, w_050_032, w_050_045, w_050_049, w_050_054, w_050_062, w_050_063, w_050_069, w_050_074, w_050_076, w_050_096, w_050_112, w_050_113;
  wire w_051_006, w_051_027, w_051_056, w_051_122, w_051_143;
  wire w_052_027, w_052_031, w_052_040, w_052_050, w_052_055;
  wire w_053_005, w_053_012, w_053_032, w_053_033, w_053_045, w_053_065;
  wire w_054_000, w_054_001, w_054_002, w_054_003, w_054_004, w_054_005, w_054_008, w_054_009;
  wire w_055_015, w_055_024, w_055_035, w_055_077, w_055_087, w_055_132, w_055_177;
  wire w_056_001, w_056_014, w_056_018, w_056_058, w_056_070, w_056_074, w_056_099, w_056_103, w_056_104;
  wire w_057_026, w_057_031, w_057_051, w_057_083;
  wire w_058_000, w_058_018, w_058_019, w_058_028, w_058_031, w_058_036, w_058_039, w_058_067, w_058_069, w_058_072, w_058_089;
  wire w_059_011, w_059_039, w_059_046, w_059_058, w_059_065, w_059_070, w_059_073, w_059_085, w_059_097, w_059_117, w_059_134, w_059_163;
  wire w_060_006, w_060_007, w_060_029, w_060_030, w_060_044, w_060_045, w_060_049, w_060_061;
  wire w_061_003, w_061_035, w_061_072, w_061_096;
  wire w_062_003, w_062_060, w_062_125, w_062_127, w_062_194;
  wire w_063_007, w_063_010, w_063_029, w_063_068, w_063_078;
  wire w_064_028, w_064_035, w_064_037, w_064_070, w_064_079, w_064_130, w_064_144, w_064_152, w_064_165;
  wire w_065_004, w_065_037, w_065_062, w_065_064;
  wire w_066_011, w_066_065, w_066_088, w_066_126, w_066_138, w_066_156;
  wire w_067_022, w_067_028, w_067_046, w_067_047;
  wire w_068_018, w_068_029, w_068_035, w_068_046;
  wire w_069_100, w_069_133, w_069_155;
  wire w_070_026, w_070_044, w_070_055, w_070_062, w_070_083, w_070_084, w_070_085, w_070_086, w_070_087, w_070_088, w_070_089, w_070_090, w_070_091, w_070_093;
  wire w_071_007, w_071_017, w_071_028, w_071_076;
  wire w_072_051, w_072_096, w_072_103, w_072_150;
  wire w_073_009, w_073_015, w_073_025, w_073_062;
  wire w_074_069, w_074_087, w_074_136, w_074_138;
  wire w_075_023, w_075_036;
  wire w_076_008, w_076_023, w_076_156, w_076_167;
  wire w_077_017, w_077_019, w_077_031, w_077_032;
  wire w_078_010, w_078_015, w_078_024, w_078_026, w_078_043, w_078_070;
  wire w_079_003, w_079_004, w_079_008, w_079_009;
  wire w_080_001, w_080_008, w_080_024, w_080_032, w_080_036;
  wire w_081_017, w_081_026, w_081_027, w_081_054, w_081_091;
  wire w_082_008, w_082_012, w_082_020, w_082_051, w_082_061, w_082_063;
  wire w_083_012, w_083_036, w_083_059, w_083_069;
  wire w_084_015, w_084_028, w_084_036, w_084_079;
  wire w_085_015, w_085_044;
  wire w_086_026, w_086_029, w_086_035;
  wire w_087_016, w_087_032;
  wire w_088_005, w_088_033;
  wire w_089_016, w_089_020, w_089_033, w_089_039;
  wire w_090_015, w_090_020, w_090_029, w_090_069;
  wire w_091_011, w_091_100, w_091_148;
  wire w_092_038, w_092_053, w_092_109, w_092_121;
  wire w_093_030, w_093_042;
  wire w_094_075, w_094_080, w_094_084, w_094_086;
  wire w_096_009, w_096_015, w_096_016, w_096_023;
  wire w_097_003, w_097_018, w_097_020, w_097_054, w_097_055, w_097_056;
  wire w_098_036, w_098_077, w_098_079;
  wire w_099_029;
  wire w_100_002, w_100_018, w_100_019, w_100_020;
  wire w_101_001, w_101_005, w_101_025;
  wire w_102_079, w_102_104, w_102_135;
  wire w_103_013, w_103_094, w_103_127, w_103_138;
  wire w_104_104, w_104_119;
  wire w_105_182;
  wire w_106_000, w_106_008;
  wire w_107_013, w_107_019, w_107_063, w_107_152;
  wire w_108_023, w_108_027;
  wire w_109_069, w_109_075, w_109_106, w_109_122;
  wire w_110_022;
  wire w_111_008, w_111_011, w_111_039;
  wire w_112_061, w_112_075, w_112_089;
  wire w_113_001;
  wire w_114_053, w_114_100, w_114_101, w_114_102, w_114_103, w_114_107, w_114_108, w_114_109, w_114_110, w_114_111, w_114_112, w_114_113, w_114_114, w_114_115;
  wire w_115_011;
  wire w_117_000, w_117_001;
  wire w_118_025, w_118_030, w_118_066;
  wire w_119_006, w_119_011;
  wire w_120_011, w_120_172;
  wire w_121_013;
  wire w_122_028, w_122_059;
  wire w_123_000, w_123_044, w_123_108;
  wire w_124_047;
  wire w_126_001, w_126_002;
  wire w_127_005;
  wire w_128_022;
  wire w_129_002, w_129_036;
  wire w_130_051, w_130_117, w_130_176;
  wire w_131_037, w_131_101;
  wire w_132_041, w_132_053, w_132_054, w_132_055, w_132_056, w_132_057, w_132_058, w_132_059, w_132_060, w_132_061, w_132_062, w_132_063, w_132_065;
  wire w_133_007, w_133_012, w_133_038, w_133_143, w_133_153, w_133_154, w_133_155, w_133_156, w_133_157, w_133_158, w_133_159, w_133_160, w_133_161, w_133_162, w_133_163, w_133_164;
  wire w_134_007, w_134_020;
  wire w_135_079;
  wire w_136_034;
  wire w_137_005;
  wire w_138_132, w_138_148;
  wire w_139_031;
  wire w_140_044;
  wire w_141_004;
  wire w_142_002, w_142_006;
  wire w_143_001;
  wire w_144_036, w_144_052, w_144_096, w_144_198, w_144_199, w_144_200, w_144_201, w_144_202, w_144_203, w_144_204, w_144_208, w_144_209, w_144_210, w_144_211, w_144_213;
  wire w_145_004, w_145_013;
  wire w_146_018, w_146_126;
  wire w_147_016, w_147_061, w_147_080;
  wire w_149_015, w_149_019;
  wire w_150_008, w_150_009, w_150_010, w_150_011, w_150_012, w_150_013, w_150_014, w_150_015, w_150_016;
  wire w_151_148;
  wire w_152_057;
  wire w_153_000, w_153_001;
  wire w_154_034, w_154_098;
  wire w_156_018, w_156_023;
  wire w_157_014, w_157_024;
  wire w_158_056;
  wire w_159_092, w_159_173;
  wire w_161_002, w_161_061, w_161_079;
  wire w_165_060;
  wire w_166_003, w_166_035;
  wire w_167_046, w_167_076, w_167_097;
  wire w_168_000, w_168_002, w_168_004, w_168_006;
  wire w_169_001, w_169_020, w_169_025, w_169_039, w_169_041;
  wire w_170_099, w_170_134;
  wire w_171_021;
  wire w_172_091;
  wire w_173_006;
  wire w_176_076, w_176_166, w_176_167, w_176_168, w_176_169, w_176_170, w_176_171, w_176_172;
  wire w_178_045;
  wire w_179_001;
  wire w_180_034, w_180_037;
  wire w_181_024;
  wire w_183_089;
  wire w_184_112;
  wire w_188_021, w_188_046, w_188_057;
  wire w_190_031;
  wire w_192_011;
  wire w_194_054;
  wire w_195_004;
  wire w_196_042;
  wire w_197_015;
  wire w_200_000, w_200_001, w_200_002, w_200_003, w_200_004, w_200_005, w_200_006, w_200_007, w_200_008, w_200_009, w_200_010, w_200_011, w_200_012, w_200_013, w_200_014, w_200_015, w_200_016, w_200_017, w_200_018, w_200_019, w_200_020, w_200_021, w_200_022, w_200_023, w_200_024, w_200_025, w_200_026, w_200_027, w_200_028, w_200_029, w_200_030, w_200_031, w_200_032, w_200_033, w_200_034, w_200_035, w_200_036, w_200_037, w_200_038, w_200_039, w_200_040, w_200_041, w_200_042, w_200_043, w_200_044, w_200_045, w_200_046, w_200_047, w_200_048, w_200_049, w_200_050, w_200_051, w_200_052, w_200_053, w_200_054, w_200_055, w_200_056, w_200_057, w_200_058, w_200_059, w_200_060, w_200_061, w_200_062, w_200_063, w_200_064, w_200_065, w_200_066, w_200_067, w_200_068, w_200_069, w_200_070, w_200_071, w_200_072, w_200_073, w_200_074, w_200_075, w_200_076, w_200_077, w_200_078, w_200_079, w_200_080, w_200_081, w_200_082, w_200_083, w_200_084, w_200_085, w_200_086, w_200_087;
  not1 I001_000(w_001_000, w_000_000);
  nand2 I001_001(w_001_001, w_000_001, w_000_002);
  not1 I001_002(w_001_002, w_000_003);
  or2  I001_003(w_001_003, w_000_004, w_000_005);
  nand2 I001_004(w_001_004, w_000_006, w_000_007);
  nand2 I001_005(w_001_005, w_000_008, w_000_009);
  not1 I001_006(w_001_006, w_000_010);
  and2 I001_007(w_001_007, w_000_011, w_000_012);
  nand2 I001_008(w_001_008, w_000_013, w_000_014);
  not1 I001_009(w_001_009, w_000_015);
  nand2 I001_010(w_001_010, w_000_016, w_000_017);
  or2  I001_011(w_001_011, w_000_002, w_000_018);
  not1 I001_012(w_001_012, w_000_019);
  nand2 I001_013(w_001_013, w_000_020, w_000_021);
  nand2 I001_014(w_001_014, w_000_022, w_000_023);
  or2  I001_015(w_001_015, w_000_021, w_000_024);
  and2 I001_016(w_001_016, w_000_025, w_000_026);
  and2 I001_017(w_001_017, w_000_027, w_000_028);
  or2  I001_018(w_001_018, w_000_029, w_000_030);
  and2 I002_000(w_002_000, w_001_005, w_000_031);
  or2  I002_001(w_002_001, w_001_011, w_000_032);
  and2 I002_002(w_002_002, w_001_008, w_001_018);
  or2  I002_003(w_002_003, w_000_033, w_000_034);
  not1 I002_004(w_002_004, w_001_015);
  and2 I002_005(w_002_005, w_001_017, w_001_008);
  and2 I002_006(w_002_006, w_000_035, w_000_003);
  nand2 I002_007(w_002_007, w_000_036, w_000_037);
  and2 I002_008(w_002_008, w_000_038, w_000_026);
  not1 I002_009(w_002_009, w_000_039);
  nand2 I002_010(w_002_010, w_000_034, w_000_040);
  or2  I002_011(w_002_011, w_001_007, w_001_016);
  and2 I002_012(w_002_012, w_000_041, w_000_042);
  and2 I002_014(w_002_014, w_001_012, w_001_002);
  nand2 I002_015(w_002_015, w_001_018, w_001_013);
  nand2 I002_016(w_002_016, w_000_043, w_001_015);
  or2  I002_017(w_002_017, w_000_044, w_001_005);
  and2 I002_018(w_002_018, w_001_018, w_001_008);
  nand2 I002_019(w_002_019, w_000_045, w_000_046);
  and2 I002_020(w_002_020, w_001_006, w_001_018);
  or2  I002_021(w_002_021, w_000_047, w_001_003);
  nand2 I002_022(w_002_022, w_000_048, w_000_041);
  not1 I002_023(w_002_023, w_001_005);
  not1 I002_024(w_002_024, w_000_049);
  not1 I002_025(w_002_025, w_001_018);
  nand2 I002_026(w_002_026, w_001_008, w_001_002);
  and2 I002_027(w_002_027, w_000_050, w_001_009);
  nand2 I002_028(w_002_028, w_001_017, w_001_001);
  nand2 I002_029(w_002_029, w_001_018, w_001_003);
  not1 I002_030(w_002_030, w_000_051);
  nand2 I002_031(w_002_031, w_000_052, w_000_004);
  nand2 I002_032(w_002_032, w_001_013, w_000_006);
  and2 I002_033(w_002_033, w_000_018, w_000_053);
  or2  I002_034(w_002_034, w_001_003, w_000_054);
  nand2 I002_035(w_002_035, w_000_055, w_000_056);
  and2 I002_036(w_002_036, w_001_006, w_000_057);
  nand2 I002_037(w_002_037, w_000_058, w_001_006);
  not1 I002_038(w_002_038, w_000_059);
  nand2 I002_039(w_002_039, w_001_004, w_000_011);
  not1 I002_040(w_002_040, w_000_060);
  nand2 I002_041(w_002_041, w_000_061, w_000_022);
  nand2 I002_042(w_002_042, w_000_005, w_001_004);
  not1 I002_043(w_002_043, w_000_062);
  and2 I002_044(w_002_044, w_000_044, w_000_063);
  or2  I002_045(w_002_045, w_000_016, w_000_058);
  and2 I002_046(w_002_046, w_001_005, w_000_000);
  and2 I002_047(w_002_047, w_000_064, w_001_017);
  and2 I002_048(w_002_048, w_001_002, w_001_005);
  not1 I002_049(w_002_049, w_001_018);
  and2 I002_050(w_002_050, w_001_009, w_001_004);
  and2 I002_051(w_002_051, w_001_002, w_001_011);
  not1 I002_052(w_002_052, w_001_012);
  not1 I002_053(w_002_053, w_000_065);
  not1 I002_054(w_002_054, w_000_066);
  not1 I002_055(w_002_055, w_000_067);
  or2  I002_056(w_002_056, w_000_068, w_000_069);
  and2 I002_057(w_002_057, w_000_070, w_001_009);
  and2 I002_058(w_002_058, w_000_071, w_001_006);
  or2  I002_059(w_002_059, w_001_001, w_001_017);
  nand2 I002_060(w_002_060, w_001_007, w_000_072);
  nand2 I002_061(w_002_061, w_000_067, w_001_009);
  nand2 I002_062(w_002_062, w_000_073, w_000_074);
  and2 I002_063(w_002_063, w_000_069, w_000_075);
  not1 I002_064(w_002_064, w_000_076);
  and2 I003_000(w_003_000, w_002_025, w_000_022);
  nand2 I003_001(w_003_001, w_001_004, w_002_048);
  not1 I003_002(w_003_002, w_002_059);
  not1 I003_003(w_003_003, w_002_051);
  nand2 I003_004(w_003_004, w_001_018, w_001_004);
  and2 I003_005(w_003_005, w_002_039, w_000_077);
  not1 I003_006(w_003_006, w_001_003);
  not1 I003_007(w_003_007, w_002_019);
  or2  I003_008(w_003_008, w_001_002, w_001_009);
  or2  I003_009(w_003_009, w_001_002, w_000_059);
  and2 I003_010(w_003_010, w_001_002, w_002_054);
  or2  I003_011(w_003_011, w_000_068, w_000_078);
  and2 I003_012(w_003_012, w_000_079, w_000_036);
  and2 I003_013(w_003_013, w_001_010, w_000_080);
  or2  I003_014(w_003_014, w_002_025, w_000_081);
  not1 I003_015(w_003_015, w_002_064);
  and2 I003_016(w_003_016, w_000_082, w_002_049);
  not1 I003_017(w_003_017, w_001_014);
  nand2 I003_018(w_003_018, w_002_053, w_001_010);
  or2  I003_019(w_003_019, w_002_001, w_001_017);
  or2  I003_020(w_003_020, w_000_036, w_000_014);
  or2  I003_021(w_003_021, w_000_083, w_002_027);
  not1 I003_022(w_003_022, w_002_026);
  not1 I003_023(w_003_023, w_002_032);
  nand2 I003_024(w_003_024, w_001_001, w_002_028);
  nand2 I003_025(w_003_025, w_002_016, w_002_008);
  nand2 I003_026(w_003_026, w_002_005, w_002_009);
  and2 I003_027(w_003_027, w_000_084, w_000_029);
  or2  I003_028(w_003_028, w_000_085, w_001_010);
  nand2 I003_029(w_003_029, w_000_086, w_001_000);
  or2  I003_030(w_003_030, w_000_087, w_001_016);
  nand2 I003_031(w_003_031, w_002_014, w_000_088);
  not1 I003_032(w_003_032, w_002_011);
  not1 I004_000(w_004_000, w_000_061);
  not1 I004_001(w_004_001, w_000_089);
  or2  I004_003(w_004_003, w_000_090, w_001_015);
  not1 I004_004(w_004_004, w_002_059);
  or2  I004_005(w_004_005, w_002_038, w_001_006);
  and2 I004_006(w_004_006, w_002_035, w_002_061);
  not1 I004_007(w_004_007, w_000_091);
  not1 I004_009(w_004_009, w_003_005);
  nand2 I004_010(w_004_010, w_000_031, w_001_000);
  nand2 I004_011(w_004_011, w_000_086, w_002_025);
  and2 I004_012(w_004_012, w_002_012, w_003_010);
  and2 I004_014(w_004_014, w_001_016, w_000_092);
  not1 I004_015(w_004_015, w_002_019);
  and2 I004_016(w_004_016, w_001_006, w_000_049);
  or2  I004_017(w_004_017, w_001_002, w_001_004);
  or2  I004_018(w_004_018, w_003_007, w_002_008);
  nand2 I004_021(w_004_021, w_002_038, w_001_017);
  not1 I004_022(w_004_022, w_001_005);
  or2  I004_023(w_004_023, w_001_006, w_002_034);
  or2  I004_024(w_004_024, w_003_004, w_003_022);
  not1 I004_025(w_004_025, w_001_009);
  nand2 I004_026(w_004_026, w_002_017, w_002_027);
  not1 I004_028(w_004_028, w_003_015);
  not1 I004_030(w_004_030, w_002_033);
  or2  I004_031(w_004_031, w_001_002, w_000_002);
  nand2 I004_032(w_004_032, w_003_031, w_000_093);
  and2 I004_033(w_004_033, w_002_021, w_002_062);
  and2 I004_034(w_004_034, w_003_012, w_001_003);
  and2 I004_035(w_004_035, w_000_083, w_003_027);
  or2  I004_036(w_004_036, w_000_094, w_003_028);
  not1 I004_037(w_004_037, w_000_095);
  not1 I004_038(w_004_038, w_001_011);
  or2  I004_039(w_004_039, w_000_096, w_001_001);
  nand2 I004_040(w_004_040, w_003_023, w_002_059);
  not1 I004_042(w_004_042, w_002_052);
  not1 I004_043(w_004_043, w_001_003);
  not1 I004_044(w_004_044, w_001_010);
  or2  I004_045(w_004_045, w_003_008, w_002_048);
  nand2 I004_046(w_004_046, w_001_010, w_003_022);
  nand2 I004_047(w_004_047, w_002_002, w_002_017);
  not1 I004_048(w_004_048, w_003_005);
  nand2 I004_049(w_004_049, w_001_010, w_001_014);
  or2  I004_050(w_004_050, w_003_011, w_002_017);
  and2 I004_051(w_004_051, w_003_022, w_002_058);
  not1 I004_052(w_004_052, w_000_097);
  or2  I004_053(w_004_053, w_001_009, w_001_016);
  or2  I004_057(w_004_057, w_000_099, w_001_008);
  and2 I004_058(w_004_058, w_003_005, w_002_011);
  not1 I004_059(w_004_059, w_000_100);
  nand2 I004_061(w_004_061, w_002_040, w_003_006);
  not1 I004_062(w_004_062, w_002_063);
  nand2 I004_063(w_004_063, w_002_030, w_001_000);
  nand2 I004_064(w_004_064, w_002_047, w_000_082);
  nand2 I004_065(w_004_065, w_000_004, w_002_043);
  not1 I004_067(w_004_067, w_003_029);
  and2 I004_069(w_004_069, w_003_025, w_000_102);
  or2  I004_071(w_004_071, w_001_014, w_003_011);
  or2  I004_072(w_004_072, w_002_036, w_003_020);
  or2  I004_073(w_004_073, w_003_027, w_000_006);
  or2  I004_074(w_004_074, w_000_084, w_000_103);
  not1 I004_076(w_004_076, w_003_019);
  nand2 I004_077(w_004_077, w_001_007, w_002_010);
  not1 I004_079(w_004_079, w_001_015);
  or2  I004_080(w_004_080, w_002_008, w_001_007);
  and2 I004_082(w_004_082, w_002_016, w_003_017);
  nand2 I004_085(w_004_085, w_000_033, w_002_051);
  or2  I004_088(w_004_088, w_000_106, w_001_011);
  not1 I004_090(w_004_090, w_001_007);
  and2 I004_092(w_004_092, w_002_021, w_002_033);
  or2  I004_094(w_004_094, w_002_060, w_003_015);
  and2 I004_096(w_004_096, w_003_026, w_002_006);
  not1 I004_098(w_004_098, w_001_015);
  and2 I004_104(w_004_104, w_002_063, w_001_014);
  and2 I004_105(w_004_105, w_003_020, w_003_021);
  or2  I004_107(w_004_107, w_001_002, w_000_098);
  not1 I004_110(w_004_110, w_001_003);
  and2 I004_111(w_004_111, w_002_045, w_000_109);
  or2  I004_112(w_004_112, w_003_012, w_003_017);
  or2  I004_115(w_004_115, w_002_042, w_001_002);
  not1 I005_000(w_005_000, w_003_015);
  not1 I005_001(w_005_001, w_001_012);
  and2 I005_003(w_005_003, w_002_007, w_004_028);
  nand2 I005_004(w_005_004, w_000_110, w_001_000);
  or2  I005_005(w_005_005, w_000_111, w_004_000);
  not1 I005_007(w_005_007, w_003_001);
  and2 I005_008(w_005_008, w_004_032, w_004_104);
  nand2 I005_009(w_005_009, w_004_024, w_002_008);
  or2  I005_010(w_005_010, w_001_018, w_001_006);
  and2 I005_011(w_005_011, w_004_014, w_000_112);
  not1 I005_012(w_005_012, w_001_012);
  nand2 I005_013(w_005_013, w_004_018, w_002_021);
  or2  I005_014(w_005_014, w_000_089, w_004_031);
  or2  I005_015(w_005_015, w_004_018, w_003_029);
  or2  I005_016(w_005_016, w_003_000, w_003_017);
  nand2 I005_017(w_005_017, w_000_113, w_003_024);
  and2 I005_018(w_005_018, w_003_023, w_001_000);
  not1 I005_019(w_005_019, w_002_010);
  or2  I005_020(w_005_020, w_001_009, w_000_114);
  nand2 I005_022(w_005_022, w_004_042, w_004_059);
  nand2 I005_023(w_005_023, w_004_044, w_004_038);
  nand2 I005_024(w_005_024, w_001_012, w_004_016);
  nand2 I005_025(w_005_025, w_004_039, w_001_018);
  not1 I005_026(w_005_026, w_001_015);
  and2 I005_027(w_005_027, w_002_064, w_002_003);
  nand2 I005_028(w_005_028, w_002_044, w_002_053);
  and2 I005_029(w_005_029, w_003_012, w_002_007);
  or2  I005_030(w_005_030, w_002_062, w_000_116);
  or2  I005_031(w_005_031, w_001_018, w_001_001);
  not1 I005_032(w_005_032, w_004_063);
  or2  I005_033(w_005_033, w_000_117, w_000_030);
  and2 I005_035(w_005_035, w_004_080, w_001_007);
  not1 I005_036(w_005_036, w_000_119);
  nand2 I005_037(w_005_037, w_004_023, w_003_024);
  not1 I005_038(w_005_038, w_002_028);
  nand2 I005_039(w_005_039, w_000_020, w_000_090);
  or2  I005_040(w_005_040, w_001_000, w_000_021);
  nand2 I005_041(w_005_041, w_004_071, w_000_120);
  nand2 I005_042(w_005_042, w_004_024, w_003_022);
  or2  I005_044(w_005_044, w_000_121, w_000_033);
  nand2 I005_045(w_005_045, w_002_014, w_004_049);
  not1 I005_047(w_005_047, w_001_001);
  or2  I005_048(w_005_048, w_000_122, w_001_011);
  not1 I005_050(w_005_050, w_002_043);
  nand2 I005_051(w_005_051, w_004_025, w_004_044);
  and2 I005_052(w_005_052, w_004_059, w_003_018);
  or2  I005_053(w_005_053, w_002_004, w_000_004);
  or2  I005_054(w_005_054, w_004_017, w_004_115);
  nand2 I005_055(w_005_055, w_002_053, w_004_050);
  nand2 I005_056(w_005_056, w_002_037, w_002_024);
  and2 I005_058(w_005_058, w_001_005, w_004_003);
  nand2 I005_060(w_005_060, w_004_044, w_003_013);
  nand2 I005_061(w_005_061, w_000_045, w_002_057);
  nand2 I005_062(w_005_062, w_001_018, w_001_001);
  not1 I005_063(w_005_063, w_003_029);
  and2 I005_064(w_005_064, w_001_012, w_002_017);
  and2 I005_065(w_005_065, w_001_001, w_000_124);
  not1 I005_066(w_005_066, w_004_006);
  nand2 I005_068(w_005_068, w_002_044, w_000_125);
  and2 I005_069(w_005_069, w_004_028, w_000_022);
  nand2 I005_070(w_005_070, w_000_126, w_004_001);
  and2 I005_071(w_005_071, w_002_041, w_000_125);
  and2 I006_000(w_006_000, w_001_013, w_003_001);
  not1 I006_001(w_006_001, w_000_050);
  and2 I006_002(w_006_002, w_002_003, w_001_015);
  nand2 I006_003(w_006_003, w_004_077, w_004_115);
  or2  I006_004(w_006_004, w_004_039, w_005_063);
  not1 I006_005(w_006_005, w_002_009);
  not1 I006_006(w_006_006, w_005_031);
  nand2 I006_008(w_006_008, w_004_025, w_005_068);
  or2  I006_009(w_006_009, w_000_026, w_002_028);
  nand2 I006_012(w_006_012, w_003_028, w_005_070);
  and2 I006_013(w_006_013, w_005_030, w_004_079);
  or2  I006_015(w_006_015, w_003_020, w_002_050);
  and2 I006_016(w_006_016, w_002_011, w_001_000);
  or2  I006_017(w_006_017, w_005_023, w_004_107);
  or2  I006_018(w_006_018, w_003_005, w_000_127);
  or2  I006_020(w_006_020, w_002_040, w_005_019);
  nand2 I006_021(w_006_021, w_002_008, w_002_034);
  nand2 I006_022(w_006_022, w_001_016, w_003_031);
  nand2 I006_023(w_006_023, w_004_048, w_002_037);
  or2  I006_024(w_006_024, w_003_026, w_005_007);
  nand2 I006_027(w_006_027, w_001_009, w_002_057);
  nand2 I006_028(w_006_028, w_003_005, w_002_064);
  and2 I006_029(w_006_029, w_002_033, w_000_018);
  or2  I006_031(w_006_031, w_001_009, w_000_098);
  or2  I006_032(w_006_032, w_000_128, w_001_014);
  or2  I006_033(w_006_033, w_004_030, w_002_051);
  not1 I006_034(w_006_034, w_000_129);
  or2  I006_035(w_006_035, w_002_023, w_003_000);
  nand2 I006_038(w_006_038, w_003_019, w_000_130);
  or2  I006_043(w_006_043, w_003_000, w_002_000);
  not1 I006_044(w_006_044, w_000_016);
  or2  I006_045(w_006_045, w_001_000, w_005_022);
  nand2 I006_047(w_006_047, w_003_026, w_004_062);
  not1 I006_048(w_006_048, w_003_031);
  and2 I006_049(w_006_049, w_004_080, w_002_045);
  not1 I006_050(w_006_050, w_004_023);
  and2 I006_051(w_006_051, w_004_001, w_001_004);
  not1 I006_053(w_006_053, w_001_010);
  not1 I006_054(w_006_054, w_000_131);
  nand2 I006_055(w_006_055, w_000_034, w_001_006);
  nand2 I006_056(w_006_056, w_002_031, w_004_065);
  or2  I006_058(w_006_058, w_003_028, w_004_064);
  and2 I006_059(w_006_059, w_004_079, w_004_024);
  or2  I006_060(w_006_060, w_000_028, w_001_013);
  not1 I006_061(w_006_061, w_002_005);
  and2 I006_062(w_006_062, w_001_009, w_003_001);
  nand2 I006_065(w_006_065, w_004_094, w_003_013);
  not1 I006_066(w_006_066, w_002_044);
  or2  I006_068(w_006_068, w_005_065, w_002_016);
  or2  I006_069(w_006_069, w_001_004, w_001_002);
  not1 I006_070(w_006_070, w_000_132);
  nand2 I006_072(w_006_072, w_004_011, w_003_022);
  and2 I006_074(w_006_074, w_002_041, w_005_018);
  and2 I006_075(w_006_075, w_002_018, w_002_037);
  or2  I006_078(w_006_078, w_001_014, w_002_017);
  and2 I006_080(w_006_080, w_003_022, w_003_001);
  or2  I006_081(w_006_081, w_004_053, w_004_052);
  and2 I006_083(w_006_083, w_003_026, w_005_005);
  nand2 I006_084(w_006_084, w_000_128, w_005_026);
  and2 I006_086(w_006_086, w_001_016, w_001_004);
  and2 I006_090(w_006_090, w_001_002, w_005_015);
  or2  I006_092(w_006_092, w_003_030, w_002_044);
  not1 I006_093(w_006_093, w_004_012);
  or2  I006_094(w_006_094, w_001_014, w_004_049);
  not1 I006_096(w_006_096, w_005_001);
  not1 I006_097(w_006_097, w_003_013);
  and2 I006_099(w_006_099, w_005_061, w_004_063);
  nand2 I006_100(w_006_100, w_005_003, w_002_055);
  and2 I006_101(w_006_101, w_002_022, w_000_104);
  or2  I006_103(w_006_103, w_002_036, w_004_043);
  not1 I006_104(w_006_104, w_000_135);
  or2  I006_106(w_006_106, w_005_000, w_004_069);
  and2 I006_107(w_006_107, w_001_001, w_000_127);
  or2  I006_109(w_006_109, w_000_136, w_002_044);
  not1 I006_112(w_006_112, w_000_038);
  or2  I006_116(w_006_118, w_005_039, w_006_117);
  nand2 I006_117(w_006_119, w_001_001, w_006_118);
  nand2 I006_118(w_006_120, w_002_051, w_006_119);
  or2  I006_119(w_006_121, w_004_031, w_006_120);
  or2  I006_120(w_006_117, w_006_121, w_005_070);
  not1 I007_000(w_007_000, w_003_020);
  and2 I007_001(w_007_001, w_004_025, w_001_000);
  nand2 I007_002(w_007_002, w_005_000, w_004_021);
  or2  I007_003(w_007_003, w_001_006, w_003_008);
  not1 I007_004(w_007_004, w_006_009);
  nand2 I007_005(w_007_005, w_006_094, w_002_030);
  nand2 I007_006(w_007_006, w_003_021, w_003_022);
  not1 I007_008(w_007_008, w_001_015);
  or2  I007_009(w_007_009, w_006_094, w_003_009);
  and2 I007_010(w_007_010, w_004_028, w_004_005);
  and2 I007_012(w_007_012, w_000_096, w_002_000);
  and2 I007_013(w_007_013, w_005_051, w_004_039);
  or2  I007_014(w_007_014, w_001_010, w_003_028);
  not1 I007_015(w_007_015, w_003_022);
  and2 I007_016(w_007_016, w_006_081, w_006_023);
  not1 I007_017(w_007_017, w_004_014);
  or2  I007_019(w_007_019, w_002_015, w_005_012);
  or2  I007_020(w_007_020, w_002_059, w_003_018);
  and2 I007_021(w_007_021, w_006_092, w_002_028);
  and2 I007_022(w_007_022, w_001_003, w_003_012);
  or2  I007_023(w_007_023, w_000_060, w_005_030);
  nand2 I007_024(w_007_024, w_000_116, w_006_065);
  nand2 I007_025(w_007_025, w_004_017, w_006_059);
  or2  I007_027(w_007_027, w_003_011, w_006_045);
  nand2 I007_029(w_007_029, w_000_137, w_001_002);
  not1 I007_031(w_007_031, w_002_037);
  or2  I007_032(w_007_032, w_006_020, w_006_093);
  or2  I007_033(w_007_033, w_003_020, w_006_012);
  and2 I007_034(w_007_034, w_003_008, w_000_095);
  not1 I007_036(w_007_036, w_004_030);
  nand2 I007_037(w_007_037, w_005_042, w_006_047);
  or2  I007_038(w_007_038, w_003_002, w_001_005);
  nand2 I007_039(w_007_039, w_000_131, w_005_036);
  and2 I007_040(w_007_040, w_001_005, w_003_028);
  and2 I007_041(w_007_041, w_004_001, w_003_003);
  and2 I007_042(w_007_042, w_000_052, w_005_025);
  not1 I007_043(w_007_043, w_000_102);
  or2  I007_044(w_007_044, w_006_033, w_006_035);
  or2  I007_046(w_007_046, w_006_028, w_004_082);
  and2 I007_047(w_007_047, w_005_013, w_003_031);
  not1 I007_048(w_007_048, w_006_068);
  not1 I007_049(w_007_049, w_005_036);
  and2 I007_050(w_007_050, w_003_005, w_000_038);
  and2 I007_051(w_007_051, w_004_022, w_000_035);
  nand2 I007_052(w_007_052, w_001_010, w_001_012);
  not1 I007_053(w_007_053, w_000_078);
  and2 I007_054(w_007_054, w_005_014, w_001_011);
  and2 I007_055(w_006_123, w_007_008, w_006_117);
  or2  I008_000(w_008_000, w_007_012, w_001_000);
  and2 I008_001(w_008_001, w_006_034, w_000_138);
  nand2 I008_002(w_008_002, w_006_065, w_000_049);
  nand2 I008_003(w_008_003, w_003_011, w_006_001);
  not1 I008_004(w_008_004, w_000_139);
  not1 I008_005(w_008_005, w_006_027);
  not1 I008_006(w_008_006, w_004_033);
  or2  I008_008(w_008_008, w_007_004, w_007_040);
  or2  I008_009(w_008_009, w_001_015, w_006_060);
  or2  I008_010(w_008_010, w_007_037, w_007_043);
  or2  I008_012(w_008_012, w_004_096, w_007_001);
  not1 I008_013(w_008_013, w_003_008);
  or2  I008_014(w_008_014, w_001_005, w_002_024);
  not1 I008_015(w_008_015, w_001_003);
  nand2 I008_018(w_008_018, w_004_010, w_004_021);
  or2  I008_020(w_008_020, w_005_050, w_006_006);
  or2  I008_021(w_008_021, w_000_047, w_003_026);
  and2 I008_025(w_008_025, w_006_008, w_002_038);
  or2  I008_026(w_008_026, w_003_027, w_003_001);
  and2 I008_028(w_008_028, w_003_014, w_000_075);
  and2 I008_031(w_008_031, w_005_020, w_000_043);
  and2 I008_033(w_008_033, w_000_096, w_003_004);
  not1 I008_036(w_008_036, w_004_039);
  or2  I008_038(w_008_038, w_007_016, w_003_014);
  and2 I008_039(w_008_039, w_007_041, w_007_044);
  nand2 I008_040(w_008_040, w_002_064, w_002_056);
  or2  I008_044(w_008_044, w_000_130, w_005_003);
  and2 I008_047(w_008_047, w_007_010, w_006_104);
  and2 I008_048(w_008_048, w_000_026, w_006_086);
  or2  I008_049(w_008_049, w_002_016, w_003_004);
  nand2 I008_050(w_008_050, w_005_029, w_001_010);
  and2 I008_051(w_008_051, w_000_069, w_000_071);
  not1 I008_052(w_008_052, w_004_064);
  nand2 I008_054(w_008_054, w_006_123, w_003_023);
  or2  I008_055(w_008_055, w_002_061, w_006_056);
  nand2 I008_056(w_008_056, w_001_015, w_007_039);
  not1 I008_057(w_008_057, w_000_057);
  not1 I008_059(w_008_059, w_000_028);
  and2 I008_062(w_008_062, w_006_044, w_007_000);
  not1 I008_063(w_008_063, w_005_045);
  nand2 I008_064(w_008_064, w_004_046, w_004_038);
  or2  I008_065(w_008_065, w_002_035, w_006_004);
  or2  I008_066(w_008_066, w_004_033, w_005_056);
  not1 I008_069(w_008_069, w_000_140);
  nand2 I008_071(w_008_071, w_003_007, w_007_008);
  or2  I008_075(w_008_075, w_005_017, w_007_053);
  nand2 I008_076(w_008_076, w_000_124, w_003_001);
  and2 I008_078(w_008_078, w_002_032, w_003_030);
  nand2 I008_080(w_008_080, w_002_021, w_006_094);
  or2  I008_081(w_008_081, w_003_017, w_002_017);
  and2 I008_084(w_008_084, w_001_006, w_004_035);
  and2 I008_086(w_008_086, w_002_044, w_001_006);
  and2 I008_088(w_008_088, w_002_020, w_003_024);
  and2 I008_090(w_008_090, w_001_018, w_002_041);
  not1 I008_091(w_008_091, w_003_015);
  not1 I008_093(w_008_093, w_002_012);
  and2 I008_099(w_008_099, w_001_013, w_002_009);
  and2 I008_100(w_008_100, w_006_050, w_000_043);
  or2  I008_104(w_008_104, w_005_037, w_005_008);
  nand2 I008_105(w_008_105, w_000_131, w_004_005);
  and2 I008_108(w_008_108, w_002_018, w_004_004);
  and2 I008_109(w_008_109, w_007_012, w_007_019);
  or2  I008_110(w_008_110, w_005_048, w_006_054);
  or2  I008_112(w_008_112, w_007_038, w_002_058);
  nand2 I008_115(w_008_115, w_003_003, w_006_003);
  and2 I008_120(w_008_120, w_007_002, w_006_016);
  or2  I009_004(w_009_004, w_000_002, w_003_006);
  not1 I009_005(w_009_005, w_004_058);
  and2 I009_006(w_009_006, w_002_016, w_008_120);
  or2  I009_010(w_009_010, w_002_035, w_008_025);
  or2  I009_012(w_009_012, w_007_038, w_005_028);
  not1 I009_015(w_009_015, w_003_010);
  and2 I009_018(w_009_018, w_007_001, w_007_049);
  not1 I009_023(w_009_023, w_006_106);
  or2  I009_026(w_009_026, w_004_018, w_005_032);
  or2  I009_027(w_009_027, w_001_018, w_000_102);
  and2 I009_028(w_009_028, w_002_004, w_002_056);
  not1 I009_030(w_009_030, w_008_075);
  or2  I009_031(w_009_031, w_001_016, w_003_014);
  and2 I009_033(w_009_033, w_002_003, w_000_061);
  and2 I009_034(w_009_034, w_001_013, w_004_036);
  nand2 I009_035(w_009_035, w_007_047, w_008_048);
  or2  I009_037(w_009_037, w_005_010, w_001_004);
  nand2 I009_038(w_009_038, w_000_124, w_004_037);
  not1 I009_040(w_009_040, w_005_070);
  or2  I009_041(w_009_041, w_003_003, w_005_032);
  not1 I009_042(w_009_042, w_000_144);
  not1 I009_043(w_009_043, w_000_145);
  not1 I009_044(w_009_044, w_006_023);
  and2 I009_046(w_009_046, w_005_005, w_001_017);
  or2  I009_047(w_009_047, w_005_048, w_007_050);
  not1 I009_052(w_009_052, w_006_109);
  not1 I009_054(w_009_054, w_008_064);
  and2 I009_055(w_009_055, w_007_029, w_008_065);
  nand2 I009_057(w_009_057, w_005_023, w_003_004);
  nand2 I009_060(w_009_060, w_002_043, w_002_027);
  not1 I009_062(w_009_062, w_003_028);
  nand2 I009_063(w_009_063, w_002_014, w_004_061);
  nand2 I009_064(w_009_064, w_007_043, w_003_011);
  not1 I009_071(w_009_071, w_000_015);
  and2 I009_077(w_009_077, w_006_051, w_002_017);
  not1 I009_078(w_009_078, w_001_003);
  nand2 I009_080(w_009_080, w_001_016, w_000_014);
  nand2 I009_081(w_009_081, w_000_138, w_007_034);
  and2 I009_082(w_009_082, w_003_017, w_006_022);
  not1 I009_083(w_009_083, w_002_014);
  not1 I009_086(w_009_086, w_000_002);
  nand2 I009_089(w_009_089, w_002_039, w_008_002);
  or2  I009_091(w_009_091, w_007_050, w_004_090);
  and2 I009_092(w_009_092, w_007_023, w_004_057);
  nand2 I009_095(w_009_095, w_007_053, w_005_029);
  not1 I009_097(w_009_097, w_006_054);
  not1 I009_105(w_009_105, w_003_030);
  and2 I009_107(w_009_107, w_004_000, w_001_004);
  and2 I009_114(w_009_114, w_001_016, w_002_039);
  and2 I009_117(w_009_117, w_006_049, w_001_016);
  and2 I009_118(w_009_118, w_000_129, w_007_003);
  nand2 I009_122(w_009_122, w_002_007, w_000_150);
  nand2 I009_123(w_009_123, w_007_029, w_001_001);
  not1 I009_125(w_009_125, w_006_021);
  nand2 I009_127(w_009_127, w_005_071, w_005_023);
  not1 I009_134(w_009_134, w_004_105);
  or2  I009_135(w_009_135, w_004_050, w_005_014);
  and2 I009_138(w_009_138, w_000_151, w_002_014);
  nand2 I009_139(w_009_139, w_003_018, w_006_053);
  or2  I010_000(w_010_000, w_004_073, w_001_008);
  and2 I010_002(w_010_002, w_008_057, w_003_030);
  or2  I010_003(w_010_003, w_004_076, w_005_035);
  nand2 I010_004(w_010_004, w_006_005, w_009_005);
  and2 I010_005(w_010_005, w_003_007, w_001_001);
  nand2 I010_006(w_010_006, w_006_075, w_007_036);
  and2 I010_007(w_010_007, w_000_022, w_005_036);
  and2 I010_008(w_010_008, w_001_012, w_009_035);
  and2 I010_009(w_010_009, w_005_009, w_003_027);
  or2  I010_010(w_010_010, w_009_139, w_006_054);
  and2 I010_011(w_010_011, w_004_023, w_000_152);
  not1 I010_012(w_010_012, w_001_004);
  or2  I010_014(w_010_014, w_006_061, w_009_080);
  nand2 I010_015(w_010_015, w_009_057, w_006_050);
  not1 I010_016(w_010_016, w_001_006);
  nand2 I010_017(w_010_017, w_002_049, w_005_024);
  and2 I010_019(w_010_019, w_007_006, w_007_051);
  or2  I010_022(w_010_022, w_006_021, w_008_105);
  or2  I010_023(w_010_023, w_006_080, w_001_006);
  and2 I010_025(w_010_025, w_005_029, w_008_051);
  nand2 I010_026(w_010_026, w_008_055, w_001_010);
  not1 I010_027(w_010_027, w_001_009);
  not1 I010_028(w_010_028, w_000_089);
  and2 I010_029(w_010_029, w_008_062, w_006_024);
  and2 I010_030(w_010_030, w_003_020, w_005_040);
  nand2 I010_032(w_010_032, w_005_004, w_003_018);
  nand2 I010_033(w_010_033, w_001_002, w_008_066);
  and2 I010_034(w_010_034, w_002_062, w_001_013);
  nand2 I010_035(w_010_035, w_007_047, w_006_027);
  not1 I010_037(w_010_037, w_007_040);
  not1 I010_038(w_010_038, w_009_027);
  and2 I010_040(w_010_040, w_008_047, w_008_055);
  or2  I010_042(w_010_042, w_001_015, w_009_054);
  not1 I010_043(w_010_043, w_002_020);
  not1 I010_044(w_010_044, w_000_070);
  or2  I010_046(w_010_046, w_000_154, w_003_005);
  or2  I010_047(w_010_047, w_003_019, w_007_053);
  and2 I010_048(w_010_048, w_005_023, w_001_001);
  or2  I010_049(w_010_049, w_002_009, w_002_016);
  not1 I011_000(w_011_000, w_001_016);
  nand2 I011_002(w_011_002, w_006_090, w_007_042);
  and2 I011_008(w_011_008, w_005_025, w_000_096);
  and2 I011_015(w_011_015, w_004_038, w_001_007);
  not1 I011_016(w_011_016, w_004_069);
  and2 I011_020(w_011_020, w_010_030, w_004_064);
  nand2 I011_023(w_011_023, w_006_097, w_008_021);
  or2  I011_024(w_011_024, w_005_020, w_000_042);
  or2  I011_026(w_011_026, w_003_003, w_001_009);
  and2 I011_029(w_011_029, w_008_038, w_006_016);
  nand2 I011_031(w_011_031, w_004_053, w_009_057);
  and2 I011_032(w_011_032, w_000_034, w_006_021);
  nand2 I011_033(w_011_033, w_007_043, w_009_054);
  not1 I011_034(w_011_034, w_005_033);
  or2  I011_040(w_011_040, w_005_033, w_006_023);
  or2  I011_042(w_011_042, w_004_072, w_009_031);
  not1 I011_043(w_011_043, w_005_052);
  nand2 I011_047(w_011_047, w_003_020, w_000_155);
  and2 I011_050(w_011_050, w_008_004, w_001_008);
  nand2 I011_051(w_011_051, w_004_079, w_006_061);
  not1 I011_052(w_011_052, w_005_018);
  nand2 I011_053(w_011_053, w_000_132, w_005_038);
  nand2 I011_054(w_011_054, w_009_083, w_001_012);
  and2 I011_055(w_011_055, w_007_009, w_009_047);
  nand2 I011_057(w_011_057, w_009_138, w_003_032);
  nand2 I011_060(w_011_060, w_003_023, w_005_001);
  nand2 I011_071(w_011_071, w_005_053, w_006_048);
  and2 I011_072(w_011_072, w_005_022, w_008_000);
  and2 I011_073(w_011_073, w_009_095, w_003_025);
  or2  I011_074(w_011_074, w_007_005, w_007_001);
  not1 I011_077(w_011_077, w_007_036);
  and2 I011_079(w_011_079, w_001_006, w_005_010);
  nand2 I011_080(w_011_080, w_004_001, w_010_040);
  nand2 I011_082(w_011_082, w_006_017, w_002_005);
  or2  I011_085(w_011_085, w_009_028, w_007_036);
  and2 I011_091(w_011_091, w_003_011, w_007_037);
  not1 I011_092(w_011_092, w_001_001);
  nand2 I011_093(w_011_093, w_010_038, w_010_043);
  and2 I011_095(w_011_095, w_002_063, w_006_051);
  not1 I011_101(w_011_101, w_002_003);
  or2  I011_106(w_011_106, w_001_003, w_007_049);
  not1 I011_108(w_011_108, w_008_081);
  not1 I011_113(w_011_113, w_010_006);
  not1 I011_115(w_011_115, w_010_009);
  not1 I011_116(w_011_116, w_009_118);
  nand2 I011_117(w_011_117, w_003_018, w_005_045);
  and2 I011_119(w_011_119, w_010_015, w_003_022);
  not1 I011_122(w_011_122, w_008_012);
  or2  I011_124(w_011_124, w_000_072, w_005_048);
  not1 I011_125(w_011_125, w_004_040);
  and2 I011_128(w_011_128, w_010_047, w_005_044);
  nand2 I011_132(w_011_132, w_008_080, w_000_159);
  and2 I011_133(w_011_133, w_005_020, w_007_012);
  and2 I011_134(w_011_134, w_007_015, w_001_011);
  or2  I011_136(w_011_136, w_000_160, w_007_014);
  or2  I011_137(w_011_137, w_000_109, w_002_027);
  and2 I011_140(w_011_140, w_010_016, w_004_040);
  nand2 I012_000(w_012_000, w_001_010, w_005_033);
  nand2 I012_001(w_012_001, w_004_069, w_003_003);
  nand2 I012_003(w_012_003, w_003_007, w_004_045);
  and2 I012_009(w_012_009, w_009_015, w_003_001);
  and2 I012_010(w_012_010, w_008_014, w_003_024);
  not1 I012_011(w_012_011, w_003_010);
  not1 I012_012(w_012_012, w_009_037);
  and2 I012_013(w_012_013, w_005_028, w_004_046);
  nand2 I012_015(w_012_015, w_001_012, w_002_016);
  and2 I012_016(w_012_016, w_003_026, w_007_024);
  and2 I012_018(w_012_018, w_010_029, w_011_079);
  and2 I012_025(w_012_025, w_011_032, w_002_063);
  or2  I012_027(w_012_027, w_006_100, w_003_000);
  or2  I012_029(w_012_029, w_005_016, w_011_020);
  not1 I012_030(w_012_030, w_000_058);
  nand2 I012_031(w_012_031, w_001_000, w_011_132);
  and2 I012_032(w_012_032, w_005_013, w_008_006);
  not1 I012_033(w_012_033, w_011_073);
  and2 I012_035(w_012_035, w_010_043, w_001_005);
  and2 I012_039(w_012_039, w_006_012, w_008_044);
  or2  I012_043(w_012_043, w_007_021, w_000_161);
  and2 I012_045(w_012_045, w_003_023, w_011_071);
  nand2 I012_048(w_012_048, w_007_002, w_008_069);
  not1 I012_049(w_012_049, w_004_049);
  and2 I012_054(w_012_054, w_000_067, w_010_016);
  nand2 I012_056(w_012_056, w_011_053, w_003_004);
  not1 I012_057(w_012_057, w_006_062);
  or2  I012_067(w_012_067, w_003_013, w_008_056);
  or2  I012_072(w_012_072, w_009_028, w_001_018);
  or2  I012_075(w_012_075, w_008_009, w_009_105);
  or2  I012_078(w_012_078, w_008_049, w_007_023);
  and2 I012_080(w_012_080, w_011_085, w_006_103);
  not1 I012_082(w_012_082, w_005_010);
  or2  I012_084(w_012_084, w_005_018, w_001_002);
  nand2 I012_086(w_012_086, w_004_009, w_003_023);
  not1 I012_087(w_012_087, w_009_078);
  and2 I012_090(w_012_090, w_001_012, w_002_064);
  not1 I012_095(w_012_095, w_006_018);
  or2  I012_103(w_012_103, w_000_021, w_000_045);
  nand2 I012_107(w_012_107, w_006_101, w_008_047);
  nand2 I012_110(w_012_110, w_000_157, w_011_133);
  and2 I012_116(w_012_116, w_005_050, w_010_012);
  not1 I012_119(w_012_119, w_008_008);
  nand2 I012_127(w_012_127, w_004_004, w_000_073);
  nand2 I012_128(w_012_128, w_002_057, w_003_008);
  and2 I013_000(w_013_000, w_005_014, w_003_000);
  or2  I013_001(w_013_001, w_011_055, w_006_075);
  not1 I013_002(w_013_002, w_000_065);
  or2  I013_003(w_013_003, w_012_116, w_007_003);
  not1 I013_008(w_013_008, w_000_162);
  and2 I013_009(w_013_009, w_006_005, w_005_038);
  not1 I013_010(w_013_010, w_004_051);
  not1 I013_012(w_013_012, w_004_036);
  or2  I013_016(w_013_016, w_000_046, w_011_053);
  nand2 I013_017(w_013_017, w_007_000, w_006_043);
  or2  I013_018(w_013_018, w_003_030, w_009_047);
  not1 I013_020(w_013_020, w_002_059);
  or2  I013_021(w_013_021, w_008_025, w_010_033);
  and2 I013_022(w_013_022, w_001_012, w_000_115);
  or2  I013_023(w_013_023, w_000_109, w_006_083);
  and2 I013_024(w_013_024, w_012_078, w_012_010);
  or2  I013_026(w_013_026, w_009_034, w_008_001);
  and2 I013_027(w_013_027, w_010_010, w_004_038);
  not1 I013_030(w_013_030, w_003_027);
  not1 I013_031(w_013_031, w_012_075);
  nand2 I013_032(w_013_032, w_012_013, w_009_010);
  and2 I013_036(w_013_036, w_012_029, w_005_019);
  nand2 I013_037(w_013_037, w_008_001, w_002_040);
  or2  I013_038(w_013_038, w_007_052, w_006_022);
  and2 I013_042(w_013_042, w_001_013, w_003_023);
  or2  I013_044(w_013_044, w_006_065, w_005_027);
  and2 I013_045(w_013_045, w_011_002, w_004_005);
  or2  I013_046(w_013_046, w_008_086, w_000_128);
  or2  I013_047(w_013_047, w_004_085, w_001_015);
  or2  I013_048(w_013_048, w_002_047, w_009_064);
  or2  I013_049(w_013_049, w_000_142, w_012_075);
  or2  I013_050(w_013_050, w_007_022, w_002_036);
  nand2 I013_057(w_013_057, w_010_043, w_003_031);
  nand2 I013_059(w_013_059, w_010_035, w_009_041);
  nand2 I013_060(w_013_060, w_011_029, w_002_019);
  or2  I013_061(w_013_061, w_000_102, w_006_053);
  not1 I013_063(w_013_063, w_007_002);
  or2  I013_064(w_013_064, w_010_038, w_006_054);
  not1 I013_067(w_013_067, w_001_000);
  not1 I013_071(w_013_071, w_009_055);
  or2  I014_004(w_014_004, w_005_014, w_008_063);
  or2  I014_005(w_014_005, w_005_001, w_012_011);
  and2 I014_007(w_014_007, w_006_068, w_011_101);
  nand2 I014_009(w_014_009, w_008_093, w_004_018);
  or2  I014_015(w_014_015, w_003_007, w_012_011);
  nand2 I014_020(w_014_020, w_011_115, w_010_037);
  or2  I014_021(w_014_021, w_008_109, w_002_017);
  or2  I014_030(w_014_030, w_012_067, w_003_012);
  and2 I014_031(w_014_031, w_004_011, w_011_042);
  or2  I014_035(w_014_035, w_006_096, w_009_038);
  nand2 I014_037(w_014_037, w_005_027, w_002_038);
  nand2 I014_038(w_014_038, w_007_002, w_010_028);
  and2 I014_040(w_014_040, w_011_023, w_013_002);
  nand2 I014_042(w_014_042, w_001_005, w_003_029);
  nand2 I014_046(w_014_046, w_003_027, w_011_053);
  not1 I014_047(w_014_047, w_012_027);
  and2 I014_052(w_014_052, w_001_000, w_005_003);
  and2 I014_053(w_014_053, w_003_020, w_008_040);
  or2  I014_055(w_014_055, w_000_027, w_000_056);
  and2 I014_056(w_014_056, w_000_027, w_004_049);
  or2  I014_057(w_014_057, w_012_011, w_000_165);
  or2  I014_058(w_014_058, w_001_003, w_008_050);
  nand2 I014_059(w_014_059, w_006_013, w_003_000);
  or2  I014_064(w_014_064, w_003_001, w_005_050);
  not1 I014_065(w_014_065, w_011_124);
  or2  I014_066(w_014_066, w_001_016, w_000_004);
  and2 I014_070(w_014_070, w_011_117, w_000_078);
  or2  I014_072(w_014_072, w_008_052, w_007_022);
  not1 I014_074(w_014_074, w_008_002);
  not1 I014_077(w_014_077, w_006_004);
  and2 I014_078(w_014_078, w_004_023, w_009_139);
  nand2 I014_080(w_014_080, w_004_090, w_005_041);
  or2  I014_081(w_014_081, w_011_060, w_000_166);
  and2 I014_093(w_014_093, w_009_077, w_006_012);
  and2 I014_100(w_014_100, w_001_008, w_010_002);
  not1 I014_102(w_014_102, w_009_023);
  or2  I014_118(w_014_118, w_008_000, w_012_056);
  or2  I014_121(w_014_121, w_013_071, w_013_061);
  or2  I014_122(w_014_122, w_005_012, w_013_059);
  not1 I014_125(w_014_125, w_010_046);
  nand2 I014_130(w_014_130, w_012_084, w_011_119);
  nand2 I014_139(w_014_139, w_003_019, w_004_011);
  nand2 I015_002(w_015_002, w_014_078, w_014_057);
  nand2 I015_003(w_015_003, w_007_039, w_007_027);
  or2  I015_005(w_015_005, w_002_031, w_008_112);
  or2  I015_012(w_015_012, w_011_050, w_011_000);
  not1 I015_015(w_015_015, w_011_052);
  or2  I015_021(w_015_021, w_002_032, w_003_025);
  or2  I015_022(w_015_022, w_009_043, w_003_029);
  or2  I015_024(w_015_024, w_004_048, w_001_016);
  not1 I015_025(w_015_025, w_006_058);
  or2  I015_027(w_015_027, w_000_013, w_013_023);
  nand2 I015_029(w_015_029, w_013_012, w_009_134);
  nand2 I015_033(w_015_033, w_011_020, w_002_018);
  nand2 I015_034(w_015_034, w_008_115, w_007_034);
  nand2 I015_036(w_015_036, w_002_061, w_004_015);
  not1 I015_037(w_015_037, w_012_057);
  or2  I015_043(w_015_043, w_005_051, w_006_112);
  not1 I015_044(w_015_044, w_011_053);
  and2 I015_047(w_015_047, w_011_092, w_000_094);
  or2  I015_050(w_015_050, w_007_010, w_008_005);
  or2  I015_053(w_015_053, w_013_003, w_010_010);
  nand2 I015_054(w_015_054, w_013_008, w_004_023);
  and2 I015_056(w_015_056, w_012_067, w_000_125);
  and2 I015_057(w_015_057, w_014_052, w_004_059);
  and2 I015_058(w_015_058, w_011_015, w_010_014);
  or2  I015_059(w_015_059, w_014_004, w_009_082);
  or2  I015_062(w_015_062, w_010_025, w_013_042);
  nand2 I015_064(w_015_064, w_012_043, w_014_038);
  nand2 I015_065(w_015_065, w_010_003, w_005_055);
  not1 I015_066(w_015_066, w_004_071);
  and2 I015_076(w_015_076, w_011_053, w_014_139);
  nand2 I015_084(w_015_084, w_013_036, w_011_091);
  and2 I015_085(w_015_085, w_006_038, w_011_140);
  not1 I015_086(w_015_086, w_008_076);
  and2 I015_092(w_015_092, w_000_131, w_011_057);
  and2 I015_106(w_015_106, w_014_077, w_011_074);
  not1 I015_113(w_015_113, w_012_045);
  or2  I015_115(w_015_115, w_011_113, w_004_082);
  or2  I015_118(w_015_118, w_014_009, w_002_064);
  or2  I015_120(w_015_120, w_000_049, w_012_043);
  or2  I015_123(w_015_123, w_012_087, w_009_012);
  not1 I015_126(w_015_126, w_003_023);
  nand2 I016_005(w_016_005, w_002_032, w_014_093);
  and2 I016_007(w_016_007, w_001_007, w_009_018);
  not1 I016_008(w_016_008, w_001_006);
  not1 I016_009(w_016_009, w_011_055);
  not1 I016_012(w_016_012, w_012_015);
  or2  I016_015(w_016_015, w_001_002, w_013_010);
  nand2 I016_016(w_016_016, w_015_012, w_005_010);
  nand2 I016_017(w_016_017, w_004_000, w_004_025);
  not1 I016_021(w_016_021, w_000_005);
  and2 I016_022(w_016_022, w_013_023, w_015_076);
  nand2 I016_023(w_016_023, w_004_065, w_002_063);
  not1 I016_025(w_016_025, w_004_112);
  and2 I016_027(w_016_027, w_006_055, w_002_010);
  not1 I016_029(w_016_029, w_010_027);
  nand2 I016_030(w_016_030, w_010_007, w_015_005);
  or2  I016_031(w_016_031, w_006_016, w_002_002);
  nand2 I016_036(w_016_036, w_000_173, w_010_030);
  nand2 I016_039(w_016_039, w_009_138, w_011_122);
  not1 I016_043(w_016_043, w_010_023);
  and2 I016_045(w_016_045, w_006_048, w_007_031);
  and2 I016_046(w_016_046, w_000_169, w_011_091);
  not1 I016_049(w_016_049, w_004_096);
  and2 I016_050(w_016_050, w_014_121, w_007_043);
  not1 I016_051(w_016_051, w_013_030);
  and2 I016_056(w_016_056, w_006_012, w_008_044);
  and2 I016_065(w_016_065, w_012_095, w_008_033);
  and2 I016_066(w_016_066, w_001_000, w_000_005);
  not1 I016_067(w_016_067, w_005_047);
  nand2 I016_070(w_016_070, w_012_054, w_005_069);
  not1 I016_071(w_016_071, w_007_015);
  not1 I016_073(w_016_073, w_013_010);
  and2 I016_074(w_016_074, w_014_122, w_013_008);
  nand2 I016_075(w_016_075, w_004_064, w_007_033);
  not1 I016_076(w_016_076, w_012_049);
  nand2 I016_079(w_016_079, w_011_015, w_011_057);
  and2 I017_002(w_017_002, w_007_021, w_015_062);
  not1 I017_004(w_017_004, w_009_040);
  and2 I017_006(w_017_006, w_014_021, w_001_005);
  or2  I017_010(w_017_010, w_008_020, w_004_061);
  not1 I017_011(w_017_011, w_013_067);
  and2 I017_022(w_017_022, w_002_028, w_014_056);
  or2  I017_026(w_017_026, w_015_065, w_009_097);
  and2 I017_027(w_017_027, w_008_059, w_000_094);
  nand2 I017_030(w_017_030, w_004_063, w_002_039);
  or2  I017_031(w_017_031, w_008_055, w_003_018);
  and2 I017_032(w_017_032, w_007_052, w_012_010);
  and2 I017_033(w_017_033, w_002_025, w_006_000);
  not1 I017_038(w_017_038, w_007_033);
  nand2 I017_041(w_017_041, w_008_063, w_002_062);
  or2  I017_042(w_017_042, w_012_000, w_005_014);
  or2  I017_045(w_017_045, w_006_048, w_011_072);
  not1 I017_047(w_017_047, w_010_035);
  and2 I017_056(w_017_056, w_016_066, w_008_104);
  nand2 I017_059(w_017_059, w_006_070, w_010_028);
  and2 I017_061(w_017_061, w_015_057, w_015_022);
  and2 I017_065(w_017_065, w_009_046, w_014_118);
  and2 I017_070(w_017_070, w_016_021, w_004_011);
  not1 I017_076(w_017_076, w_007_005);
  nand2 I017_080(w_017_080, w_004_016, w_010_028);
  or2  I017_090(w_017_090, w_013_000, w_013_049);
  not1 I017_097(w_017_097, w_007_013);
  not1 I017_100(w_017_100, w_010_022);
  and2 I017_104(w_017_104, w_005_064, w_001_003);
  and2 I017_107(w_017_107, w_011_125, w_012_015);
  and2 I017_108(w_017_108, w_016_050, w_009_035);
  and2 I017_113(w_017_113, w_000_175, w_001_001);
  and2 I017_134(w_017_134, w_005_004, w_000_070);
  nand2 I018_000(w_018_000, w_001_014, w_002_036);
  nand2 I018_012(w_018_012, w_010_034, w_008_091);
  or2  I018_017(w_018_017, w_002_012, w_009_092);
  nand2 I018_020(w_018_020, w_011_000, w_014_093);
  nand2 I018_023(w_018_023, w_011_016, w_014_081);
  or2  I018_028(w_018_028, w_006_069, w_003_013);
  or2  I018_032(w_018_032, w_016_012, w_008_048);
  nand2 I018_033(w_018_033, w_013_037, w_007_049);
  nand2 I018_035(w_018_035, w_001_005, w_012_039);
  or2  I018_037(w_018_037, w_000_049, w_014_072);
  or2  I018_046(w_018_046, w_002_064, w_014_020);
  and2 I018_051(w_018_051, w_016_046, w_000_000);
  not1 I018_052(w_018_052, w_006_107);
  and2 I018_058(w_018_058, w_000_000, w_007_005);
  not1 I018_059(w_018_059, w_013_024);
  and2 I018_061(w_018_061, w_000_130, w_006_075);
  not1 I018_062(w_018_062, w_017_002);
  or2  I018_064(w_018_064, w_009_082, w_012_103);
  not1 I018_072(w_018_072, w_000_168);
  nand2 I018_073(w_018_073, w_012_072, w_000_116);
  nand2 I018_081(w_018_081, w_000_162, w_017_059);
  not1 I018_082(w_018_082, w_006_069);
  not1 I018_083(w_018_083, w_002_022);
  not1 I018_089(w_018_089, w_007_013);
  not1 I018_110(w_018_110, w_015_085);
  and2 I018_118(w_018_118, w_012_086, w_013_032);
  or2  I018_122(w_018_122, w_013_016, w_017_108);
  and2 I019_003(w_019_003, w_013_024, w_014_055);
  not1 I019_017(w_019_017, w_018_081);
  or2  I019_020(w_019_020, w_014_015, w_008_031);
  nand2 I019_021(w_019_021, w_009_077, w_000_098);
  not1 I019_028(w_019_028, w_011_000);
  and2 I019_033(w_019_033, w_013_042, w_012_012);
  and2 I019_036(w_019_036, w_008_028, w_015_118);
  not1 I019_043(w_019_043, w_005_036);
  nand2 I019_051(w_019_051, w_014_058, w_016_015);
  nand2 I019_052(w_019_052, w_010_006, w_009_122);
  or2  I019_053(w_019_053, w_009_026, w_011_093);
  not1 I019_057(w_019_057, w_014_080);
  and2 I019_071(w_019_071, w_010_023, w_013_067);
  nand2 I019_074(w_019_074, w_005_066, w_002_002);
  nand2 I019_078(w_019_078, w_003_006, w_005_070);
  and2 I019_087(w_019_087, w_016_050, w_006_018);
  not1 I019_091(w_019_091, w_008_026);
  and2 I019_103(w_019_103, w_012_080, w_010_023);
  or2  I019_105(w_019_105, w_008_056, w_001_015);
  nand2 I019_106(w_019_106, w_018_062, w_018_122);
  nand2 I019_111(w_019_111, w_002_012, w_003_009);
  or2  I019_113(w_019_113, w_004_067, w_016_045);
  or2  I019_121(w_019_121, w_003_020, w_010_005);
  not1 I019_124(w_019_124, w_013_000);
  nand2 I019_125(w_019_125, w_015_034, w_004_033);
  and2 I019_126(w_019_126, w_015_059, w_004_098);
  and2 I019_135(w_019_135, w_000_177, w_000_075);
  and2 I019_136(w_019_136, w_000_065, w_002_005);
  nand2 I020_000(w_020_000, w_003_028, w_009_135);
  not1 I020_003(w_020_003, w_000_068);
  not1 I020_004(w_020_004, w_007_032);
  not1 I020_005(w_020_005, w_003_020);
  or2  I020_007(w_020_007, w_008_039, w_012_110);
  and2 I020_008(w_020_008, w_015_025, w_015_065);
  and2 I020_009(w_020_009, w_005_048, w_000_065);
  and2 I020_010(w_020_010, w_007_052, w_017_045);
  and2 I020_011(w_020_011, w_018_000, w_003_002);
  nand2 I020_014(w_020_014, w_018_083, w_007_023);
  and2 I020_015(w_020_015, w_014_130, w_001_005);
  not1 I021_001(w_021_001, w_003_024);
  or2  I021_003(w_021_003, w_020_008, w_013_060);
  nand2 I021_007(w_021_007, w_020_005, w_009_027);
  or2  I021_008(w_021_008, w_013_009, w_009_086);
  or2  I021_011(w_021_011, w_018_033, w_019_051);
  and2 I021_013(w_021_013, w_005_011, w_009_030);
  not1 I021_015(w_021_015, w_011_106);
  and2 I021_023(w_021_023, w_019_017, w_005_069);
  or2  I021_024(w_021_024, w_010_012, w_014_056);
  or2  I021_032(w_021_032, w_005_018, w_008_015);
  and2 I021_036(w_021_036, w_005_036, w_008_005);
  nand2 I021_043(w_021_043, w_016_039, w_019_106);
  or2  I021_044(w_021_044, w_007_033, w_008_078);
  nand2 I021_048(w_021_048, w_009_038, w_000_076);
  and2 I021_051(w_021_051, w_003_029, w_016_008);
  or2  I021_054(w_021_054, w_013_020, w_016_016);
  and2 I021_055(w_021_055, w_010_007, w_013_026);
  not1 I021_080(w_021_080, w_009_089);
  not1 I021_097(w_021_097, w_020_011);
  nand2 I021_108(w_021_108, w_001_014, w_020_010);
  nand2 I021_112(w_021_112, w_014_064, w_016_030);
  nand2 I021_113(w_021_113, w_016_023, w_018_012);
  not1 I021_114(w_021_114, w_015_044);
  not1 I021_121(w_021_121, w_012_027);
  not1 I021_139(w_021_139, w_000_180);
  not1 I021_155(w_021_157, w_021_156);
  and2 I021_156(w_021_158, w_021_157, w_021_176);
  not1 I021_157(w_021_159, w_021_158);
  nand2 I021_158(w_021_160, w_021_159, w_009_134);
  nand2 I021_159(w_021_161, w_021_160, w_016_016);
  and2 I021_160(w_021_162, w_004_074, w_021_161);
  or2  I021_161(w_021_156, w_010_012, w_021_162);
  nand2 I021_162(w_021_167, w_014_066, w_021_166);
  not1 I021_163(w_021_168, w_021_167);
  and2 I021_164(w_021_169, w_011_080, w_021_168);
  not1 I021_165(w_021_170, w_021_169);
  or2  I021_166(w_021_171, w_021_170, w_001_018);
  not1 I021_167(w_021_172, w_021_171);
  not1 I021_168(w_021_173, w_021_172);
  or2  I021_169(w_021_174, w_021_173, w_020_009);
  not1 I021_170(w_021_166, w_021_158);
  and2 I021_171(w_021_176, w_002_049, w_021_174);
  and2 I021_172(w_021_179, w_021_178, w_003_002);
  not1 I021_173(w_021_180, w_021_179);
  and2 I021_174(w_021_181, w_001_003, w_021_180);
  nand2 I021_175(w_021_182, w_021_181, w_020_008);
  or2  I021_176(w_021_183, w_008_071, w_021_182);
  nand2 I021_177(w_021_178, w_021_183, w_002_060);
  or2  I022_000(w_022_000, w_003_031, w_002_006);
  not1 I022_008(w_022_008, w_021_043);
  not1 I022_009(w_022_009, w_001_003);
  and2 I022_015(w_022_015, w_000_145, w_015_027);
  or2  I022_018(w_022_018, w_004_003, w_001_003);
  and2 I022_019(w_022_019, w_008_120, w_008_044);
  not1 I022_022(w_022_022, w_016_071);
  and2 I022_026(w_022_026, w_010_028, w_016_070);
  nand2 I022_027(w_022_027, w_016_007, w_016_029);
  not1 I022_030(w_022_030, w_010_017);
  not1 I022_033(w_022_033, w_012_030);
  or2  I022_034(w_022_034, w_004_044, w_017_056);
  or2  I022_045(w_022_045, w_015_086, w_005_048);
  nand2 I022_054(w_022_054, w_014_040, w_013_064);
  nand2 I022_055(w_022_055, w_016_027, w_008_110);
  not1 I022_071(w_022_071, w_013_057);
  or2  I022_075(w_022_075, w_010_014, w_017_011);
  and2 I022_078(w_022_078, w_006_032, w_000_021);
  not1 I022_079(w_022_079, w_010_042);
  nand2 I022_088(w_022_088, w_002_032, w_001_006);
  and2 I022_094(w_022_094, w_015_092, w_021_097);
  not1 I022_101(w_022_101, w_014_037);
  not1 I023_013(w_023_013, w_014_059);
  not1 I023_015(w_023_015, w_000_052);
  and2 I023_018(w_023_018, w_016_027, w_002_042);
  and2 I023_028(w_023_028, w_011_122, w_002_046);
  or2  I023_030(w_023_030, w_018_020, w_006_028);
  not1 I023_033(w_023_033, w_016_073);
  and2 I023_036(w_023_036, w_022_045, w_000_069);
  not1 I023_038(w_023_038, w_021_055);
  and2 I023_039(w_023_039, w_004_088, w_009_023);
  not1 I023_041(w_023_041, w_000_143);
  nand2 I023_044(w_023_044, w_017_030, w_013_047);
  or2  I023_048(w_023_048, w_007_017, w_019_071);
  and2 I023_053(w_023_053, w_019_033, w_006_059);
  and2 I023_056(w_023_056, w_007_027, w_006_018);
  and2 I023_060(w_023_060, w_011_136, w_018_046);
  not1 I023_061(w_023_061, w_005_008);
  not1 I023_067(w_023_067, w_003_007);
  nand2 I023_087(w_023_087, w_004_007, w_020_010);
  not1 I023_091(w_023_091, w_006_061);
  nand2 I023_098(w_023_098, w_003_027, w_006_028);
  and2 I023_116(w_023_116, w_015_106, w_005_044);
  not1 I023_118(w_023_118, w_005_041);
  not1 I024_000(w_024_000, w_009_052);
  and2 I024_001(w_024_001, w_003_032, w_001_004);
  not1 I024_002(w_024_002, w_018_073);
  or2  I024_003(w_024_003, w_017_042, w_001_004);
  and2 I024_005(w_024_005, w_013_017, w_017_010);
  or2  I024_006(w_024_006, w_019_125, w_016_079);
  or2  I024_008(w_024_008, w_017_004, w_007_020);
  or2  I024_009(w_024_009, w_004_012, w_008_044);
  not1 I024_010(w_024_010, w_020_011);
  nand2 I025_004(w_025_004, w_003_001, w_023_018);
  nand2 I025_009(w_025_009, w_016_071, w_013_022);
  or2  I025_027(w_025_027, w_024_001, w_004_059);
  not1 I025_028(w_025_028, w_017_027);
  and2 I025_033(w_025_033, w_024_001, w_007_043);
  not1 I025_036(w_025_036, w_002_063);
  or2  I025_050(w_025_050, w_009_091, w_023_015);
  nand2 I025_065(w_025_065, w_008_071, w_008_026);
  and2 I025_068(w_025_068, w_010_046, w_021_036);
  nand2 I025_072(w_025_072, w_021_024, w_002_049);
  or2  I025_082(w_025_082, w_014_021, w_008_065);
  and2 I025_087(w_025_087, w_011_034, w_004_031);
  not1 I025_093(w_025_093, w_005_054);
  not1 I025_096(w_025_096, w_018_089);
  or2  I025_106(w_025_106, w_023_056, w_008_075);
  or2  I025_109(w_025_109, w_006_112, w_023_041);
  or2  I025_111(w_025_111, w_005_020, w_003_015);
  or2  I025_123(w_025_123, w_001_012, w_024_006);
  or2  I025_128(w_025_128, w_001_010, w_022_009);
  not1 I025_132(w_025_132, w_009_052);
  nand2 I026_001(w_026_001, w_005_016, w_005_012);
  and2 I026_004(w_026_004, w_019_136, w_022_055);
  or2  I026_005(w_026_005, w_007_014, w_000_082);
  not1 I026_006(w_026_006, w_015_037);
  nand2 I026_012(w_026_012, w_007_008, w_025_027);
  nand2 I026_015(w_026_015, w_006_021, w_018_052);
  or2  I026_017(w_026_017, w_010_014, w_003_031);
  or2  I026_029(w_026_029, w_014_058, w_005_040);
  nand2 I026_035(w_026_035, w_008_008, w_012_031);
  or2  I026_040(w_026_040, w_007_012, w_004_033);
  nand2 I026_042(w_026_042, w_001_016, w_012_119);
  nand2 I026_053(w_026_053, w_015_126, w_011_116);
  nand2 I026_054(w_026_054, w_011_077, w_002_053);
  not1 I026_069(w_026_069, w_001_010);
  nand2 I026_070(w_026_070, w_006_060, w_002_009);
  or2  I026_074(w_026_074, w_005_054, w_015_002);
  not1 I026_077(w_026_077, w_020_009);
  and2 I026_085(w_026_085, w_020_015, w_000_074);
  not1 I026_087(w_026_087, w_014_037);
  and2 I026_088(w_026_088, w_021_001, w_004_034);
  nand2 I026_091(w_026_093, w_021_008, w_026_092);
  or2  I026_092(w_026_094, w_026_093, w_021_139);
  or2  I026_093(w_026_095, w_015_065, w_026_094);
  nand2 I026_094(w_026_092, w_003_021, w_026_095);
  not1 I027_005(w_027_005, w_011_043);
  and2 I027_006(w_027_006, w_001_006, w_001_008);
  not1 I027_014(w_027_014, w_023_091);
  or2  I027_020(w_027_020, w_000_105, w_018_073);
  or2  I027_030(w_027_030, w_025_132, w_009_127);
  and2 I027_031(w_027_031, w_020_015, w_005_039);
  not1 I027_032(w_027_032, w_009_125);
  and2 I027_037(w_027_037, w_017_022, w_026_035);
  not1 I027_043(w_027_043, w_004_007);
  and2 I027_048(w_027_048, w_000_060, w_016_021);
  nand2 I027_050(w_027_050, w_025_072, w_006_031);
  not1 I027_051(w_027_051, w_026_069);
  and2 I027_054(w_027_054, w_017_033, w_026_054);
  or2  I027_055(w_027_055, w_015_050, w_009_077);
  not1 I027_058(w_027_058, w_011_020);
  not1 I027_060(w_027_060, w_009_080);
  nand2 I027_062(w_027_062, w_006_066, w_025_009);
  and2 I027_063(w_027_063, w_011_054, w_021_013);
  and2 I028_000(w_028_000, w_021_113, w_017_076);
  not1 I028_001(w_028_001, w_015_120);
  not1 I028_007(w_028_007, w_017_061);
  or2  I028_009(w_028_009, w_020_010, w_018_028);
  or2  I028_010(w_028_010, w_008_100, w_004_036);
  nand2 I028_011(w_028_011, w_025_111, w_000_186);
  nand2 I028_013(w_028_013, w_006_083, w_009_107);
  and2 I028_018(w_028_018, w_003_011, w_018_035);
  not1 I028_026(w_028_026, w_005_050);
  not1 I028_029(w_028_029, w_007_043);
  not1 I028_034(w_028_034, w_014_074);
  not1 I028_039(w_028_039, w_020_009);
  not1 I028_041(w_028_041, w_000_073);
  or2  I028_045(w_028_045, w_010_010, w_015_054);
  not1 I028_056(w_028_056, w_007_036);
  not1 I028_066(w_028_066, w_011_055);
  and2 I028_070(w_028_070, w_023_028, w_001_015);
  not1 I028_080(w_028_080, w_000_170);
  and2 I028_086(w_028_086, w_010_032, w_016_023);
  and2 I028_087(w_028_087, w_022_088, w_016_065);
  not1 I028_091(w_028_091, w_010_032);
  and2 I028_101(w_028_101, w_009_044, w_003_025);
  not1 I028_113(w_028_113, w_004_096);
  and2 I028_132(w_028_132, w_008_003, w_012_082);
  or2  I028_138(w_028_138, w_005_017, w_010_049);
  nand2 I028_159(w_028_161, w_028_160, w_017_113);
  or2  I028_160(w_028_162, w_028_161, w_015_086);
  not1 I028_161(w_028_163, w_028_162);
  nand2 I028_162(w_028_164, w_028_163, w_004_082);
  nand2 I028_163(w_028_165, w_028_164, w_008_020);
  or2  I028_164(w_028_166, w_015_043, w_028_165);
  nand2 I028_165(w_028_167, w_027_020, w_028_166);
  nand2 I028_166(w_028_168, w_002_054, w_028_167);
  nand2 I028_167(w_028_169, w_028_168, w_007_039);
  or2  I028_168(w_028_160, w_022_075, w_028_169);
  or2  I028_169(w_028_174, w_028_173, w_011_095);
  and2 I028_170(w_028_175, w_020_005, w_028_174);
  not1 I028_171(w_028_176, w_028_175);
  or2  I028_172(w_028_177, w_028_176, w_023_087);
  not1 I028_173(w_028_173, w_028_177);
  and2 I029_000(w_029_000, w_005_070, w_008_108);
  or2  I029_001(w_029_001, w_013_012, w_019_113);
  and2 I029_003(w_029_003, w_010_049, w_003_017);
  not1 I029_004(w_029_004, w_027_048);
  or2  I029_005(w_029_005, w_004_085, w_016_005);
  not1 I029_006(w_029_006, w_017_038);
  not1 I029_007(w_029_007, w_023_060);
  or2  I029_008(w_029_008, w_023_098, w_006_033);
  or2  I029_009(w_029_009, w_020_014, w_017_042);
  and2 I029_010(w_028_171, w_013_044, w_028_160);
  nand2 I029_011(w_029_012, w_016_067, w_029_011);
  and2 I029_012(w_029_013, w_005_058, w_029_012);
  not1 I029_013(w_029_014, w_029_013);
  not1 I029_014(w_029_015, w_029_014);
  not1 I029_015(w_029_016, w_029_015);
  nand2 I029_016(w_029_017, w_027_006, w_029_016);
  not1 I029_017(w_029_018, w_029_017);
  nand2 I029_018(w_029_019, w_029_018, w_028_132);
  not1 I029_019(w_029_020, w_029_019);
  nand2 I029_020(w_029_011, w_029_020, w_002_029);
  and2 I030_003(w_030_003, w_000_012, w_004_064);
  nand2 I030_005(w_030_005, w_021_051, w_028_086);
  and2 I030_022(w_030_022, w_028_171, w_026_074);
  not1 I030_026(w_030_026, w_014_031);
  or2  I030_033(w_030_033, w_006_062, w_007_046);
  nand2 I030_061(w_030_061, w_020_004, w_028_113);
  nand2 I030_063(w_030_063, w_018_059, w_010_028);
  not1 I031_002(w_031_002, w_004_073);
  nand2 I031_005(w_031_005, w_009_006, w_008_014);
  and2 I031_009(w_031_009, w_026_017, w_016_017);
  nand2 I031_014(w_031_014, w_015_021, w_022_027);
  nand2 I031_016(w_031_016, w_005_050, w_029_009);
  or2  I031_021(w_031_021, w_013_001, w_027_014);
  and2 I031_022(w_031_022, w_008_028, w_024_000);
  not1 I031_036(w_031_036, w_008_090);
  nand2 I031_039(w_031_039, w_015_084, w_015_015);
  nand2 I031_044(w_031_044, w_021_013, w_011_079);
  and2 I031_045(w_031_045, w_011_047, w_011_033);
  not1 I031_054(w_031_054, w_010_027);
  not1 I031_057(w_031_057, w_000_115);
  not1 I031_068(w_031_068, w_021_044);
  and2 I031_076(w_031_076, w_014_058, w_030_022);
  nand2 I031_087(w_031_087, w_020_008, w_004_045);
  nand2 I031_089(w_031_089, w_003_023, w_023_030);
  or2  I031_093(w_031_093, w_013_001, w_005_010);
  and2 I031_097(w_031_097, w_020_007, w_027_031);
  or2  I031_103(w_031_103, w_003_003, w_020_014);
  not1 I031_105(w_031_105, w_005_004);
  or2  I031_118(w_031_118, w_019_103, w_014_035);
  and2 I031_129(w_031_129, w_014_046, w_010_019);
  or2  I031_131(w_031_131, w_013_046, w_014_030);
  not1 I031_135(w_031_135, w_007_027);
  not1 I032_001(w_032_001, w_020_004);
  or2  I032_011(w_032_011, w_000_062, w_028_039);
  or2  I032_019(w_032_019, w_020_000, w_004_024);
  nand2 I032_024(w_032_024, w_003_018, w_028_034);
  or2  I032_029(w_032_029, w_000_172, w_005_064);
  not1 I032_033(w_032_033, w_018_023);
  not1 I032_039(w_032_039, w_022_008);
  not1 I032_054(w_032_054, w_008_056);
  or2  I032_062(w_032_062, w_024_009, w_000_189);
  and2 I032_065(w_032_065, w_029_005, w_024_002);
  not1 I032_067(w_032_067, w_010_027);
  and2 I032_069(w_032_069, w_025_123, w_000_056);
  not1 I032_082(w_032_082, w_012_033);
  and2 I032_103(w_032_103, w_009_042, w_029_000);
  and2 I032_105(w_032_105, w_031_045, w_022_018);
  not1 I032_122(w_032_122, w_027_043);
  and2 I033_005(w_033_005, w_032_054, w_031_016);
  not1 I033_006(w_033_006, w_013_063);
  and2 I033_007(w_033_007, w_017_090, w_015_053);
  and2 I033_008(w_033_008, w_013_023, w_028_007);
  nand2 I033_012(w_033_012, w_023_038, w_021_015);
  and2 I033_014(w_033_014, w_008_088, w_015_123);
  and2 I033_018(w_033_018, w_026_035, w_018_037);
  nand2 I033_029(w_033_029, w_013_030, w_005_016);
  and2 I033_030(w_033_030, w_027_063, w_008_040);
  and2 I033_031(w_033_031, w_017_031, w_005_023);
  or2  I033_034(w_033_034, w_002_042, w_032_062);
  or2  I033_035(w_033_035, w_006_075, w_021_003);
  not1 I033_037(w_033_037, w_031_022);
  nand2 I033_040(w_033_040, w_005_033, w_003_023);
  not1 I033_044(w_033_044, w_001_012);
  not1 I033_049(w_033_049, w_032_105);
  not1 I034_001(w_034_001, w_016_025);
  not1 I034_002(w_034_002, w_028_001);
  or2  I034_014(w_034_014, w_005_065, w_011_008);
  or2  I034_017(w_034_017, w_033_018, w_001_006);
  and2 I034_018(w_034_018, w_004_092, w_029_007);
  and2 I034_030(w_034_030, w_021_108, w_033_005);
  not1 I034_041(w_034_041, w_010_023);
  nand2 I034_050(w_034_050, w_016_022, w_028_000);
  or2  I034_065(w_034_065, w_033_012, w_024_000);
  nand2 I034_069(w_034_069, w_029_004, w_029_006);
  and2 I034_072(w_034_072, w_011_082, w_002_052);
  not1 I034_074(w_034_074, w_012_013);
  nand2 I034_088(w_034_088, w_007_048, w_025_096);
  nand2 I034_105(w_034_105, w_014_065, w_002_024);
  nand2 I034_117(w_034_117, w_017_041, w_003_032);
  nand2 I034_128(w_034_128, w_022_009, w_031_068);
  nand2 I034_134(w_034_134, w_032_067, w_022_071);
  or2  I034_136(w_034_136, w_019_087, w_016_073);
  not1 I035_005(w_035_005, w_011_031);
  and2 I035_018(w_035_018, w_017_097, w_005_069);
  not1 I035_027(w_035_027, w_011_024);
  or2  I035_031(w_035_031, w_028_018, w_029_003);
  or2  I035_040(w_035_040, w_018_017, w_033_049);
  nand2 I035_042(w_035_042, w_008_044, w_022_078);
  nand2 I035_044(w_035_044, w_001_006, w_015_085);
  not1 I035_052(w_035_052, w_016_076);
  nand2 I035_057(w_035_057, w_017_006, w_016_008);
  nand2 I035_070(w_035_070, w_003_003, w_002_060);
  and2 I035_073(w_035_073, w_015_043, w_005_042);
  or2  I035_076(w_035_076, w_031_097, w_031_009);
  and2 I035_079(w_035_079, w_016_029, w_007_001);
  and2 I035_082(w_035_082, w_020_000, w_010_006);
  nand2 I035_083(w_035_083, w_018_058, w_034_050);
  or2  I036_000(w_036_000, w_002_054, w_021_121);
  not1 I036_002(w_036_002, w_003_002);
  or2  I036_003(w_036_003, w_021_114, w_001_009);
  not1 I036_004(w_036_004, w_025_068);
  and2 I036_005(w_036_005, w_015_056, w_004_064);
  not1 I036_006(w_036_006, w_005_022);
  or2  I036_008(w_036_008, w_009_081, w_022_022);
  or2  I036_012(w_036_012, w_001_011, w_009_057);
  nand2 I037_000(w_037_000, w_019_121, w_029_009);
  or2  I037_003(w_037_003, w_005_051, w_009_071);
  and2 I037_004(w_037_004, w_028_101, w_001_009);
  nand2 I037_012(w_037_012, w_019_135, w_000_064);
  nand2 I037_075(w_037_075, w_017_070, w_033_007);
  not1 I037_090(w_037_090, w_005_060);
  or2  I037_126(w_037_126, w_021_011, w_016_050);
  or2  I037_128(w_037_128, w_034_014, w_000_178);
  and2 I037_153(w_037_153, w_021_054, w_012_128);
  not1 I038_000(w_038_000, w_013_000);
  not1 I038_002(w_038_002, w_018_051);
  not1 I038_003(w_038_003, w_016_009);
  nand2 I038_004(w_038_004, w_026_054, w_036_000);
  nand2 I038_005(w_038_005, w_035_018, w_003_027);
  or2  I038_006(w_038_006, w_023_048, w_037_000);
  and2 I038_007(w_038_007, w_025_004, w_002_003);
  or2  I038_012(w_038_012, w_017_042, w_018_020);
  or2  I038_013(w_038_013, w_018_118, w_017_107);
  not1 I038_014(w_038_014, w_019_105);
  and2 I038_016(w_038_016, w_004_039, w_007_013);
  not1 I038_017(w_038_017, w_026_069);
  nand2 I038_019(w_038_021, w_009_060, w_038_020);
  or2  I038_020(w_038_022, w_038_021, w_037_128);
  not1 I038_021(w_038_023, w_038_022);
  or2  I038_022(w_038_024, w_038_023, w_021_080);
  or2  I038_023(w_038_020, w_038_024, w_032_039);
  and2 I039_000(w_039_000, w_017_032, w_003_016);
  not1 I039_001(w_039_001, w_038_012);
  not1 I039_002(w_039_002, w_018_028);
  or2  I039_004(w_039_004, w_030_033, w_009_041);
  or2  I039_005(w_039_005, w_036_003, w_023_116);
  not1 I039_006(w_039_006, w_017_047);
  not1 I039_007(w_039_007, w_006_083);
  nand2 I039_011(w_039_012, w_039_011, w_039_036);
  and2 I039_012(w_039_013, w_039_012, w_033_006);
  not1 I039_013(w_039_014, w_039_013);
  and2 I039_014(w_039_015, w_039_014, w_012_090);
  or2  I039_015(w_039_016, w_039_015, w_010_044);
  and2 I039_016(w_039_017, w_039_016, w_010_003);
  not1 I039_017(w_039_018, w_039_017);
  and2 I039_018(w_039_019, w_011_032, w_039_018);
  not1 I039_019(w_039_020, w_039_019);
  not1 I039_020(w_039_021, w_039_020);
  not1 I039_021(w_039_011, w_039_021);
  nand2 I039_022(w_039_026, w_039_025, w_028_010);
  not1 I039_023(w_039_027, w_039_026);
  nand2 I039_024(w_039_028, w_039_027, w_007_013);
  and2 I039_025(w_039_029, w_039_028, w_029_009);
  or2  I039_026(w_039_030, w_039_029, w_023_036);
  or2  I039_027(w_039_031, w_007_013, w_039_030);
  nand2 I039_028(w_039_032, w_035_070, w_039_031);
  and2 I039_029(w_039_033, w_039_032, w_028_066);
  not1 I039_030(w_039_034, w_039_033);
  not1 I039_031(w_039_025, w_039_012);
  and2 I039_032(w_039_036, w_028_138, w_039_034);
  nand2 I040_009(w_040_009, w_026_029, w_022_054);
  nand2 I040_016(w_040_016, w_010_010, w_031_014);
  not1 I040_018(w_040_018, w_013_050);
  and2 I040_037(w_040_037, w_039_005, w_001_004);
  and2 I040_043(w_040_043, w_035_082, w_024_008);
  or2  I040_047(w_040_047, w_026_053, w_000_095);
  not1 I040_053(w_040_053, w_034_088);
  nand2 I040_059(w_040_059, w_013_059, w_012_072);
  nand2 I040_069(w_040_069, w_012_018, w_004_051);
  or2  I040_082(w_040_082, w_008_064, w_010_012);
  or2  I040_106(w_040_106, w_028_034, w_011_128);
  nand2 I040_115(w_040_115, w_003_029, w_013_061);
  or2  I041_023(w_041_023, w_040_037, w_035_079);
  nand2 I041_029(w_041_029, w_023_061, w_035_057);
  and2 I041_035(w_041_035, w_010_048, w_031_005);
  or2  I041_059(w_041_059, w_016_016, w_035_044);
  not1 I041_081(w_041_081, w_013_042);
  not1 I041_116(w_041_116, w_012_025);
  not1 I042_011(w_042_011, w_021_023);
  or2  I042_015(w_042_015, w_006_074, w_031_054);
  not1 I042_016(w_042_016, w_027_062);
  not1 I042_034(w_042_034, w_028_011);
  not1 I042_041(w_042_041, w_004_026);
  or2  I042_049(w_042_049, w_014_038, w_038_000);
  and2 I042_054(w_042_054, w_021_032, w_030_026);
  nand2 I043_016(w_043_016, w_028_013, w_006_084);
  and2 I043_020(w_043_020, w_026_040, w_035_027);
  and2 I043_025(w_043_025, w_036_004, w_029_009);
  not1 I043_030(w_043_030, w_029_007);
  not1 I043_036(w_043_036, w_026_087);
  or2  I043_053(w_043_053, w_028_029, w_036_002);
  or2  I043_062(w_043_062, w_019_052, w_015_043);
  or2  I044_000(w_044_000, w_005_040, w_008_005);
  not1 I044_013(w_044_013, w_028_041);
  nand2 I044_040(w_044_040, w_039_007, w_002_060);
  nand2 I044_058(w_044_058, w_000_115, w_006_086);
  nand2 I044_099(w_044_099, w_006_018, w_017_080);
  and2 I044_139(w_044_139, w_005_013, w_029_000);
  not1 I044_159(w_044_159, w_029_001);
  nand2 I044_161(w_044_161, w_034_030, w_018_061);
  and2 I044_166(w_044_166, w_034_069, w_019_021);
  and2 I044_170(w_044_170, w_013_038, w_005_068);
  nand2 I044_180(w_044_180, w_024_006, w_033_044);
  or2  I045_009(w_045_009, w_013_050, w_040_053);
  and2 I045_013(w_045_013, w_035_044, w_007_054);
  not1 I045_038(w_045_038, w_004_036);
  nand2 I045_039(w_045_039, w_022_034, w_034_041);
  nand2 I045_041(w_045_041, w_024_003, w_026_001);
  nand2 I045_042(w_045_042, w_031_089, w_008_020);
  and2 I045_051(w_045_051, w_007_040, w_006_099);
  or2  I046_010(w_046_010, w_009_114, w_007_012);
  or2  I046_020(w_046_020, w_011_108, w_033_035);
  or2  I046_028(w_046_028, w_024_009, w_029_009);
  and2 I046_030(w_046_030, w_045_041, w_040_069);
  or2  I046_051(w_046_051, w_036_005, w_019_124);
  or2  I046_055(w_046_055, w_034_065, w_020_008);
  not1 I046_056(w_046_056, w_029_005);
  not1 I046_090(w_046_090, w_027_037);
  nand2 I046_092(w_046_092, w_011_060, w_035_042);
  or2  I046_103(w_046_103, w_027_060, w_000_153);
  or2  I046_130(w_046_130, w_027_058, w_009_027);
  and2 I047_006(w_047_006, w_021_112, w_026_006);
  not1 I047_012(w_047_012, w_044_139);
  and2 I047_013(w_047_013, w_031_039, w_002_022);
  nand2 I047_021(w_047_021, w_000_109, w_014_047);
  nand2 I047_027(w_047_027, w_003_004, w_011_093);
  and2 I047_030(w_047_030, w_028_070, w_004_005);
  nand2 I047_033(w_047_033, w_011_026, w_038_000);
  and2 I047_035(w_047_035, w_024_008, w_000_150);
  nand2 I047_048(w_047_048, w_008_080, w_006_078);
  not1 I048_008(w_048_008, w_036_006);
  not1 I048_017(w_048_017, w_003_000);
  nand2 I048_051(w_048_051, w_025_082, w_033_034);
  and2 I048_058(w_048_058, w_022_079, w_011_137);
  and2 I048_076(w_048_076, w_007_039, w_029_008);
  not1 I048_109(w_048_109, w_013_045);
  nand2 I048_136(w_048_136, w_027_030, w_020_011);
  nand2 I048_157(w_048_157, w_019_020, w_008_009);
  or2  I049_008(w_049_008, w_012_003, w_011_082);
  not1 I049_036(w_049_036, w_021_114);
  and2 I049_045(w_049_045, w_035_031, w_016_036);
  or2  I049_046(w_049_046, w_034_001, w_034_128);
  nand2 I049_059(w_049_059, w_044_166, w_029_003);
  not1 I049_069(w_049_069, w_038_017);
  and2 I049_103(w_049_103, w_006_027, w_003_007);
  not1 I049_107(w_049_107, w_019_036);
  and2 I049_125(w_049_125, w_008_020, w_024_008);
  or2  I049_126(w_049_126, w_034_074, w_017_100);
  and2 I049_129(w_049_129, w_046_030, w_042_016);
  not1 I050_006(w_050_006, w_035_005);
  or2  I050_020(w_050_020, w_034_050, w_022_026);
  nand2 I050_025(w_050_025, w_031_021, w_008_084);
  nand2 I050_032(w_050_032, w_003_002, w_011_122);
  nand2 I050_045(w_050_045, w_006_061, w_014_072);
  and2 I050_049(w_050_049, w_046_055, w_031_076);
  not1 I050_054(w_050_054, w_027_005);
  or2  I050_062(w_050_062, w_047_035, w_048_058);
  and2 I050_063(w_050_063, w_004_018, w_047_048);
  and2 I050_069(w_050_069, w_048_136, w_045_038);
  not1 I050_074(w_050_074, w_004_110);
  and2 I050_076(w_050_076, w_023_036, w_032_011);
  or2  I050_096(w_050_096, w_008_099, w_008_018);
  or2  I050_112(w_050_112, w_008_054, w_037_153);
  not1 I050_113(w_050_113, w_040_082);
  and2 I051_006(w_051_006, w_008_078, w_042_011);
  not1 I051_027(w_051_027, w_027_050);
  or2  I051_056(w_051_056, w_005_031, w_031_044);
  and2 I051_122(w_051_122, w_039_004, w_023_013);
  or2  I051_143(w_051_143, w_019_124, w_006_060);
  or2  I052_027(w_052_027, w_015_024, w_019_126);
  and2 I052_031(w_052_031, w_034_018, w_049_046);
  nand2 I052_040(w_052_040, w_029_003, w_037_075);
  and2 I052_050(w_052_050, w_026_004, w_012_016);
  or2  I052_055(w_052_055, w_000_148, w_040_082);
  and2 I053_005(w_053_005, w_008_093, w_022_033);
  not1 I053_012(w_053_012, w_012_048);
  nand2 I053_032(w_053_032, w_049_125, w_043_016);
  and2 I053_033(w_053_033, w_031_036, w_038_016);
  or2  I053_045(w_053_045, w_047_030, w_013_067);
  not1 I053_065(w_053_065, w_031_131);
  and2 I054_000(w_054_000, w_045_009, w_041_059);
  and2 I054_001(w_054_001, w_001_012, w_023_039);
  and2 I054_002(w_054_002, w_002_047, w_034_117);
  and2 I054_003(w_054_003, w_002_020, w_050_032);
  and2 I054_004(w_054_004, w_010_004, w_030_022);
  or2  I054_005(w_054_005, w_038_004, w_000_032);
  not1 I054_008(w_054_008, w_004_050);
  not1 I054_009(w_054_009, w_038_005);
  nand2 I055_015(w_055_015, w_038_006, w_005_016);
  or2  I055_024(w_055_024, w_027_062, w_033_031);
  or2  I055_035(w_055_035, w_001_002, w_010_000);
  and2 I055_077(w_055_077, w_040_018, w_009_043);
  and2 I055_087(w_055_087, w_024_002, w_001_016);
  nand2 I055_132(w_055_132, w_053_012, w_042_054);
  or2  I055_177(w_055_177, w_028_080, w_051_143);
  and2 I056_001(w_056_001, w_010_027, w_000_122);
  or2  I056_014(w_056_014, w_023_033, w_028_056);
  and2 I056_018(w_056_018, w_003_030, w_000_100);
  nand2 I056_058(w_056_058, w_004_048, w_011_125);
  and2 I056_070(w_056_070, w_051_006, w_018_064);
  not1 I056_074(w_056_074, w_020_004);
  or2  I056_099(w_056_099, w_030_003, w_033_040);
  and2 I056_103(w_056_103, w_037_126, w_044_170);
  and2 I056_104(w_056_104, w_039_001, w_054_004);
  nand2 I057_026(w_057_026, w_011_122, w_006_002);
  or2  I057_031(w_057_031, w_049_059, w_049_036);
  nand2 I057_051(w_057_051, w_010_026, w_044_159);
  or2  I057_083(w_057_083, w_050_020, w_025_065);
  nand2 I058_000(w_058_000, w_050_113, w_046_051);
  nand2 I058_018(w_058_018, w_045_013, w_054_002);
  or2  I058_019(w_058_019, w_052_050, w_010_033);
  not1 I058_028(w_058_028, w_001_000);
  not1 I058_031(w_058_031, w_038_004);
  and2 I058_036(w_058_036, w_029_003, w_014_053);
  not1 I058_039(w_058_039, w_050_025);
  and2 I058_067(w_058_067, w_050_076, w_009_063);
  nand2 I058_069(w_058_069, w_024_010, w_056_018);
  and2 I058_072(w_058_072, w_040_115, w_003_021);
  not1 I058_089(w_058_089, w_022_088);
  not1 I059_011(w_059_011, w_038_006);
  not1 I059_039(w_059_039, w_056_104);
  and2 I059_046(w_059_046, w_042_049, w_043_025);
  and2 I059_058(w_059_058, w_025_033, w_002_059);
  and2 I059_065(w_059_065, w_008_044, w_022_094);
  not1 I059_070(w_059_070, w_030_022);
  nand2 I059_073(w_059_073, w_010_008, w_007_020);
  nand2 I059_085(w_059_085, w_031_118, w_019_078);
  not1 I059_097(w_059_097, w_001_017);
  or2  I059_117(w_059_117, w_056_014, w_017_004);
  not1 I059_134(w_059_134, w_003_007);
  or2  I059_163(w_059_163, w_005_039, w_042_034);
  and2 I060_006(w_060_006, w_031_087, w_043_030);
  not1 I060_007(w_060_007, w_005_062);
  not1 I060_029(w_060_029, w_019_121);
  or2  I060_030(w_060_030, w_058_019, w_038_002);
  or2  I060_044(w_060_044, w_054_009, w_050_006);
  not1 I060_045(w_060_045, w_012_035);
  nand2 I060_049(w_060_049, w_032_067, w_028_091);
  or2  I060_061(w_060_061, w_015_115, w_015_058);
  nand2 I061_003(w_061_003, w_006_093, w_009_031);
  not1 I061_035(w_061_035, w_008_020);
  and2 I061_072(w_061_072, w_059_070, w_024_005);
  and2 I061_096(w_061_096, w_054_000, w_048_008);
  nand2 I062_003(w_062_003, w_033_012, w_037_004);
  and2 I062_060(w_062_060, w_055_024, w_017_026);
  or2  I062_125(w_062_125, w_006_029, w_030_005);
  nand2 I062_127(w_062_127, w_037_003, w_017_065);
  not1 I062_194(w_062_194, w_060_045);
  or2  I063_007(w_063_007, w_044_040, w_031_036);
  nand2 I063_010(w_063_010, w_016_074, w_020_010);
  nand2 I063_029(w_063_029, w_014_042, w_020_003);
  not1 I063_068(w_063_068, w_024_008);
  not1 I063_078(w_063_078, w_048_051);
  nand2 I064_028(w_064_028, w_029_005, w_038_017);
  not1 I064_035(w_064_035, w_014_031);
  and2 I064_037(w_064_037, w_019_003, w_016_021);
  not1 I064_070(w_064_070, w_022_015);
  and2 I064_079(w_064_079, w_029_003, w_054_003);
  not1 I064_130(w_064_130, w_052_031);
  not1 I064_144(w_064_144, w_055_132);
  or2  I064_152(w_064_152, w_012_032, w_043_020);
  and2 I064_165(w_064_165, w_046_020, w_050_045);
  or2  I065_004(w_065_004, w_054_008, w_013_018);
  or2  I065_037(w_065_037, w_049_103, w_038_007);
  nand2 I065_062(w_065_062, w_031_057, w_036_000);
  and2 I065_064(w_065_064, w_052_055, w_058_018);
  not1 I066_011(w_066_011, w_020_009);
  or2  I066_065(w_066_065, w_032_019, w_049_107);
  not1 I066_088(w_066_088, w_017_104);
  or2  I066_126(w_066_126, w_041_029, w_033_029);
  and2 I066_138(w_066_138, w_000_080, w_055_035);
  and2 I066_156(w_066_156, w_061_072, w_065_037);
  or2  I067_022(w_067_022, w_026_088, w_033_030);
  not1 I067_028(w_067_028, w_041_116);
  and2 I067_046(w_067_046, w_002_024, w_015_092);
  not1 I067_047(w_067_047, w_020_010);
  and2 I068_018(w_068_018, w_032_001, w_000_115);
  nand2 I068_029(w_068_029, w_052_040, w_023_060);
  or2  I068_035(w_068_035, w_046_028, w_008_010);
  or2  I068_046(w_068_046, w_022_000, w_039_001);
  or2  I069_100(w_069_100, w_063_029, w_065_037);
  and2 I069_133(w_069_133, w_003_026, w_027_030);
  and2 I069_155(w_069_155, w_007_029, w_022_019);
  or2  I070_026(w_070_026, w_047_013, w_058_036);
  and2 I070_044(w_070_044, w_052_027, w_017_134);
  not1 I070_055(w_070_055, w_059_163);
  not1 I070_062(w_070_062, w_016_051);
  nand2 I070_082(w_070_084, w_070_083, w_033_037);
  or2  I070_083(w_070_085, w_070_084, w_050_054);
  nand2 I070_084(w_070_086, w_069_100, w_070_085);
  or2  I070_085(w_070_087, w_025_033, w_070_086);
  nand2 I070_086(w_070_088, w_019_087, w_070_087);
  and2 I070_087(w_070_089, w_070_088, w_018_032);
  nand2 I070_088(w_070_090, w_039_006, w_070_089);
  or2  I070_089(w_070_091, w_070_090, w_013_048);
  and2 I070_090(w_070_083, w_044_058, w_070_091);
  or2  I071_007(w_071_007, w_013_021, w_032_122);
  and2 I071_017(w_071_017, w_016_056, w_029_005);
  not1 I071_028(w_071_028, w_036_000);
  or2  I071_076(w_071_076, w_003_005, w_048_017);
  and2 I071_129(w_070_093, w_018_000, w_070_083);
  nand2 I072_051(w_072_051, w_056_104, w_025_093);
  or2  I072_096(w_072_096, w_070_093, w_047_033);
  nand2 I072_103(w_072_103, w_026_015, w_070_062);
  or2  I072_150(w_072_150, w_005_023, w_009_035);
  not1 I073_009(w_073_009, w_026_077);
  or2  I073_015(w_073_015, w_048_109, w_001_014);
  or2  I073_025(w_073_025, w_035_040, w_036_006);
  or2  I073_062(w_073_062, w_001_013, w_028_087);
  not1 I074_069(w_074_069, w_059_065);
  or2  I074_087(w_074_087, w_066_138, w_039_007);
  and2 I074_136(w_074_136, w_063_078, w_049_045);
  and2 I074_138(w_074_138, w_067_028, w_066_156);
  and2 I075_023(w_075_023, w_050_096, w_038_014);
  and2 I075_036(w_075_036, w_065_004, w_073_062);
  nand2 I076_008(w_076_008, w_058_069, w_019_074);
  or2  I076_023(w_076_023, w_032_024, w_015_047);
  and2 I076_156(w_076_156, w_012_009, w_001_015);
  or2  I076_167(w_076_167, w_064_144, w_056_099);
  not1 I077_017(w_077_017, w_015_066);
  or2  I077_019(w_077_019, w_003_006, w_046_103);
  or2  I077_031(w_077_031, w_039_004, w_025_050);
  or2  I077_032(w_077_032, w_024_008, w_066_088);
  or2  I078_010(w_078_010, w_043_053, w_039_002);
  and2 I078_015(w_078_015, w_006_083, w_063_007);
  and2 I078_024(w_078_024, w_003_009, w_045_009);
  nand2 I078_026(w_078_026, w_055_077, w_049_008);
  or2  I078_043(w_078_043, w_056_070, w_053_033);
  nand2 I078_070(w_078_070, w_003_010, w_028_026);
  not1 I079_003(w_079_003, w_019_111);
  or2  I079_004(w_079_004, w_038_003, w_047_027);
  not1 I079_008(w_079_008, w_034_002);
  and2 I079_009(w_079_009, w_077_019, w_068_046);
  and2 I080_001(w_080_001, w_004_018, w_034_072);
  not1 I080_008(w_080_008, w_023_067);
  and2 I080_024(w_080_024, w_060_007, w_015_003);
  and2 I080_032(w_080_032, w_070_044, w_074_069);
  and2 I080_036(w_080_036, w_078_026, w_032_065);
  and2 I081_017(w_081_017, w_066_065, w_009_114);
  not1 I081_026(w_081_026, w_060_006);
  not1 I081_027(w_081_027, w_001_007);
  and2 I081_054(w_081_054, w_016_076, w_049_069);
  or2  I081_091(w_081_091, w_015_113, w_038_000);
  nand2 I082_008(w_082_008, w_021_007, w_007_013);
  or2  I082_012(w_082_012, w_058_067, w_007_032);
  or2  I082_020(w_082_020, w_054_001, w_022_101);
  and2 I082_051(w_082_051, w_081_026, w_055_087);
  and2 I082_061(w_082_061, w_011_134, w_045_051);
  nand2 I082_063(w_082_063, w_019_053, w_005_054);
  nand2 I083_012(w_083_012, w_050_063, w_057_031);
  nand2 I083_036(w_083_036, w_025_028, w_018_072);
  or2  I083_059(w_083_059, w_078_043, w_077_032);
  and2 I083_069(w_083_069, w_015_029, w_064_130);
  or2  I084_015(w_084_015, w_083_036, w_017_002);
  or2  I084_028(w_084_028, w_051_122, w_059_046);
  not1 I084_036(w_084_036, w_040_106);
  not1 I084_079(w_084_079, w_009_033);
  or2  I085_015(w_085_015, w_012_018, w_056_074);
  and2 I085_044(w_085_044, w_055_177, w_007_036);
  and2 I086_026(w_086_026, w_046_092, w_003_004);
  not1 I086_029(w_086_029, w_053_045);
  not1 I086_035(w_086_035, w_047_006);
  and2 I087_016(w_087_016, w_041_023, w_019_043);
  or2  I087_032(w_087_032, w_046_130, w_076_156);
  and2 I088_005(w_088_005, w_031_039, w_083_059);
  and2 I088_033(w_088_033, w_086_026, w_059_039);
  and2 I089_016(w_089_016, w_086_029, w_026_042);
  nand2 I089_020(w_089_020, w_064_028, w_078_010);
  not1 I089_033(w_089_033, w_071_028);
  not1 I089_039(w_089_039, w_009_023);
  not1 I090_015(w_090_015, w_007_029);
  nand2 I090_020(w_090_020, w_045_039, w_023_033);
  or2  I090_029(w_090_029, w_079_004, w_032_082);
  not1 I090_069(w_090_069, w_051_056);
  not1 I091_011(w_091_011, w_042_041);
  or2  I091_100(w_091_100, w_010_011, w_002_039);
  not1 I091_148(w_091_148, w_062_125);
  not1 I092_038(w_092_038, w_035_052);
  and2 I092_053(w_092_053, w_026_004, w_004_111);
  not1 I092_109(w_092_109, w_025_106);
  or2  I092_121(w_092_121, w_040_016, w_058_000);
  or2  I093_030(w_093_030, w_014_005, w_083_059);
  or2  I093_042(w_093_042, w_092_038, w_054_003);
  nand2 I094_075(w_094_075, w_009_004, w_092_109);
  nand2 I094_080(w_094_080, w_032_103, w_068_029);
  not1 I094_084(w_094_084, w_047_013);
  and2 I094_086(w_094_086, w_040_059, w_025_036);
  not1 I096_009(w_096_009, w_053_065);
  not1 I096_015(w_096_015, w_075_023);
  nand2 I096_016(w_096_016, w_009_062, w_000_016);
  nand2 I096_023(w_096_023, w_031_129, w_002_008);
  or2  I097_003(w_097_003, w_054_002, w_016_049);
  nand2 I097_018(w_097_018, w_076_008, w_034_105);
  not1 I097_020(w_097_020, w_009_123);
  not1 I097_054(w_097_054, w_022_030);
  not1 I097_055(w_097_055, w_039_000);
  not1 I097_056(w_097_056, w_067_046);
  not1 I098_036(w_098_036, w_019_028);
  and2 I098_077(w_098_077, w_090_020, w_094_075);
  or2  I098_079(w_098_079, w_072_051, w_038_002);
  not1 I099_029(w_099_029, w_034_136);
  not1 I100_002(w_100_002, w_054_002);
  not1 I100_018(w_100_018, w_026_085);
  or2  I100_019(w_100_019, w_025_087, w_032_033);
  nand2 I100_020(w_100_020, w_030_003, w_040_009);
  nand2 I101_001(w_101_001, w_100_018, w_073_015);
  not1 I101_005(w_101_005, w_088_033);
  or2  I101_025(w_101_025, w_006_001, w_043_036);
  not1 I102_079(w_102_079, w_082_020);
  or2  I102_104(w_102_104, w_056_001, w_082_063);
  and2 I102_135(w_102_135, w_072_096, w_076_167);
  not1 I103_013(w_103_013, w_019_091);
  or2  I103_094(w_103_094, w_050_112, w_041_035);
  not1 I103_127(w_103_127, w_000_097);
  and2 I103_138(w_103_138, w_004_047, w_085_044);
  and2 I104_104(w_104_104, w_097_054, w_007_049);
  nand2 I104_119(w_104_119, w_054_004, w_077_017);
  nand2 I105_182(w_105_182, w_012_001, w_001_011);
  not1 I106_000(w_106_000, w_087_032);
  or2  I106_008(w_106_008, w_005_064, w_097_018);
  and2 I107_013(w_107_013, w_087_016, w_102_104);
  not1 I107_019(w_107_019, w_010_046);
  not1 I107_063(w_107_063, w_023_067);
  and2 I107_152(w_107_152, w_097_003, w_026_070);
  nand2 I108_023(w_108_023, w_029_009, w_083_069);
  or2  I108_027(w_108_027, w_064_152, w_065_062);
  nand2 I109_069(w_109_069, w_082_012, w_098_036);
  and2 I109_075(w_109_075, w_089_016, w_016_043);
  not1 I109_106(w_109_106, w_005_007);
  not1 I109_122(w_109_122, w_062_127);
  or2  I110_022(w_110_022, w_062_003, w_073_009);
  nand2 I111_008(w_111_008, w_038_000, w_081_091);
  or2  I111_011(w_111_011, w_076_023, w_110_022);
  nand2 I111_039(w_111_039, w_074_138, w_028_045);
  nand2 I112_061(w_112_061, w_092_053, w_097_056);
  not1 I112_075(w_112_075, w_003_003);
  or2  I112_089(w_112_089, w_033_008, w_070_026);
  or2  I113_001(w_113_001, w_064_037, w_104_104);
  nand2 I114_053(w_114_053, w_098_077, w_034_014);
  nand2 I114_099(w_114_101, w_114_100, w_031_093);
  and2 I114_100(w_114_102, w_109_106, w_114_101);
  or2  I114_101(w_114_103, w_114_102, w_060_030);
  not1 I114_102(w_114_100, w_114_103);
  nand2 I114_103(w_114_108, w_114_107, w_054_000);
  not1 I114_104(w_114_109, w_114_108);
  and2 I114_105(w_114_110, w_114_109, w_077_031);
  not1 I114_106(w_114_111, w_114_110);
  and2 I114_107(w_114_112, w_114_111, w_005_063);
  and2 I114_108(w_114_113, w_014_070, w_114_112);
  nand2 I114_109(w_114_114, w_114_113, w_070_055);
  not1 I114_110(w_114_115, w_114_114);
  or2  I114_111(w_114_107, w_114_115, w_093_030);
  nand2 I115_011(w_115_011, w_028_009, w_092_121);
  or2  I117_000(w_117_000, w_060_044, w_084_036);
  nand2 I117_001(w_117_001, w_084_028, w_107_063);
  nand2 I118_025(w_118_025, w_035_044, w_108_023);
  and2 I118_030(w_118_030, w_090_029, w_048_076);
  not1 I118_066(w_118_066, w_067_022);
  nand2 I119_006(w_119_006, w_064_035, w_118_066);
  or2  I119_011(w_119_011, w_058_072, w_079_003);
  not1 I120_011(w_120_011, w_025_109);
  or2  I120_172(w_120_172, w_108_027, w_084_015);
  or2  I121_013(w_121_013, w_107_013, w_040_043);
  and2 I122_028(w_122_028, w_105_182, w_081_027);
  and2 I122_059(w_122_059, w_016_075, w_048_157);
  or2  I123_000(w_123_000, w_045_042, w_004_016);
  not1 I123_044(w_123_044, w_091_148);
  not1 I123_108(w_123_108, w_032_122);
  nand2 I124_047(w_124_047, w_026_005, w_117_001);
  nand2 I126_001(w_126_001, w_027_055, w_120_172);
  and2 I126_002(w_126_002, w_083_012, w_082_061);
  nand2 I127_005(w_127_005, w_060_029, w_031_135);
  and2 I128_022(w_128_022, w_126_001, w_101_025);
  or2  I129_002(w_129_002, w_066_126, w_111_039);
  and2 I129_036(w_129_036, w_127_005, w_096_023);
  nand2 I130_051(w_130_051, w_112_075, w_059_085);
  or2  I130_117(w_130_117, w_041_081, w_002_011);
  and2 I130_176(w_130_176, w_101_005, w_020_003);
  not1 I131_037(w_131_037, w_011_040);
  nand2 I131_101(w_131_101, w_100_020, w_085_015);
  not1 I132_041(w_132_041, w_059_117);
  or2  I132_052(w_132_054, w_009_080, w_132_053);
  and2 I132_053(w_132_055, w_132_054, w_101_001);
  or2  I132_054(w_132_056, w_067_047, w_132_055);
  not1 I132_055(w_132_057, w_132_056);
  or2  I132_056(w_132_058, w_132_057, w_046_010);
  or2  I132_057(w_132_059, w_103_094, w_132_058);
  or2  I132_058(w_132_060, w_109_069, w_132_059);
  not1 I132_059(w_132_061, w_132_060);
  nand2 I132_060(w_132_062, w_132_061, w_097_055);
  nand2 I132_061(w_132_063, w_047_021, w_132_062);
  and2 I132_062(w_132_053, w_132_063, w_012_127);
  not1 I133_007(w_133_007, w_050_062);
  and2 I133_012(w_133_012, w_019_057, w_044_180);
  or2  I133_038(w_133_038, w_081_054, w_018_110);
  and2 I133_143(w_133_143, w_057_051, w_013_024);
  and2 I133_152(w_132_065, w_106_008, w_132_053);
  nand2 I133_153(w_133_154, w_075_036, w_133_153);
  nand2 I133_154(w_133_155, w_133_154, w_106_000);
  nand2 I133_155(w_133_156, w_032_029, w_133_155);
  nand2 I133_156(w_133_157, w_133_156, w_072_103);
  nand2 I133_157(w_133_158, w_133_157, w_015_064);
  or2  I133_158(w_133_159, w_133_158, w_078_024);
  not1 I133_159(w_133_160, w_133_159);
  and2 I133_160(w_133_161, w_133_160, w_096_015);
  not1 I133_161(w_133_162, w_133_161);
  nand2 I133_162(w_133_163, w_036_006, w_133_162);
  not1 I133_163(w_133_164, w_133_163);
  and2 I133_164(w_133_153, w_133_164, w_053_032);
  nand2 I134_007(w_134_007, w_074_136, w_011_002);
  nand2 I134_020(w_134_020, w_132_065, w_037_090);
  or2  I135_079(w_135_079, w_036_003, w_103_138);
  not1 I136_034(w_136_034, w_079_008);
  or2  I137_005(w_137_005, w_008_055, w_120_011);
  or2  I138_132(w_138_132, w_074_087, w_123_044);
  or2  I138_148(w_138_148, w_132_041, w_015_036);
  and2 I139_031(w_139_031, w_038_004, w_039_007);
  nand2 I140_044(w_140_044, w_091_011, w_062_194);
  and2 I141_004(w_141_004, w_032_069, w_137_005);
  nand2 I142_002(w_142_002, w_007_025, w_059_011);
  not1 I142_006(w_142_006, w_111_008);
  nand2 I143_001(w_143_001, w_091_100, w_049_126);
  and2 I144_036(w_144_036, w_082_008, w_090_069);
  or2  I144_052(w_144_052, w_058_039, w_008_013);
  not1 I144_096(w_144_096, w_068_035);
  nand2 I144_197(w_144_199, w_093_042, w_144_198);
  not1 I144_198(w_144_200, w_144_199);
  not1 I144_199(w_144_201, w_144_200);
  and2 I144_200(w_144_202, w_144_201, w_144_213);
  and2 I144_201(w_144_203, w_144_202, w_057_083);
  not1 I144_202(w_144_204, w_144_203);
  nand2 I144_203(w_144_198, w_144_204, w_016_031);
  not1 I144_204(w_144_209, w_144_208);
  nand2 I144_205(w_144_210, w_144_209, w_059_073);
  or2  I144_206(w_144_211, w_144_210, w_061_096);
  not1 I144_207(w_144_208, w_144_202);
  and2 I144_208(w_144_213, w_088_005, w_144_211);
  or2  I145_004(w_145_004, w_034_134, w_037_012);
  not1 I145_013(w_145_013, w_002_006);
  or2  I146_018(w_146_018, w_010_007, w_072_150);
  and2 I146_126(w_146_126, w_133_007, w_098_079);
  not1 I147_016(w_147_016, w_008_006);
  and2 I147_061(w_147_061, w_136_034, w_119_011);
  nand2 I147_080(w_147_080, w_146_018, w_082_051);
  not1 I149_015(w_149_015, w_021_044);
  nand2 I149_019(w_149_019, w_033_030, w_099_029);
  not1 I150_007(w_150_009, w_150_008);
  not1 I150_008(w_150_010, w_150_009);
  or2  I150_009(w_150_011, w_006_015, w_150_010);
  not1 I150_010(w_150_012, w_150_011);
  not1 I150_011(w_150_013, w_150_012);
  and2 I150_012(w_150_014, w_150_013, w_060_049);
  nand2 I150_013(w_150_015, w_150_014, w_130_176);
  or2  I150_014(w_150_016, w_071_017, w_150_015);
  or2  I150_015(w_150_008, w_096_009, w_150_016);
  and2 I151_148(w_151_148, w_133_012, w_103_013);
  nand2 I152_057(w_152_057, w_059_134, w_027_032);
  and2 I153_000(w_153_000, w_061_003, w_142_002);
  and2 I153_001(w_153_001, w_035_073, w_094_084);
  and2 I154_034(w_154_034, w_053_005, w_031_105);
  not1 I154_098(w_154_098, w_089_033);
  nand2 I156_018(w_156_018, w_003_017, w_027_051);
  nand2 I156_023(w_156_023, w_153_000, w_121_013);
  not1 I157_014(w_157_014, w_030_063);
  nand2 I157_024(w_157_024, w_023_118, w_138_148);
  not1 I158_056(w_158_056, w_122_059);
  not1 I159_092(w_159_092, w_066_011);
  nand2 I159_173(w_159_173, w_071_007, w_103_127);
  not1 I161_002(w_161_002, w_144_036);
  or2  I161_061(w_161_061, w_036_008, w_159_173);
  not1 I161_079(w_161_079, w_001_011);
  nand2 I165_060(w_165_060, w_042_015, w_113_001);
  nand2 I166_003(w_166_003, w_068_018, w_046_090);
  or2  I166_035(w_166_035, w_159_092, w_147_061);
  or2  I167_046(w_167_046, w_013_031, w_069_155);
  not1 I167_076(w_167_076, w_138_132);
  or2  I167_097(w_167_097, w_080_008, w_050_049);
  and2 I168_000(w_168_000, w_023_044, w_006_018);
  and2 I168_002(w_168_002, w_039_004, w_026_012);
  or2  I168_004(w_168_004, w_154_034, w_035_083);
  not1 I168_006(w_168_006, w_049_129);
  or2  I169_001(w_169_001, w_158_056, w_091_100);
  or2  I169_020(w_169_020, w_089_039, w_131_037);
  or2  I169_025(w_169_025, w_002_050, w_002_000);
  and2 I169_039(w_169_039, w_118_030, w_153_001);
  and2 I169_041(w_169_041, w_128_022, w_112_061);
  or2  I170_099(w_170_099, w_133_143, w_166_035);
  and2 I170_134(w_170_134, w_080_032, w_102_135);
  or2  I171_021(w_171_021, w_043_062, w_170_134);
  nand2 I172_091(w_172_091, w_015_033, w_080_036);
  and2 I173_006(w_173_006, w_030_061, w_165_060);
  or2  I176_076(w_176_076, w_171_021, w_172_091);
  or2  I176_165(w_176_167, w_176_166, w_050_074);
  or2  I176_166(w_176_168, w_018_082, w_176_167);
  and2 I176_167(w_176_169, w_069_133, w_176_168);
  not1 I176_168(w_176_170, w_176_169);
  or2  I176_169(w_176_171, w_143_001, w_176_170);
  and2 I176_170(w_176_172, w_086_035, w_176_171);
  not1 I176_171(w_176_166, w_176_172);
  or2  I178_045(w_178_045, w_130_117, w_124_047);
  or2  I179_001(w_179_001, w_133_038, w_123_000);
  and2 I180_034(w_180_034, w_167_097, w_102_079);
  not1 I180_037(w_180_037, w_097_020);
  or2  I181_024(w_181_024, w_100_019, w_047_012);
  or2  I183_089(w_183_089, w_147_080, w_134_020);
  nand2 I184_112(w_184_112, w_119_006, w_146_126);
  not1 I188_021(w_188_021, w_014_125);
  or2  I188_046(w_188_046, w_096_016, w_056_103);
  nand2 I188_057(w_188_057, w_014_100, w_112_089);
  not1 I190_031(w_190_031, w_139_031);
  nand2 I192_011(w_192_011, w_063_068, w_167_046);
  nand2 I194_054(w_194_054, w_035_076, w_055_015);
  or2  I195_004(w_195_004, w_031_002, w_161_079);
  and2 I196_042(w_196_042, w_059_097, w_107_019);
  and2 I197_015(w_197_015, w_188_057, w_062_060);
  nand2 I200_000(w_200_000, w_025_128, w_156_023);
  nand2 I200_001(w_200_001, w_002_059, w_161_061);
  or2  I200_002(w_200_002, w_141_004, w_144_052);
  or2  I200_003(w_200_003, w_050_069, w_031_103);
  or2  I200_004(w_200_004, w_063_010, w_056_058);
  not1 I200_005(w_200_005, w_142_006);
  nand2 I200_006(w_200_006, w_003_006, w_094_080);
  not1 I200_007(w_200_007, w_003_027);
  or2  I200_008(w_200_008, w_005_017, w_170_099);
  not1 I200_009(w_200_009, w_064_165);
  nand2 I200_010(w_200_010, w_068_046, w_157_024);
  or2  I200_011(w_200_011, w_012_107, w_044_000);
  and2 I200_012(w_200_012, w_038_013, w_010_034);
  and2 I200_013(w_200_013, w_013_024, w_054_005);
  not1 I200_014(w_200_014, w_057_026);
  and2 I200_015(w_200_015, w_015_058, w_126_002);
  and2 I200_016(w_200_016, w_190_031, w_059_058);
  not1 I200_017(w_200_017, w_168_000);
  nand2 I200_018(w_200_018, w_180_037, w_104_119);
  and2 I200_019(w_200_019, w_094_084, w_058_028);
  and2 I200_020(w_200_020, w_023_053, w_002_038);
  nand2 I200_021(w_200_021, w_060_061, w_051_027);
  not1 I200_022(w_200_022, w_178_045);
  not1 I200_023(w_200_023, w_168_004);
  or2  I200_024(w_200_024, w_179_001, w_013_027);
  not1 I200_025(w_200_025, w_145_004);
  not1 I200_026(w_200_026, w_064_079);
  and2 I200_027(w_200_027, w_100_002, w_144_096);
  and2 I200_028(w_200_028, w_149_015, w_080_001);
  nand2 I200_029(w_200_029, w_021_048, w_090_015);
  not1 I200_030(w_200_030, w_183_089);
  nand2 I200_031(w_200_031, w_011_134, w_078_070);
  nand2 I200_032(w_200_032, w_129_036, w_044_161);
  not1 I200_033(w_200_033, w_061_035);
  not1 I200_034(w_200_034, w_161_002);
  not1 I200_035(w_200_035, w_058_089);
  and2 I200_036(w_200_036, w_109_075, w_169_020);
  and2 I200_037(w_200_037, w_169_025, w_151_148);
  or2  I200_038(w_200_038, w_040_047, w_008_005);
  or2  I200_039(w_200_039, w_078_015, w_054_004);
  or2  I200_040(w_200_040, w_167_076, w_034_017);
  not1 I200_041(w_200_041, w_196_042);
  or2  I200_042(w_200_042, w_006_072, w_197_015);
  nand2 I200_043(w_200_043, w_166_003, w_111_011);
  or2  I200_044(w_200_044, w_014_035, w_194_054);
  not1 I200_045(w_200_045, w_002_002);
  nand2 I200_046(w_200_046, w_081_017, w_014_007);
  nand2 I200_047(w_200_047, w_181_024, w_117_000);
  not1 I200_048(w_200_048, w_065_064);
  nand2 I200_049(w_200_049, w_071_076, w_000_138);
  nand2 I200_050(w_200_050, w_118_025, w_003_006);
  not1 I200_051(w_200_051, w_169_041);
  and2 I200_052(w_200_052, w_176_076, w_123_108);
  nand2 I200_053(w_200_053, w_156_018, w_001_017);
  or2  I200_054(w_200_054, w_135_079, w_122_028);
  not1 I200_055(w_200_055, w_188_021);
  or2  I200_056(w_200_056, w_011_051, w_014_102);
  nand2 I200_057(w_200_057, w_084_079, w_038_004);
  not1 I200_058(w_200_058, w_008_036);
  not1 I200_059(w_200_059, w_184_112);
  or2  I200_060(w_200_060, w_044_099, w_157_014);
  or2  I200_061(w_200_061, w_013_067, w_140_044);
  not1 I200_062(w_200_062, w_168_006);
  not1 I200_063(w_200_063, w_036_012);
  or2  I200_064(w_200_064, w_180_034, w_147_016);
  not1 I200_065(w_200_065, w_027_054);
  or2  I200_066(w_200_066, w_033_014, w_149_019);
  not1 I200_067(w_200_067, w_013_017);
  nand2 I200_068(w_200_068, w_064_070, w_009_117);
  nand2 I200_069(w_200_069, w_029_009, w_080_024);
  not1 I200_070(w_200_070, w_134_007);
  not1 I200_071(w_200_071, w_154_098);
  nand2 I200_072(w_200_072, w_188_046, w_115_011);
  or2  I200_073(w_200_073, w_169_039, w_058_031);
  or2  I200_074(w_200_074, w_169_001, w_038_006);
  or2  I200_075(w_200_075, w_054_003, w_195_004);
  and2 I200_076(w_200_076, w_024_001, w_020_011);
  nand2 I200_077(w_200_077, w_107_152, w_030_061);
  not1 I200_078(w_200_078, w_129_002);
  and2 I200_079(w_200_079, w_044_013, w_073_025);
  or2  I200_080(w_200_080, w_131_101, w_114_053);
  and2 I200_081(w_200_081, w_152_057, w_173_006);
  and2 I200_082(w_200_082, w_168_002, w_029_004);
  and2 I200_083(w_200_083, w_001_005, w_079_009);
  nand2 I200_084(w_200_084, w_109_122, w_046_056);
  and2 I200_085(w_200_085, w_094_086, w_089_020);
  and2 I200_086(w_200_086, w_130_051, w_005_044);
  and2 I200_087(w_200_087, w_145_013, w_192_011);

  initial begin
    $get_module_info();
  end
endmodule

// ****** Combined Logic Module Defination ******

// ****** TestBench Module Defination ******

/*
module tb();
  wire  w_000_000, w_000_001, w_000_002, w_000_003, w_000_004, w_000_005, w_000_006, w_000_007, w_000_008, w_000_009, w_000_010, w_000_011, w_000_012, w_000_013, w_000_014, w_000_015, w_000_016, w_000_017, w_000_018, w_000_019, w_000_020, w_000_021, w_000_022, w_000_023, w_000_024, w_000_025, w_000_026, w_000_027, w_000_028, w_000_029, w_000_030, w_000_031, w_000_032, w_000_033, w_000_034, w_000_035, w_000_036, w_000_037, w_000_038, w_000_039, w_000_040, w_000_041, w_000_042, w_000_043, w_000_044, w_000_045, w_000_046, w_000_047, w_000_048, w_000_049, w_000_050, w_000_051, w_000_052, w_000_053, w_000_054, w_000_055, w_000_056, w_000_057, w_000_058, w_000_059, w_000_060, w_000_061, w_000_062, w_000_063, w_000_064, w_000_065, w_000_066, w_000_067, w_000_068, w_000_069, w_000_070, w_000_071, w_000_072, w_000_073, w_000_074, w_000_075, w_000_076, w_000_077, w_000_078, w_000_079, w_000_080, w_000_081, w_000_082, w_000_083, w_000_084, w_000_085, w_000_086, w_000_087, w_000_088, w_000_089, w_000_090, w_000_091, w_000_092, w_000_093, w_000_094, w_000_095, w_000_096, w_000_097, w_000_098, w_000_099, w_000_100, w_000_102, w_000_103, w_000_104, w_000_105, w_000_106, w_000_109, w_000_110, w_000_111, w_000_112, w_000_113, w_000_114, w_000_115, w_000_116, w_000_117, w_000_119, w_000_120, w_000_121, w_000_122, w_000_124, w_000_125, w_000_126, w_000_127, w_000_128, w_000_129, w_000_130, w_000_131, w_000_132, w_000_135, w_000_136, w_000_137, w_000_138, w_000_139, w_000_140, w_000_142, w_000_143, w_000_144, w_000_145, w_000_148, w_000_150, w_000_151, w_000_152, w_000_153, w_000_154, w_000_155, w_000_157, w_000_159, w_000_160, w_000_161, w_000_162, w_000_165, w_000_166, w_000_168, w_000_169, w_000_170, w_000_172, w_000_173, w_000_175, w_000_177, w_000_178, w_000_180, w_000_186, w_000_189, w_200_000, w_200_001, w_200_002, w_200_003, w_200_004, w_200_005, w_200_006, w_200_007, w_200_008, w_200_009, w_200_010, w_200_011, w_200_012, w_200_013, w_200_014, w_200_015, w_200_016, w_200_017, w_200_018, w_200_019, w_200_020, w_200_021, w_200_022, w_200_023, w_200_024, w_200_025, w_200_026, w_200_027, w_200_028, w_200_029, w_200_030, w_200_031, w_200_032, w_200_033, w_200_034, w_200_035, w_200_036, w_200_037, w_200_038, w_200_039, w_200_040, w_200_041, w_200_042, w_200_043, w_200_044, w_200_045, w_200_046, w_200_047, w_200_048, w_200_049, w_200_050, w_200_051, w_200_052, w_200_053, w_200_054, w_200_055, w_200_056, w_200_057, w_200_058, w_200_059, w_200_060, w_200_061, w_200_062, w_200_063, w_200_064, w_200_065, w_200_066, w_200_067, w_200_068, w_200_069, w_200_070, w_200_071, w_200_072, w_200_073, w_200_074, w_200_075, w_200_076, w_200_077, w_200_078, w_200_079, w_200_080, w_200_081, w_200_082, w_200_083, w_200_084, w_200_085, w_200_086, w_200_087 ;
  combLogic I0(  w_000_000, w_000_001, w_000_002, w_000_003, w_000_004, w_000_005, w_000_006, w_000_007, w_000_008, w_000_009, w_000_010, w_000_011, w_000_012, w_000_013, w_000_014, w_000_015, w_000_016, w_000_017, w_000_018, w_000_019, w_000_020, w_000_021, w_000_022, w_000_023, w_000_024, w_000_025, w_000_026, w_000_027, w_000_028, w_000_029, w_000_030, w_000_031, w_000_032, w_000_033, w_000_034, w_000_035, w_000_036, w_000_037, w_000_038, w_000_039, w_000_040, w_000_041, w_000_042, w_000_043, w_000_044, w_000_045, w_000_046, w_000_047, w_000_048, w_000_049, w_000_050, w_000_051, w_000_052, w_000_053, w_000_054, w_000_055, w_000_056, w_000_057, w_000_058, w_000_059, w_000_060, w_000_061, w_000_062, w_000_063, w_000_064, w_000_065, w_000_066, w_000_067, w_000_068, w_000_069, w_000_070, w_000_071, w_000_072, w_000_073, w_000_074, w_000_075, w_000_076, w_000_077, w_000_078, w_000_079, w_000_080, w_000_081, w_000_082, w_000_083, w_000_084, w_000_085, w_000_086, w_000_087, w_000_088, w_000_089, w_000_090, w_000_091, w_000_092, w_000_093, w_000_094, w_000_095, w_000_096, w_000_097, w_000_098, w_000_099, w_000_100, w_000_102, w_000_103, w_000_104, w_000_105, w_000_106, w_000_109, w_000_110, w_000_111, w_000_112, w_000_113, w_000_114, w_000_115, w_000_116, w_000_117, w_000_119, w_000_120, w_000_121, w_000_122, w_000_124, w_000_125, w_000_126, w_000_127, w_000_128, w_000_129, w_000_130, w_000_131, w_000_132, w_000_135, w_000_136, w_000_137, w_000_138, w_000_139, w_000_140, w_000_142, w_000_143, w_000_144, w_000_145, w_000_148, w_000_150, w_000_151, w_000_152, w_000_153, w_000_154, w_000_155, w_000_157, w_000_159, w_000_160, w_000_161, w_000_162, w_000_165, w_000_166, w_000_168, w_000_169, w_000_170, w_000_172, w_000_173, w_000_175, w_000_177, w_000_178, w_000_180, w_000_186, w_000_189, w_200_000, w_200_001, w_200_002, w_200_003, w_200_004, w_200_005, w_200_006, w_200_007, w_200_008, w_200_009, w_200_010, w_200_011, w_200_012, w_200_013, w_200_014, w_200_015, w_200_016, w_200_017, w_200_018, w_200_019, w_200_020, w_200_021, w_200_022, w_200_023, w_200_024, w_200_025, w_200_026, w_200_027, w_200_028, w_200_029, w_200_030, w_200_031, w_200_032, w_200_033, w_200_034, w_200_035, w_200_036, w_200_037, w_200_038, w_200_039, w_200_040, w_200_041, w_200_042, w_200_043, w_200_044, w_200_045, w_200_046, w_200_047, w_200_048, w_200_049, w_200_050, w_200_051, w_200_052, w_200_053, w_200_054, w_200_055, w_200_056, w_200_057, w_200_058, w_200_059, w_200_060, w_200_061, w_200_062, w_200_063, w_200_064, w_200_065, w_200_066, w_200_067, w_200_068, w_200_069, w_200_070, w_200_071, w_200_072, w_200_073, w_200_074, w_200_075, w_200_076, w_200_077, w_200_078, w_200_079, w_200_080, w_200_081, w_200_082, w_200_083, w_200_084, w_200_085, w_200_086, w_200_087  );

  reg r0, r1, r2, r3, r4, r5, r6, r7, r8, r9, r10, r11, r12, r13, r14, r15, r16, r17, r18, r19, r20, r21, r22, r23, r24, r25, r26, r27, r28, r29, r30, r31, r32, r33, r34, r35, r36, r37, r38, r39, r40, r41, r42, r43, r44, r45, r46, r47, r48, r49, r50, r51, r52, r53, r54, r55, r56, r57, r58, r59, r60, r61, r62, r63, r64, r65, r66, r67, r68, r69, r70, r71, r72, r73, r74, r75, r76, r77, r78, r79, r80, r81, r82, r83, r84, r85, r86, r87, r88, r89, r90, r91, r92, r93, r94, r95, r96, r97, r98, r99, r100, r101, r102, r103, r104, r105, r106, r107, r108, r109, r110, r111, r112, r113, r114, r115, r116, r117, r118, r119, r120, r121, r122, r123, r124, r125, r126, r127, r128, r129, r130, r131, r132, r133, r134, r135, r136, r137, r138, r139, r140, r141, r142, r143, r144, r145, r146, r147, r148, r149, r150, r151, r152, r153, r154, r155, r156, r157, r158, r159, r160, r161, r162, r163, r164, r165, r166, r167, r168, r169, r170, r171, r172, r173, r174, r175, r176, r177, r178, r179, r180, r181, r182, r183, r184, r185, r186, r187, r188, r189, r190, r191, r192, r193, r194, r195, r196, r197, r198, rEnd; 

  assign w_000_000 = r0;
  assign w_000_001 = r1;
  assign w_000_002 = r2;
  assign w_000_003 = r3;
  assign w_000_004 = r4;
  assign w_000_005 = r5;
  assign w_000_006 = r6;
  assign w_000_007 = r7;
  assign w_000_008 = r8;
  assign w_000_009 = r9;
  assign w_000_010 = r10;
  assign w_000_011 = r11;
  assign w_000_012 = r12;
  assign w_000_013 = r13;
  assign w_000_014 = r14;
  assign w_000_015 = r15;
  assign w_000_016 = r16;
  assign w_000_017 = r17;
  assign w_000_018 = r18;
  assign w_000_019 = r19;
  assign w_000_020 = r20;
  assign w_000_021 = r21;
  assign w_000_022 = r22;
  assign w_000_023 = r23;
  assign w_000_024 = r24;
  assign w_000_025 = r25;
  assign w_000_026 = r26;
  assign w_000_027 = r27;
  assign w_000_028 = r28;
  assign w_000_029 = r29;
  assign w_000_030 = r30;
  assign w_000_031 = r31;
  assign w_000_032 = r32;
  assign w_000_033 = r33;
  assign w_000_034 = r34;
  assign w_000_035 = r35;
  assign w_000_036 = r36;
  assign w_000_037 = r37;
  assign w_000_038 = r38;
  assign w_000_039 = r39;
  assign w_000_040 = r40;
  assign w_000_041 = r41;
  assign w_000_042 = r42;
  assign w_000_043 = r43;
  assign w_000_044 = r44;
  assign w_000_045 = r45;
  assign w_000_046 = r46;
  assign w_000_047 = r47;
  assign w_000_048 = r48;
  assign w_000_049 = r49;
  assign w_000_050 = r50;
  assign w_000_051 = r51;
  assign w_000_052 = r52;
  assign w_000_053 = r53;
  assign w_000_054 = r54;
  assign w_000_055 = r55;
  assign w_000_056 = r56;
  assign w_000_057 = r57;
  assign w_000_058 = r58;
  assign w_000_059 = r59;
  assign w_000_060 = r60;
  assign w_000_061 = r61;
  assign w_000_062 = r62;
  assign w_000_063 = r63;
  assign w_000_064 = r64;
  assign w_000_065 = r65;
  assign w_000_066 = r66;
  assign w_000_067 = r67;
  assign w_000_068 = r68;
  assign w_000_069 = r69;
  assign w_000_070 = r70;
  assign w_000_071 = r71;
  assign w_000_072 = r72;
  assign w_000_073 = r73;
  assign w_000_074 = r74;
  assign w_000_075 = r75;
  assign w_000_076 = r76;
  assign w_000_077 = r77;
  assign w_000_078 = r78;
  assign w_000_079 = r79;
  assign w_000_080 = r80;
  assign w_000_081 = r81;
  assign w_000_082 = r82;
  assign w_000_083 = r83;
  assign w_000_084 = r84;
  assign w_000_085 = r85;
  assign w_000_086 = r86;
  assign w_000_087 = r87;
  assign w_000_088 = r88;
  assign w_000_089 = r89;
  assign w_000_090 = r90;
  assign w_000_091 = r91;
  assign w_000_092 = r92;
  assign w_000_093 = r93;
  assign w_000_094 = r94;
  assign w_000_095 = r95;
  assign w_000_096 = r96;
  assign w_000_097 = r97;
  assign w_000_098 = r98;
  assign w_000_099 = r99;
  assign w_000_100 = r100;
  assign w_000_101 = r101;
  assign w_000_102 = r102;
  assign w_000_103 = r103;
  assign w_000_104 = r104;
  assign w_000_105 = r105;
  assign w_000_106 = r106;
  assign w_000_107 = r107;
  assign w_000_108 = r108;
  assign w_000_109 = r109;
  assign w_000_110 = r110;
  assign w_000_111 = r111;
  assign w_000_112 = r112;
  assign w_000_113 = r113;
  assign w_000_114 = r114;
  assign w_000_115 = r115;
  assign w_000_116 = r116;
  assign w_000_117 = r117;
  assign w_000_118 = r118;
  assign w_000_119 = r119;
  assign w_000_120 = r120;
  assign w_000_121 = r121;
  assign w_000_122 = r122;
  assign w_000_123 = r123;
  assign w_000_124 = r124;
  assign w_000_125 = r125;
  assign w_000_126 = r126;
  assign w_000_127 = r127;
  assign w_000_128 = r128;
  assign w_000_129 = r129;
  assign w_000_130 = r130;
  assign w_000_131 = r131;
  assign w_000_132 = r132;
  assign w_000_133 = r133;
  assign w_000_134 = r134;
  assign w_000_135 = r135;
  assign w_000_136 = r136;
  assign w_000_137 = r137;
  assign w_000_138 = r138;
  assign w_000_139 = r139;
  assign w_000_140 = r140;
  assign w_000_141 = r141;
  assign w_000_142 = r142;
  assign w_000_143 = r143;
  assign w_000_144 = r144;
  assign w_000_145 = r145;
  assign w_000_146 = r146;
  assign w_000_147 = r147;
  assign w_000_148 = r148;
  assign w_000_149 = r149;
  assign w_000_150 = r150;
  assign w_000_151 = r151;
  assign w_000_152 = r152;
  assign w_000_153 = r153;
  assign w_000_154 = r154;
  assign w_000_155 = r155;
  assign w_000_156 = r156;
  assign w_000_157 = r157;
  assign w_000_158 = r158;
  assign w_000_159 = r159;
  assign w_000_160 = r160;
  assign w_000_161 = r161;
  assign w_000_162 = r162;
  assign w_000_163 = r163;
  assign w_000_164 = r164;
  assign w_000_165 = r165;
  assign w_000_166 = r166;
  assign w_000_167 = r167;
  assign w_000_168 = r168;
  assign w_000_169 = r169;
  assign w_000_170 = r170;
  assign w_000_171 = r171;
  assign w_000_172 = r172;
  assign w_000_173 = r173;
  assign w_000_174 = r174;
  assign w_000_175 = r175;
  assign w_000_176 = r176;
  assign w_000_177 = r177;
  assign w_000_178 = r178;
  assign w_000_179 = r179;
  assign w_000_180 = r180;
  assign w_000_181 = r181;
  assign w_000_182 = r182;
  assign w_000_183 = r183;
  assign w_000_184 = r184;
  assign w_000_185 = r185;
  assign w_000_186 = r186;
  assign w_000_187 = r187;
  assign w_000_188 = r188;
  assign w_000_189 = r189;
  assign w_000_190 = r190;
  assign w_000_191 = r191;
  assign w_000_192 = r192;
  assign w_000_193 = r193;
  assign w_000_194 = r194;
  assign w_000_195 = r195;
  assign w_000_196 = r196;
  assign w_000_197 = r197;
  assign w_000_198 = r198;

  initial begin 
    r0 = 1'b0; 
    r1 = 1'b0; 
    r2 = 1'b0; 
    r3 = 1'b0; 
    r4 = 1'b0; 
    r5 = 1'b0; 
    r6 = 1'b0; 
    r7 = 1'b0; 
    r8 = 1'b0; 
    r9 = 1'b0; 
    r10 = 1'b0; 
    r11 = 1'b0; 
    r12 = 1'b0; 
    r13 = 1'b0; 
    r14 = 1'b0; 
    r15 = 1'b0; 
    r16 = 1'b0; 
    r17 = 1'b0; 
    r18 = 1'b0; 
    r19 = 1'b0; 
    r20 = 1'b0; 
    r21 = 1'b0; 
    r22 = 1'b0; 
    r23 = 1'b0; 
    r24 = 1'b0; 
    r25 = 1'b0; 
    r26 = 1'b0; 
    r27 = 1'b0; 
    r28 = 1'b0; 
    r29 = 1'b0; 
    r30 = 1'b0; 
    r31 = 1'b0; 
    r32 = 1'b0; 
    r33 = 1'b0; 
    r34 = 1'b0; 
    r35 = 1'b0; 
    r36 = 1'b0; 
    r37 = 1'b0; 
    r38 = 1'b0; 
    r39 = 1'b0; 
    r40 = 1'b0; 
    r41 = 1'b0; 
    r42 = 1'b0; 
    r43 = 1'b0; 
    r44 = 1'b0; 
    r45 = 1'b0; 
    r46 = 1'b0; 
    r47 = 1'b0; 
    r48 = 1'b0; 
    r49 = 1'b0; 
    r50 = 1'b0; 
    r51 = 1'b0; 
    r52 = 1'b0; 
    r53 = 1'b0; 
    r54 = 1'b0; 
    r55 = 1'b0; 
    r56 = 1'b0; 
    r57 = 1'b0; 
    r58 = 1'b0; 
    r59 = 1'b0; 
    r60 = 1'b0; 
    r61 = 1'b0; 
    r62 = 1'b0; 
    r63 = 1'b0; 
    r64 = 1'b0; 
    r65 = 1'b0; 
    r66 = 1'b0; 
    r67 = 1'b0; 
    r68 = 1'b0; 
    r69 = 1'b0; 
    r70 = 1'b0; 
    r71 = 1'b0; 
    r72 = 1'b0; 
    r73 = 1'b0; 
    r74 = 1'b0; 
    r75 = 1'b0; 
    r76 = 1'b0; 
    r77 = 1'b0; 
    r78 = 1'b0; 
    r79 = 1'b0; 
    r80 = 1'b0; 
    r81 = 1'b0; 
    r82 = 1'b0; 
    r83 = 1'b0; 
    r84 = 1'b0; 
    r85 = 1'b0; 
    r86 = 1'b0; 
    r87 = 1'b0; 
    r88 = 1'b0; 
    r89 = 1'b0; 
    r90 = 1'b0; 
    r91 = 1'b0; 
    r92 = 1'b0; 
    r93 = 1'b0; 
    r94 = 1'b0; 
    r95 = 1'b0; 
    r96 = 1'b0; 
    r97 = 1'b0; 
    r98 = 1'b0; 
    r99 = 1'b0; 
    r100 = 1'b0; 
    r101 = 1'b0; 
    r102 = 1'b0; 
    r103 = 1'b0; 
    r104 = 1'b0; 
    r105 = 1'b0; 
    r106 = 1'b0; 
    r107 = 1'b0; 
    r108 = 1'b0; 
    r109 = 1'b0; 
    r110 = 1'b0; 
    r111 = 1'b0; 
    r112 = 1'b0; 
    r113 = 1'b0; 
    r114 = 1'b0; 
    r115 = 1'b0; 
    r116 = 1'b0; 
    r117 = 1'b0; 
    r118 = 1'b0; 
    r119 = 1'b0; 
    r120 = 1'b0; 
    r121 = 1'b0; 
    r122 = 1'b0; 
    r123 = 1'b0; 
    r124 = 1'b0; 
    r125 = 1'b0; 
    r126 = 1'b0; 
    r127 = 1'b0; 
    r128 = 1'b0; 
    r129 = 1'b0; 
    r130 = 1'b0; 
    r131 = 1'b0; 
    r132 = 1'b0; 
    r133 = 1'b0; 
    r134 = 1'b0; 
    r135 = 1'b0; 
    r136 = 1'b0; 
    r137 = 1'b0; 
    r138 = 1'b0; 
    r139 = 1'b0; 
    r140 = 1'b0; 
    r141 = 1'b0; 
    r142 = 1'b0; 
    r143 = 1'b0; 
    r144 = 1'b0; 
    r145 = 1'b0; 
    r146 = 1'b0; 
    r147 = 1'b0; 
    r148 = 1'b0; 
    r149 = 1'b0; 
    r150 = 1'b0; 
    r151 = 1'b0; 
    r152 = 1'b0; 
    r153 = 1'b0; 
    r154 = 1'b0; 
    r155 = 1'b0; 
    r156 = 1'b0; 
    r157 = 1'b0; 
    r158 = 1'b0; 
    r159 = 1'b0; 
    r160 = 1'b0; 
    r161 = 1'b0; 
    r162 = 1'b0; 
    r163 = 1'b0; 
    r164 = 1'b0; 
    r165 = 1'b0; 
    r166 = 1'b0; 
    r167 = 1'b0; 
    r168 = 1'b0; 
    r169 = 1'b0; 
    r170 = 1'b0; 
    r171 = 1'b0; 
    r172 = 1'b0; 
    r173 = 1'b0; 
    r174 = 1'b0; 
    r175 = 1'b0; 
    r176 = 1'b0; 
    r177 = 1'b0; 
    r178 = 1'b0; 
    r179 = 1'b0; 
    r180 = 1'b0; 
    r181 = 1'b0; 
    r182 = 1'b0; 
    r183 = 1'b0; 
    r184 = 1'b0; 
    r185 = 1'b0; 
    r186 = 1'b0; 
    r187 = 1'b0; 
    r188 = 1'b0; 
    r189 = 1'b0; 
    r190 = 1'b0; 
    r191 = 1'b0; 
    r192 = 1'b0; 
    r193 = 1'b0; 
    r194 = 1'b0; 
    r195 = 1'b0; 
    r196 = 1'b0; 
    r197 = 1'b0; 
    r198 = 1'b0; 
    $monitor("%t %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b  ", $time, w_000_000, w_000_001, w_000_002, w_000_003, w_000_004, w_000_005, w_000_006, w_000_007, w_000_008, w_000_009, w_000_010, w_000_011, w_000_012, w_000_013, w_000_014, w_000_015, w_000_016, w_000_017, w_000_018, w_000_019, w_000_020, w_000_021, w_000_022, w_000_023, w_000_024, w_000_025, w_000_026, w_000_027, w_000_028, w_000_029, w_000_030, w_000_031, w_000_032, w_000_033, w_000_034, w_000_035, w_000_036, w_000_037, w_000_038, w_000_039, w_000_040, w_000_041, w_000_042, w_000_043, w_000_044, w_000_045, w_000_046, w_000_047, w_000_048, w_000_049, w_000_050, w_000_051, w_000_052, w_000_053, w_000_054, w_000_055, w_000_056, w_000_057, w_000_058, w_000_059, w_000_060, w_000_061, w_000_062, w_000_063, w_000_064, w_000_065, w_000_066, w_000_067, w_000_068, w_000_069, w_000_070, w_000_071, w_000_072, w_000_073, w_000_074, w_000_075, w_000_076, w_000_077, w_000_078, w_000_079, w_000_080, w_000_081, w_000_082, w_000_083, w_000_084, w_000_085, w_000_086, w_000_087, w_000_088, w_000_089, w_000_090, w_000_091, w_000_092, w_000_093, w_000_094, w_000_095, w_000_096, w_000_097, w_000_098, w_000_099, w_000_100, w_000_101, w_000_102, w_000_103, w_000_104, w_000_105, w_000_106, w_000_107, w_000_108, w_000_109, w_000_110, w_000_111, w_000_112, w_000_113, w_000_114, w_000_115, w_000_116, w_000_117, w_000_118, w_000_119, w_000_120, w_000_121, w_000_122, w_000_123, w_000_124, w_000_125, w_000_126, w_000_127, w_000_128, w_000_129, w_000_130, w_000_131, w_000_132, w_000_133, w_000_134, w_000_135, w_000_136, w_000_137, w_000_138, w_000_139, w_000_140, w_000_141, w_000_142, w_000_143, w_000_144, w_000_145, w_000_146, w_000_147, w_000_148, w_000_149, w_000_150, w_000_151, w_000_152, w_000_153, w_000_154, w_000_155, w_000_156, w_000_157, w_000_158, w_000_159, w_000_160, w_000_161, w_000_162, w_000_163, w_000_164, w_000_165, w_000_166, w_000_167, w_000_168, w_000_169, w_000_170, w_000_171, w_000_172, w_000_173, w_000_174, w_000_175, w_000_176, w_000_177, w_000_178, w_000_179, w_000_180, w_000_181, w_000_182, w_000_183, w_000_184, w_000_185, w_000_186, w_000_187, w_000_188, w_000_189, w_000_190, w_000_191, w_000_192, w_000_193, w_000_194, w_000_195, w_000_196, w_000_197, w_000_198, w_200_000, w_200_001, w_200_002, w_200_003, w_200_004, w_200_005, w_200_006, w_200_007, w_200_008, w_200_009, w_200_010, w_200_011, w_200_012, w_200_013, w_200_014, w_200_015, w_200_016, w_200_017, w_200_018, w_200_019, w_200_020, w_200_021, w_200_022, w_200_023, w_200_024, w_200_025, w_200_026, w_200_027, w_200_028, w_200_029, w_200_030, w_200_031, w_200_032, w_200_033, w_200_034, w_200_035, w_200_036, w_200_037, w_200_038, w_200_039, w_200_040, w_200_041, w_200_042, w_200_043, w_200_044, w_200_045, w_200_046, w_200_047, w_200_048, w_200_049, w_200_050, w_200_051, w_200_052, w_200_053, w_200_054, w_200_055, w_200_056, w_200_057, w_200_058, w_200_059, w_200_060, w_200_061, w_200_062, w_200_063, w_200_064, w_200_065, w_200_066, w_200_067, w_200_068, w_200_069, w_200_070, w_200_071, w_200_072, w_200_073, w_200_074, w_200_075, w_200_076, w_200_077, w_200_078, w_200_079, w_200_080, w_200_081, w_200_082, w_200_083, w_200_084, w_200_085, w_200_086, w_200_087);
    #100;
    $finish;
  end
  always #1 r0 = ~r0;
  always #2 r1 = ~r1;
  always #4 r2 = ~r2;
  always #8 r3 = ~r3;
  always #16 r4 = ~r4;
  always #32 r5 = ~r5;
  always #64 r6 = ~r6;
  always #128 r7 = ~r7;
  always #256 r8 = ~r8;
  always #512 r9 = ~r9;
  always #1024 r10 = ~r10;
  always #2048 r11 = ~r11;
  always #4096 r12 = ~r12;
  always #8192 r13 = ~r13;
  always #16384 r14 = ~r14;
  always #32768 r15 = ~r15;
  always #65536 r16 = ~r16;
  always #131072 r17 = ~r17;
  always #262144 r18 = ~r18;
  always #524288 r19 = ~r19;
  always #1048576 r20 = ~r20;
  always #2097152 r21 = ~r21;
  always #4194304 r22 = ~r22;
  always #8388608 r23 = ~r23;
  always #16777216 r24 = ~r24;
  always #33554432 r25 = ~r25;
  always #67108864 r26 = ~r26;
  always #134217728 r27 = ~r27;
  always #268435456 r28 = ~r28;
  always #536870912 r29 = ~r29;
  always #1073741824 r30 = ~r30;
  always #2147483648 r31 = ~r31;
  always #4294967296 r32 = ~r32;
  always #8589934592 r33 = ~r33;
  always #17179869184 r34 = ~r34;
  always #34359738368 r35 = ~r35;
  always #68719476736 r36 = ~r36;
  always #137438953472 r37 = ~r37;
  always #274877906944 r38 = ~r38;
  always #549755813888 r39 = ~r39;
  always #1099511627776 r40 = ~r40;
  always #2199023255552 r41 = ~r41;
  always #4398046511104 r42 = ~r42;
  always #8796093022208 r43 = ~r43;
  always #17592186044416 r44 = ~r44;
  always #35184372088832 r45 = ~r45;
  always #70368744177664 r46 = ~r46;
  always #140737488355328 r47 = ~r47;
  always #281474976710656 r48 = ~r48;
  always #562949953421312 r49 = ~r49;
  always #1125899906842624 r50 = ~r50;
  always #2251799813685248 r51 = ~r51;
  always #4503599627370496 r52 = ~r52;
  always #9007199254740992 r53 = ~r53;
  always #18014398509481984 r54 = ~r54;
  always #36028797018963968 r55 = ~r55;
  always #72057594037927936 r56 = ~r56;
  always #144115188075855872 r57 = ~r57;
  always #288230376151711744 r58 = ~r58;
  always #576460752303423488 r59 = ~r59;
  always #1152921504606846976 r60 = ~r60;
  always #2305843009213693952 r61 = ~r61;
  always #4611686018427387904 r62 = ~r62;
  always #9223372036854775808 r63 = ~r63;
  always #1 r64 = ~r64;
  always #2 r65 = ~r65;
  always #4 r66 = ~r66;
  always #8 r67 = ~r67;
  always #16 r68 = ~r68;
  always #32 r69 = ~r69;
  always #64 r70 = ~r70;
  always #128 r71 = ~r71;
  always #256 r72 = ~r72;
  always #512 r73 = ~r73;
  always #1024 r74 = ~r74;
  always #2048 r75 = ~r75;
  always #4096 r76 = ~r76;
  always #8192 r77 = ~r77;
  always #16384 r78 = ~r78;
  always #32768 r79 = ~r79;
  always #65536 r80 = ~r80;
  always #131072 r81 = ~r81;
  always #262144 r82 = ~r82;
  always #524288 r83 = ~r83;
  always #1048576 r84 = ~r84;
  always #2097152 r85 = ~r85;
  always #4194304 r86 = ~r86;
  always #8388608 r87 = ~r87;
  always #16777216 r88 = ~r88;
  always #33554432 r89 = ~r89;
  always #67108864 r90 = ~r90;
  always #134217728 r91 = ~r91;
  always #268435456 r92 = ~r92;
  always #536870912 r93 = ~r93;
  always #1073741824 r94 = ~r94;
  always #2147483648 r95 = ~r95;
  always #4294967296 r96 = ~r96;
  always #8589934592 r97 = ~r97;
  always #17179869184 r98 = ~r98;
  always #34359738368 r99 = ~r99;
  always #68719476736 r100 = ~r100;
  always #137438953472 r101 = ~r101;
  always #274877906944 r102 = ~r102;
  always #549755813888 r103 = ~r103;
  always #1099511627776 r104 = ~r104;
  always #2199023255552 r105 = ~r105;
  always #4398046511104 r106 = ~r106;
  always #8796093022208 r107 = ~r107;
  always #17592186044416 r108 = ~r108;
  always #35184372088832 r109 = ~r109;
  always #70368744177664 r110 = ~r110;
  always #140737488355328 r111 = ~r111;
  always #281474976710656 r112 = ~r112;
  always #562949953421312 r113 = ~r113;
  always #1125899906842624 r114 = ~r114;
  always #2251799813685248 r115 = ~r115;
  always #4503599627370496 r116 = ~r116;
  always #9007199254740992 r117 = ~r117;
  always #18014398509481984 r118 = ~r118;
  always #36028797018963968 r119 = ~r119;
  always #72057594037927936 r120 = ~r120;
  always #144115188075855872 r121 = ~r121;
  always #288230376151711744 r122 = ~r122;
  always #576460752303423488 r123 = ~r123;
  always #1152921504606846976 r124 = ~r124;
  always #2305843009213693952 r125 = ~r125;
  always #4611686018427387904 r126 = ~r126;
  always #9223372036854775808 r127 = ~r127;
  always #1 r128 = ~r128;
  always #2 r129 = ~r129;
  always #4 r130 = ~r130;
  always #8 r131 = ~r131;
  always #16 r132 = ~r132;
  always #32 r133 = ~r133;
  always #64 r134 = ~r134;
  always #128 r135 = ~r135;
  always #256 r136 = ~r136;
  always #512 r137 = ~r137;
  always #1024 r138 = ~r138;
  always #2048 r139 = ~r139;
  always #4096 r140 = ~r140;
  always #8192 r141 = ~r141;
  always #16384 r142 = ~r142;
  always #32768 r143 = ~r143;
  always #65536 r144 = ~r144;
  always #131072 r145 = ~r145;
  always #262144 r146 = ~r146;
  always #524288 r147 = ~r147;
  always #1048576 r148 = ~r148;
  always #2097152 r149 = ~r149;
  always #4194304 r150 = ~r150;
  always #8388608 r151 = ~r151;
  always #16777216 r152 = ~r152;
  always #33554432 r153 = ~r153;
  always #67108864 r154 = ~r154;
  always #134217728 r155 = ~r155;
  always #268435456 r156 = ~r156;
  always #536870912 r157 = ~r157;
  always #1073741824 r158 = ~r158;
  always #2147483648 r159 = ~r159;
  always #4294967296 r160 = ~r160;
  always #8589934592 r161 = ~r161;
  always #17179869184 r162 = ~r162;
  always #34359738368 r163 = ~r163;
  always #68719476736 r164 = ~r164;
  always #137438953472 r165 = ~r165;
  always #274877906944 r166 = ~r166;
  always #549755813888 r167 = ~r167;
  always #1099511627776 r168 = ~r168;
  always #2199023255552 r169 = ~r169;
  always #4398046511104 r170 = ~r170;
  always #8796093022208 r171 = ~r171;
  always #17592186044416 r172 = ~r172;
  always #35184372088832 r173 = ~r173;
  always #70368744177664 r174 = ~r174;
  always #140737488355328 r175 = ~r175;
  always #281474976710656 r176 = ~r176;
  always #562949953421312 r177 = ~r177;
  always #1125899906842624 r178 = ~r178;
  always #2251799813685248 r179 = ~r179;
  always #4503599627370496 r180 = ~r180;
  always #9007199254740992 r181 = ~r181;
  always #18014398509481984 r182 = ~r182;
  always #36028797018963968 r183 = ~r183;
  always #72057594037927936 r184 = ~r184;
  always #144115188075855872 r185 = ~r185;
  always #288230376151711744 r186 = ~r186;
  always #576460752303423488 r187 = ~r187;
  always #1152921504606846976 r188 = ~r188;
  always #2305843009213693952 r189 = ~r189;
  always #4611686018427387904 r190 = ~r190;
  always #9223372036854775808 r191 = ~r191;
  always #1 r192 = ~r192;
  always #2 r193 = ~r193;
  always #4 r194 = ~r194;
  always #8 r195 = ~r195;
  always #16 r196 = ~r196;
  always #32 r197 = ~r197;
  always #64 r198 = ~r198;
endmodule
*/
// ****** TestBench Module Defination End ******

/*
// ******* The results for this case *********
******* result_1.txt *********
1)
  Loop Signals: w_070_083, w_070_084, w_070_085, w_070_086, w_070_087, w_070_088, w_070_089, w_070_090, w_070_091, 
  Loop Gates: I070_082.port1, I070_083.port1, I070_084.port2, I070_085.port2, I070_086.port2, I070_087.port1, I070_088.port2, I070_089.port1, I070_090.port2, 

2)
  Loop Signals: w_114_100, w_114_101, w_114_102, w_114_103, 
  Loop Gates: I114_099.port1, I114_100.port2, I114_101.port1, I114_102.port1, 

3)
  Loop Signals: w_028_160, w_028_161, w_028_162, w_028_163, w_028_164, w_028_165, w_028_166, w_028_167, w_028_168, w_028_169, 
  Loop Gates: I028_159.port1, I028_160.port1, I028_161.port1, I028_162.port1, I028_163.port1, I028_164.port2, I028_165.port2, I028_166.port2, I028_167.port1, I028_168.port2, 

4)
  Loop Signals: w_114_107, w_114_108, w_114_109, w_114_110, w_114_111, w_114_112, w_114_113, w_114_114, w_114_115, 
  Loop Gates: I114_103.port1, I114_104.port1, I114_105.port1, I114_106.port1, I114_107.port1, I114_108.port2, I114_109.port1, I114_110.port1, I114_111.port1, 

5)
  Loop Signals: w_038_020, w_038_021, w_038_022, w_038_023, w_038_024, 
  Loop Gates: I038_019.port2, I038_020.port1, I038_021.port1, I038_022.port1, I038_023.port1, 

6)
  Loop Signals: w_021_156, w_021_157, w_021_158, w_021_159, w_021_160, w_021_161, w_021_162, 
  Loop Gates: I021_155.port1, I021_156.port1, I021_157.port1, I021_158.port1, I021_159.port1, I021_160.port2, I021_161.port2, 

7)
  Loop Signals: w_021_158, w_021_166, w_021_167, w_021_168, w_021_169, w_021_170, w_021_171, w_021_172, w_021_173, w_021_174, w_021_176, 
  Loop Gates: I021_156.port2, I021_162.port2, I021_163.port1, I021_164.port2, I021_165.port1, I021_166.port1, I021_167.port1, I021_168.port1, I021_169.port1, I021_170.port1, I021_171.port2, 

8)
  Loop Signals: w_144_198, w_144_199, w_144_200, w_144_201, w_144_202, w_144_203, w_144_204, 
  Loop Gates: I144_197.port2, I144_198.port1, I144_199.port1, I144_200.port1, I144_201.port1, I144_202.port1, I144_203.port1, 

9)
  Loop Signals: w_144_202, w_144_208, w_144_209, w_144_210, w_144_211, w_144_213, 
  Loop Gates: I144_200.port2, I144_204.port1, I144_205.port1, I144_206.port1, I144_207.port1, I144_208.port2, 

10)
  Loop Signals: w_132_053, w_132_054, w_132_055, w_132_056, w_132_057, w_132_058, w_132_059, w_132_060, w_132_061, w_132_062, w_132_063, 
  Loop Gates: I132_052.port2, I132_053.port1, I132_054.port2, I132_055.port1, I132_056.port1, I132_057.port2, I132_058.port2, I132_059.port1, I132_060.port1, I132_061.port2, I132_062.port1, 

11)
  Loop Signals: w_029_011, w_029_012, w_029_013, w_029_014, w_029_015, w_029_016, w_029_017, w_029_018, w_029_019, w_029_020, 
  Loop Gates: I029_011.port2, I029_012.port2, I029_013.port1, I029_014.port1, I029_015.port1, I029_016.port2, I029_017.port1, I029_018.port1, I029_019.port1, I029_020.port1, 

12)
  Loop Signals: w_006_117, w_006_118, w_006_119, w_006_120, w_006_121, 
  Loop Gates: I006_116.port2, I006_117.port2, I006_118.port2, I006_119.port2, I006_120.port1, 

13)
  Loop Signals: w_176_166, w_176_167, w_176_168, w_176_169, w_176_170, w_176_171, w_176_172, 
  Loop Gates: I176_165.port1, I176_166.port2, I176_167.port2, I176_168.port1, I176_169.port2, I176_170.port2, I176_171.port1, 

14)
  Loop Signals: w_026_092, w_026_093, w_026_094, w_026_095, 
  Loop Gates: I026_091.port2, I026_092.port1, I026_093.port2, I026_094.port2, 

15)
  Loop Signals: w_028_173, w_028_174, w_028_175, w_028_176, w_028_177, 
  Loop Gates: I028_169.port1, I028_170.port2, I028_171.port1, I028_172.port1, I028_173.port1, 

16)
  Loop Signals: w_021_178, w_021_179, w_021_180, w_021_181, w_021_182, w_021_183, 
  Loop Gates: I021_172.port1, I021_173.port1, I021_174.port2, I021_175.port1, I021_176.port2, I021_177.port1, 

17)
  Loop Signals: w_133_153, w_133_154, w_133_155, w_133_156, w_133_157, w_133_158, w_133_159, w_133_160, w_133_161, w_133_162, w_133_163, w_133_164, 
  Loop Gates: I133_153.port2, I133_154.port1, I133_155.port2, I133_156.port1, I133_157.port1, I133_158.port1, I133_159.port1, I133_160.port1, I133_161.port1, I133_162.port2, I133_163.port1, I133_164.port1, 

18)
  Loop Signals: w_039_011, w_039_012, w_039_013, w_039_014, w_039_015, w_039_016, w_039_017, w_039_018, w_039_019, w_039_020, w_039_021, 
  Loop Gates: I039_011.port1, I039_012.port1, I039_013.port1, I039_014.port1, I039_015.port1, I039_016.port1, I039_017.port1, I039_018.port2, I039_019.port1, I039_020.port1, I039_021.port1, 

19)
  Loop Signals: w_039_012, w_039_025, w_039_026, w_039_027, w_039_028, w_039_029, w_039_030, w_039_031, w_039_032, w_039_033, w_039_034, w_039_036, 
  Loop Gates: I039_011.port2, I039_022.port1, I039_023.port1, I039_024.port1, I039_025.port1, I039_026.port1, I039_027.port2, I039_028.port2, I039_029.port1, I039_030.port1, I039_031.port1, I039_032.port2, 

20)
  Loop Signals: w_150_008, w_150_009, w_150_010, w_150_011, w_150_012, w_150_013, w_150_014, w_150_015, w_150_016, 
  Loop Gates: I150_007.port1, I150_008.port1, I150_009.port2, I150_010.port1, I150_011.port1, I150_012.port1, I150_013.port1, I150_014.port2, I150_015.port2, 

******* result_2.txt *********
1)
  Loop Signals: w_070_083, w_070_084, w_070_085, w_070_086, w_070_087, w_070_088, w_070_089, w_070_090, w_070_091, 
  Loop Gates: I070_082.port1, I070_083.port1, I070_084.port2, I070_085.port2, I070_086.port2, I070_087.port1, I070_088.port2, I070_089.port1, I070_090.port2, 

2)
  Loop Signals: w_114_100, w_114_101, w_114_102, w_114_103, 
  Loop Gates: I114_099.port1, I114_100.port2, I114_101.port1, I114_102.port1, 

3)
  Loop Signals: w_038_020, w_038_021, w_038_022, w_038_023, w_038_024, 
  Loop Gates: I038_019.port2, I038_020.port1, I038_021.port1, I038_022.port1, I038_023.port1, 

4)
  Loop Signals: w_021_156, w_021_157, w_021_158, w_021_159, w_021_160, w_021_161, w_021_162, 
  Loop Gates: I021_155.port1, I021_156.port1, I021_157.port1, I021_158.port1, I021_159.port1, I021_160.port2, I021_161.port2, 

5)
  Loop Signals: w_021_158, w_021_166, w_021_167, w_021_168, w_021_169, w_021_170, w_021_171, w_021_172, w_021_173, w_021_174, w_021_176, 
  Loop Gates: I021_156.port2, I021_162.port2, I021_163.port1, I021_164.port2, I021_165.port1, I021_166.port1, I021_167.port1, I021_168.port1, I021_169.port1, I021_170.port1, I021_171.port2, 

6)
  Loop Signals: w_132_053, w_132_054, w_132_055, w_132_056, w_132_057, w_132_058, w_132_059, w_132_060, w_132_061, w_132_062, w_132_063, 
  Loop Gates: I132_052.port2, I132_053.port1, I132_054.port2, I132_055.port1, I132_056.port1, I132_057.port2, I132_058.port2, I132_059.port1, I132_060.port1, I132_061.port2, I132_062.port1, 

7)
  Loop Signals: w_006_117, w_006_118, w_006_119, w_006_120, w_006_121, 
  Loop Gates: I006_116.port2, I006_117.port2, I006_118.port2, I006_119.port2, I006_120.port1, 

8)
  Loop Signals: w_176_166, w_176_167, w_176_168, w_176_169, w_176_170, w_176_171, w_176_172, 
  Loop Gates: I176_165.port1, I176_166.port2, I176_167.port2, I176_168.port1, I176_169.port2, I176_170.port2, I176_171.port1, 

9)
  Loop Signals: w_026_092, w_026_093, w_026_094, w_026_095, 
  Loop Gates: I026_091.port2, I026_092.port1, I026_093.port2, I026_094.port2, 

10)
  Loop Signals: w_028_173, w_028_174, w_028_175, w_028_176, w_028_177, 
  Loop Gates: I028_169.port1, I028_170.port2, I028_171.port1, I028_172.port1, I028_173.port1, 

11)
  Loop Signals: w_039_011, w_039_012, w_039_013, w_039_014, w_039_015, w_039_016, w_039_017, w_039_018, w_039_019, w_039_020, w_039_021, 
  Loop Gates: I039_011.port1, I039_012.port1, I039_013.port1, I039_014.port1, I039_015.port1, I039_016.port1, I039_017.port1, I039_018.port2, I039_019.port1, I039_020.port1, I039_021.port1, 

******* result_3.txt *********
1)
  Loop Signals: w_028_160, w_028_161, w_028_162, w_028_163, w_028_164, w_028_165, w_028_166, w_028_167, w_028_168, w_028_169, 
  Loop Gates: I028_159.port1, I028_160.port1, I028_161.port1, I028_162.port1, I028_163.port1, I028_164.port2, I028_165.port2, I028_166.port2, I028_167.port1, I028_168.port2, 
  Loop Conditions: I028_159.port2=1, I028_160.port2=0, I028_162.port2=1, I028_163.port2=1, I028_164.port1=0, I028_165.port1=1, I028_166.port1=1, I028_167.port2=1, I028_168.port1=0, 
  (Signal Values: w_002_054=1, w_004_082=1, w_007_039=1, w_008_020=1, w_015_086=0, w_015_043=0, w_017_113=1, w_022_075=0, w_027_020=1, )

2)
  Loop Signals: w_114_107, w_114_108, w_114_109, w_114_110, w_114_111, w_114_112, w_114_113, w_114_114, w_114_115, 
  Loop Gates: I114_103.port1, I114_104.port1, I114_105.port1, I114_106.port1, I114_107.port1, I114_108.port2, I114_109.port1, I114_110.port1, I114_111.port1, 
  Loop Conditions: I114_103.port2=1, I114_105.port2=1, I114_107.port2=1, I114_108.port1=1, I114_109.port2=1, I114_111.port2=0, 
  (Signal Values: w_005_063=1, w_014_070=1, w_054_000=1, w_070_055=1, w_077_031=1, w_093_030=0, )

3)
  Loop Signals: w_144_198, w_144_199, w_144_200, w_144_201, w_144_202, w_144_203, w_144_204, 
  Loop Gates: I144_197.port2, I144_198.port1, I144_199.port1, I144_200.port1, I144_201.port1, I144_202.port1, I144_203.port1, 
  Loop Conditions: I144_197.port1=1, I144_200.port2=1, I144_201.port2=1, I144_203.port2=1, 
  (Signal Values: w_016_031=1, w_057_083=1, w_093_042=1, w_144_213=1, )

4)
  Loop Signals: w_144_202, w_144_208, w_144_209, w_144_210, w_144_211, w_144_213, 
  Loop Gates: I144_200.port2, I144_204.port1, I144_205.port1, I144_206.port1, I144_207.port1, I144_208.port2, 
  Loop Conditions: I144_200.port2=1, I144_205.port2=1, I144_206.port2=0, I144_208.port2=1, 
  (Signal Values: w_059_073=1, w_061_096=0, w_144_213=1, w_144_211=1, )

5)
  Loop Signals: w_029_011, w_029_012, w_029_013, w_029_014, w_029_015, w_029_016, w_029_017, w_029_018, w_029_019, w_029_020, 
  Loop Gates: I029_011.port2, I029_012.port2, I029_013.port1, I029_014.port1, I029_015.port1, I029_016.port2, I029_017.port1, I029_018.port1, I029_019.port1, I029_020.port1, 
  Loop Conditions: I029_011.port1=1, I029_012.port1=1, I029_016.port1=1, I029_018.port2=1, I029_020.port2=1, 
  (Signal Values: w_002_029=1, w_005_058=1, w_016_067=1, w_027_006=1, w_028_132=1, )

6)
  Loop Signals: w_021_178, w_021_179, w_021_180, w_021_181, w_021_182, w_021_183, 
  Loop Gates: I021_172.port1, I021_173.port1, I021_174.port2, I021_175.port1, I021_176.port2, I021_177.port1, 
  Loop Conditions: I021_172.port2=1, I021_174.port1=1, I021_175.port2=1, I021_176.port1=0, I021_177.port2=1, 
  (Signal Values: w_001_003=1, w_003_002=1, w_002_060=1, w_008_071=0, w_020_008=1, )

7)
  Loop Signals: w_133_153, w_133_154, w_133_155, w_133_156, w_133_157, w_133_158, w_133_159, w_133_160, w_133_161, w_133_162, w_133_163, w_133_164, 
  Loop Gates: I133_153.port2, I133_154.port1, I133_155.port2, I133_156.port1, I133_157.port1, I133_158.port1, I133_159.port1, I133_160.port1, I133_161.port1, I133_162.port2, I133_163.port1, I133_164.port1, 
  Loop Conditions: I133_153.port1=1, I133_154.port2=1, I133_155.port1=1, I133_156.port2=1, I133_157.port2=1, I133_158.port2=0, I133_160.port2=1, I133_162.port1=1, I133_164.port2=1, 
  (Signal Values: w_015_064=1, w_032_029=1, w_036_006=1, w_053_032=1, w_072_103=1, w_075_036=1, w_078_024=0, w_096_015=1, w_106_000=1, )

8)
  Loop Signals: w_039_012, w_039_025, w_039_026, w_039_027, w_039_028, w_039_029, w_039_030, w_039_031, w_039_032, w_039_033, w_039_034, w_039_036, 
  Loop Gates: I039_011.port2, I039_022.port1, I039_023.port1, I039_024.port1, I039_025.port1, I039_026.port1, I039_027.port2, I039_028.port2, I039_029.port1, I039_030.port1, I039_031.port1, I039_032.port2, 
  Loop Conditions: I039_011.port2=1, I039_022.port2=1, I039_024.port2=1, I039_025.port2=1, I039_026.port2=0, I039_027.port1=0, I039_028.port1=1, I039_029.port2=1, I039_032.port2=1, 
  (Signal Values: w_007_013=1, w_023_036=0, w_028_010=1, w_028_066=1, w_029_009=1, w_035_070=1, w_039_034=1, w_039_036=1, )** The loop condition cannot be reached.


9)
  Loop Signals: w_150_008, w_150_009, w_150_010, w_150_011, w_150_012, w_150_013, w_150_014, w_150_015, w_150_016, 
  Loop Gates: I150_007.port1, I150_008.port1, I150_009.port2, I150_010.port1, I150_011.port1, I150_012.port1, I150_013.port1, I150_014.port2, I150_015.port2, 
  Loop Conditions: I150_009.port1=0, I150_012.port2=1, I150_013.port2=1, I150_014.port1=0, I150_015.port1=0, 
  (Signal Values: w_006_015=0, w_060_049=1, w_071_017=0, w_096_009=0, w_130_176=1, )

******* result_4.txt *********
1)
  Loop Breaker: I028_159.port0-w_028_161-Register-w_028_161'-I028_160.port1 

2)
  Loop Breaker: I114_103.port0-w_114_108-Register-w_114_108'-I114_104.port1 

3)
  Loop Breaker: I144_200.port0-w_144_202-Register-w_144_202'-I144_201.port1 

4)
  Loop Breaker: I144_200.port0-w_144_202-Register-w_144_202'-I144_207.port1 

5)
  Loop Breaker: I029_011.port0-w_029_012-Register-w_029_012'-I029_012.port2 

6)
  Loop Breaker: I021_172.port0-w_021_179-Register-w_021_179'-I021_173.port1 

7)
  Loop Breaker: I133_153.port0-w_133_154-Register-w_133_154'-I133_154.port1 

8)
  Loop Breaker: I039_011.port0-w_039_012-Register-w_039_012'-I039_031.port1 

9)
  Loop Breaker: I150_007.port0-w_150_009-Register-w_150_009'-I150_008.port1 

// ******* The results for this case End *********
*/

// Gate Level Verilog Code Generated!
// GateLvl:1000 GateNum:1000 GateInputNum:2
// ****** Basic Gate Module Defination ******
module or2(out, in1, in2);
  output out;
  input in1, in2;
  wire in1, in2, out;
  assign out = in1 || in2;
endmodule

module and2(out, in1, in2);
  output out;
  input in1, in2;
  wire in1, in2, out;
  assign out = in1 && in2;
endmodule

module not1(out, in);
  output out;
  input in;
  wire in,out;
  assign out = ~in;
endmodule

module nand2(out, in1, in2);
  output out;
  input in1, in2;
  wire in1, in2, out;
  assign out = ~(in1 && in2);
endmodule
// ****** Basic Gate Module Defination End ******

// ****** Combined Logic Module Defination ******
module combLogic( w_000_000, w_000_001, w_000_002, w_000_003, w_000_004, w_000_005, w_000_006, w_000_007, w_000_008, w_000_009, w_000_010, w_000_011, w_000_012, w_000_013, w_000_014, w_000_015, w_000_016, w_000_017, w_000_018, w_000_019, w_000_020, w_000_021, w_000_022, w_000_023, w_000_024, w_000_025, w_000_026, w_000_027, w_000_028, w_000_029, w_000_030, w_000_031, w_000_032, w_000_033, w_000_034, w_000_035, w_000_036, w_000_037, w_000_038, w_000_039, w_000_040, w_000_041, w_000_042, w_000_043, w_000_044, w_000_045, w_000_046, w_000_047, w_000_048, w_000_049, w_000_050, w_000_051, w_000_052, w_000_053, w_000_054, w_000_055, w_000_056, w_000_057, w_000_058, w_000_059, w_000_060, w_000_061, w_000_062, w_000_063, w_000_064, w_000_065, w_000_066, w_000_067, w_000_068, w_000_069, w_000_070, w_000_071, w_000_072, w_000_073, w_000_074, w_000_075, w_000_076, w_000_077, w_000_078, w_000_079, w_000_080, w_000_081, w_000_082, w_000_083, w_000_084, w_000_085, w_000_086, w_000_087, w_000_088, w_000_089, w_000_090, w_000_091, w_000_092, w_000_093, w_000_094, w_000_095, w_000_096, w_000_097, w_000_098, w_000_099, w_000_100, w_000_101, w_000_102, w_000_103, w_000_104, w_000_105, w_000_106, w_000_107, w_000_108, w_000_109, w_000_110, w_000_111, w_000_112, w_000_113, w_000_114, w_000_115, w_000_116, w_000_117, w_000_118, w_000_119, w_000_120, w_000_121, w_000_122, w_000_123, w_000_124, w_000_125, w_000_126, w_000_127, w_000_128, w_000_129, w_000_130, w_000_131, w_000_132, w_000_133, w_000_134, w_000_135, w_000_136, w_000_137, w_000_138, w_000_139, w_000_140, w_000_141, w_000_142, w_000_143, w_000_144, w_000_145, w_000_146, w_000_147, w_000_148, w_000_149, w_000_150, w_000_151, w_000_152, w_000_153, w_000_154, w_000_155, w_000_156, w_000_157, w_000_158, w_000_159, w_000_160, w_000_161, w_000_162, w_000_163, w_000_164, w_000_165, w_000_166, w_000_167, w_000_168, w_000_169, w_000_170, w_000_171, w_000_172, w_000_173, w_000_174, w_000_175, w_000_176, w_000_177, w_000_178, w_000_179, w_000_180, w_000_181, w_000_182, w_000_183, w_000_184, w_000_185, w_000_186, w_000_187, w_000_188, w_000_189, w_000_190, w_000_191, w_000_192, w_000_193, w_000_194, w_000_195, w_000_196, w_000_197, w_000_198, w_000_199, w_000_200, w_000_201, w_000_202, w_000_203, w_000_204, w_000_205, w_000_206, w_000_207, w_000_208, w_000_209, w_000_210, w_000_211, w_000_212, w_000_213, w_000_214, w_000_215, w_000_216, w_000_217, w_000_218, w_000_219, w_000_220, w_000_221, w_000_222, w_000_223, w_000_224, w_000_225, w_000_226, w_000_227, w_000_228, w_000_230, w_000_231, w_000_232, w_000_233, w_000_234, w_000_235, w_000_236, w_000_237, w_000_238, w_000_239, w_000_240, w_000_241, w_000_242, w_000_243, w_000_244, w_000_245, w_000_246, w_000_247, w_000_248, w_000_249, w_000_250, w_000_251, w_000_252, w_000_253, w_000_254, w_000_255, w_000_256, w_000_257, w_000_258, w_000_259, w_000_260, w_000_262, w_000_263, w_000_264, w_000_265, w_000_266, w_000_267, w_000_268, w_000_269, w_000_270, w_000_271, w_000_272, w_000_273, w_000_274, w_000_275, w_000_276, w_000_277, w_000_278, w_000_279, w_000_280, w_000_281, w_000_282, w_000_283, w_000_284, w_000_285, w_000_286, w_000_287, w_000_288, w_000_289, w_000_290, w_000_291, w_000_292, w_000_293, w_000_294, w_000_295, w_000_296, w_000_297, w_000_298, w_000_299, w_000_300, w_000_301, w_000_302, w_000_303, w_000_304, w_000_305, w_000_306, w_000_307, w_000_308, w_000_309, w_000_310, w_000_311, w_000_312, w_000_313, w_000_314, w_000_315, w_000_316, w_000_317, w_000_318, w_000_319, w_000_320, w_000_321, w_000_322, w_000_323, w_000_324, w_000_325, w_000_326, w_000_327, w_000_328, w_000_329, w_000_330, w_000_331, w_000_332, w_000_333, w_000_334, w_000_335, w_000_336, w_000_337, w_000_338, w_000_339, w_000_340, w_000_341, w_000_342, w_000_343, w_000_344, w_000_345, w_000_346, w_000_347, w_000_348, w_000_349, w_000_350, w_000_351, w_000_352, w_000_353, w_000_354, w_000_355, w_000_356, w_000_357, w_000_358, w_000_359, w_000_360, w_000_361, w_000_362, w_000_364, w_000_365, w_000_366, w_000_367, w_000_369, w_000_370, w_000_371, w_000_372, w_000_373, w_000_374, w_000_375, w_000_376, w_000_377, w_000_378, w_000_379, w_000_380, w_000_381, w_000_382, w_000_383, w_000_384, w_000_385, w_000_386, w_000_387, w_000_388, w_000_389, w_000_390, w_000_391, w_000_392, w_000_393, w_000_394, w_000_395, w_000_396, w_000_397, w_000_398, w_000_399, w_000_400, w_000_401, w_000_402, w_000_403, w_000_404, w_000_405, w_000_406, w_000_407, w_000_408, w_000_409, w_000_410, w_000_411, w_000_412, w_000_413, w_000_414, w_000_415, w_000_416, w_000_417, w_000_418, w_000_419, w_000_420, w_000_421, w_000_422, w_000_423, w_000_424, w_000_425, w_000_426, w_000_427, w_000_428, w_000_429, w_000_430, w_000_431, w_000_432, w_000_433, w_000_434, w_000_435, w_000_436, w_000_437, w_000_438, w_000_439, w_000_440, w_000_441, w_000_442, w_000_443, w_000_444, w_000_445, w_000_446, w_000_447, w_000_448, w_000_449, w_000_450, w_000_451, w_000_452, w_000_453, w_000_454, w_000_455, w_000_456, w_000_457, w_000_458, w_000_459, w_000_460, w_000_461, w_000_462, w_000_463, w_000_464, w_000_465, w_000_466, w_000_467, w_000_468, w_000_469, w_000_470, w_000_471, w_000_472, w_000_473, w_000_474, w_000_475, w_000_476, w_000_477, w_000_478, w_000_479, w_000_480, w_000_481, w_000_482, w_000_483, w_000_484, w_000_485, w_000_486, w_000_487, w_000_488, w_000_489, w_000_490, w_000_491, w_000_492, w_000_493, w_000_494, w_000_495, w_000_496, w_000_497, w_000_498, w_000_499, w_000_500, w_000_501, w_000_502, w_000_503, w_000_504, w_000_505, w_000_506, w_000_507, w_000_508, w_000_509, w_000_510, w_000_511, w_000_512, w_000_513, w_000_514, w_000_515, w_000_516, w_000_517, w_000_518, w_000_519, w_000_520, w_000_521, w_000_522, w_000_523, w_000_524, w_000_525, w_000_526, w_000_527, w_000_528, w_000_529, w_000_530, w_000_531, w_000_532, w_000_533, w_000_534, w_000_535, w_000_536, w_000_537, w_000_538, w_000_539, w_000_540, w_000_541, w_000_542, w_000_543, w_000_544, w_000_545, w_000_546, w_000_547, w_000_548, w_000_549, w_000_550, w_000_551, w_000_552, w_000_553, w_000_554, w_000_555, w_000_556, w_000_557, w_000_558, w_000_559, w_000_560, w_000_561, w_000_562, w_000_563, w_000_564, w_000_565, w_000_566, w_000_567, w_000_568, w_000_569, w_000_570, w_000_571, w_000_572, w_000_573, w_000_574, w_000_575, w_000_576, w_000_577, w_000_578, w_000_579, w_000_580, w_000_581, w_000_582, w_000_583, w_000_584, w_000_585, w_000_586, w_000_587, w_000_588, w_000_589, w_000_590, w_000_591, w_000_592, w_000_593, w_000_594, w_000_595, w_000_596, w_000_597, w_000_598, w_000_599, w_000_600, w_000_601, w_000_602, w_000_603, w_000_604, w_000_605, w_000_606, w_000_607, w_000_608, w_000_609, w_000_610, w_000_611, w_000_612, w_000_613, w_000_614, w_000_615, w_000_616, w_000_617, w_000_618, w_000_619, w_000_620, w_000_621, w_000_622, w_000_623, w_000_624, w_000_625, w_000_626, w_000_627, w_000_628, w_000_629, w_000_630, w_000_631, w_000_632, w_000_633, w_000_634, w_000_635, w_000_636, w_000_637, w_000_638, w_000_639, w_000_640, w_000_641, w_000_642, w_000_643, w_000_644, w_000_645, w_000_646, w_000_647, w_000_648, w_000_649, w_000_650, w_000_651, w_000_652, w_000_653, w_000_654, w_000_655, w_000_656, w_000_657, w_000_658, w_000_659, w_000_660, w_000_661, w_000_662, w_000_663, w_000_664, w_000_665, w_000_666, w_000_667, w_000_669, w_000_670, w_000_671, w_000_672, w_000_673, w_000_674, w_000_675, w_000_676, w_000_677, w_000_678, w_000_679, w_000_680, w_000_681, w_000_682, w_000_683, w_000_684, w_000_685, w_000_686, w_000_687, w_000_688, w_000_689, w_000_690, w_000_691, w_000_692, w_000_693, w_000_694, w_000_695, w_000_696, w_000_697, w_000_698, w_000_699, w_000_700, w_000_701, w_000_702, w_000_703, w_000_704, w_000_705, w_000_706, w_000_707, w_000_708, w_000_709, w_000_710, w_000_711, w_000_712, w_000_713, w_000_714, w_000_715, w_000_716, w_000_717, w_000_718, w_000_719, w_000_720, w_000_721, w_000_722, w_000_723, w_000_724, w_000_725, w_000_726, w_000_727, w_000_728, w_000_729, w_000_730, w_000_731, w_000_732, w_000_733, w_000_734, w_000_735, w_000_736, w_000_737, w_000_738, w_000_739, w_000_740, w_000_741, w_000_742, w_000_743, w_000_744, w_000_745, w_000_746, w_000_747, w_000_748, w_000_749, w_000_750, w_000_751, w_000_752, w_000_753, w_000_754, w_000_755, w_000_756, w_000_757, w_000_758, w_000_759, w_000_760, w_000_761, w_000_762, w_000_763, w_000_765, w_000_766, w_000_767, w_000_769, w_000_770, w_000_772, w_000_773, w_000_774, w_000_775, w_000_776, w_000_777, w_000_779, w_000_780, w_000_781, w_000_782, w_000_783, w_000_784, w_000_785, w_000_786, w_000_787, w_000_788, w_000_789, w_000_790, w_000_791, w_000_792, w_000_793, w_000_794, w_000_795, w_000_796, w_000_797, w_000_798, w_000_799, w_000_801, w_000_802, w_000_803, w_000_804, w_000_805, w_000_806, w_000_807, w_000_808, w_000_809, w_000_810, w_000_811, w_000_812, w_000_813, w_000_814, w_000_815, w_000_816, w_000_817, w_000_818, w_000_819, w_000_820, w_000_821, w_000_822, w_000_823, w_000_824, w_000_825, w_000_826, w_000_827, w_000_828, w_000_829, w_000_830, w_000_831, w_000_832, w_000_833, w_000_834, w_000_835, w_000_836, w_000_837, w_000_838, w_000_839, w_000_840, w_000_841, w_000_842, w_000_843, w_000_844, w_000_845, w_000_846, w_000_847, w_000_848, w_000_849, w_000_850, w_000_851, w_000_852, w_000_853, w_000_854, w_000_855, w_000_856, w_000_857, w_000_858, w_000_859, w_000_860, w_000_861, w_000_862, w_000_863, w_000_864, w_000_865, w_000_866, w_000_867, w_000_868, w_000_869, w_000_870, w_000_871, w_000_872, w_000_873, w_000_874, w_000_875, w_000_876, w_000_877, w_000_878, w_000_879, w_000_880, w_000_881, w_000_882, w_000_883, w_000_885, w_000_886, w_000_887, w_000_889, w_000_890, w_000_891, w_000_893, w_000_894, w_000_895, w_000_896, w_000_897, w_000_898, w_000_899, w_000_900, w_000_901, w_000_903, w_000_904, w_000_905, w_000_906, w_000_907, w_000_908, w_000_909, w_000_910, w_000_912, w_000_914, w_000_915, w_000_916, w_000_917, w_000_918, w_000_919, w_000_923, w_000_924, w_000_925, w_000_926, w_000_928, w_000_929, w_000_930, w_000_931, w_000_932, w_000_934, w_000_935, w_000_936, w_000_937, w_000_938, w_000_939, w_000_943, w_000_944, w_000_945, w_000_947, w_000_949, w_000_950, w_000_952, w_000_953, w_000_954, w_000_955, w_000_956, w_000_958, w_000_959, w_000_960, w_000_963, w_000_964, w_000_965, w_000_967, w_000_968, w_000_969, w_000_970, w_000_971, w_000_977, w_000_979, w_000_980, w_000_981, w_000_982, w_000_983, w_1000_000, w_1000_001, w_1000_002, w_1000_003, w_1000_004, w_1000_005, w_1000_006, w_1000_007, w_1000_008, w_1000_009, w_1000_010, w_1000_011, w_1000_012, w_1000_013, w_1000_014, w_1000_015, w_1000_016, w_1000_017, w_1000_018, w_1000_019, w_1000_020, w_1000_021, w_1000_022, w_1000_023, w_1000_024, w_1000_025, w_1000_026, w_1000_027, w_1000_028, w_1000_029, w_1000_030, w_1000_031, w_1000_032, w_1000_033, w_1000_034, w_1000_035, w_1000_036, w_1000_037, w_1000_038, w_1000_039, w_1000_040, w_1000_041, w_1000_042, w_1000_043, w_1000_044, w_1000_045, w_1000_046, w_1000_047, w_1000_048, w_1000_049, w_1000_050, w_1000_051, w_1000_052, w_1000_053, w_1000_054, w_1000_055, w_1000_056, w_1000_057, w_1000_058, w_1000_059, w_1000_060, w_1000_061, w_1000_062, w_1000_063, w_1000_064, w_1000_065, w_1000_066, w_1000_067, w_1000_068, w_1000_069, w_1000_070, w_1000_071, w_1000_072, w_1000_073, w_1000_074, w_1000_075, w_1000_076, w_1000_077, w_1000_078, w_1000_079, w_1000_080, w_1000_081, w_1000_082, w_1000_083, w_1000_084, w_1000_085, w_1000_086, w_1000_087, w_1000_088, w_1000_089, w_1000_090, w_1000_091, w_1000_092, w_1000_093, w_1000_094, w_1000_095, w_1000_096, w_1000_097, w_1000_098, w_1000_099, w_1000_100, w_1000_101, w_1000_102, w_1000_103, w_1000_104, w_1000_105, w_1000_106, w_1000_107, w_1000_108, w_1000_109, w_1000_110, w_1000_111, w_1000_112, w_1000_113, w_1000_114, w_1000_115, w_1000_116, w_1000_117, w_1000_118, w_1000_119, w_1000_120, w_1000_121, w_1000_122, w_1000_123, w_1000_124, w_1000_125, w_1000_126, w_1000_127, w_1000_128, w_1000_129, w_1000_130, w_1000_131, w_1000_132, w_1000_133, w_1000_134, w_1000_135, w_1000_136, w_1000_137, w_1000_138, w_1000_139, w_1000_140, w_1000_141, w_1000_142, w_1000_143, w_1000_144, w_1000_145, w_1000_146, w_1000_147, w_1000_148, w_1000_149, w_1000_150, w_1000_151, w_1000_152, w_1000_153, w_1000_154, w_1000_155, w_1000_156, w_1000_157, w_1000_158, w_1000_159, w_1000_160, w_1000_161, w_1000_162, w_1000_163, w_1000_164, w_1000_165, w_1000_166, w_1000_167, w_1000_168, w_1000_169, w_1000_170, w_1000_171, w_1000_172, w_1000_173, w_1000_174, w_1000_175, w_1000_176, w_1000_177, w_1000_178, w_1000_179, w_1000_180, w_1000_181, w_1000_182, w_1000_183, w_1000_184, w_1000_185 );
  inout w_000_000, w_000_001, w_000_002, w_000_003, w_000_004, w_000_005, w_000_006, w_000_007, w_000_008, w_000_009, w_000_010, w_000_011, w_000_012, w_000_013, w_000_014, w_000_015, w_000_016, w_000_017, w_000_018, w_000_019, w_000_020, w_000_021, w_000_022, w_000_023, w_000_024, w_000_025, w_000_026, w_000_027, w_000_028, w_000_029, w_000_030, w_000_031, w_000_032, w_000_033, w_000_034, w_000_035, w_000_036, w_000_037, w_000_038, w_000_039, w_000_040, w_000_041, w_000_042, w_000_043, w_000_044, w_000_045, w_000_046, w_000_047, w_000_048, w_000_049, w_000_050, w_000_051, w_000_052, w_000_053, w_000_054, w_000_055, w_000_056, w_000_057, w_000_058, w_000_059, w_000_060, w_000_061, w_000_062, w_000_063, w_000_064, w_000_065, w_000_066, w_000_067, w_000_068, w_000_069, w_000_070, w_000_071, w_000_072, w_000_073, w_000_074, w_000_075, w_000_076, w_000_077, w_000_078, w_000_079, w_000_080, w_000_081, w_000_082, w_000_083, w_000_084, w_000_085, w_000_086, w_000_087, w_000_088, w_000_089, w_000_090, w_000_091, w_000_092, w_000_093, w_000_094, w_000_095, w_000_096, w_000_097, w_000_098, w_000_099, w_000_100, w_000_101, w_000_102, w_000_103, w_000_104, w_000_105, w_000_106, w_000_107, w_000_108, w_000_109, w_000_110, w_000_111, w_000_112, w_000_113, w_000_114, w_000_115, w_000_116, w_000_117, w_000_118, w_000_119, w_000_120, w_000_121, w_000_122, w_000_123, w_000_124, w_000_125, w_000_126, w_000_127, w_000_128, w_000_129, w_000_130, w_000_131, w_000_132, w_000_133, w_000_134, w_000_135, w_000_136, w_000_137, w_000_138, w_000_139, w_000_140, w_000_141, w_000_142, w_000_143, w_000_144, w_000_145, w_000_146, w_000_147, w_000_148, w_000_149, w_000_150, w_000_151, w_000_152, w_000_153, w_000_154, w_000_155, w_000_156, w_000_157, w_000_158, w_000_159, w_000_160, w_000_161, w_000_162, w_000_163, w_000_164, w_000_165, w_000_166, w_000_167, w_000_168, w_000_169, w_000_170, w_000_171, w_000_172, w_000_173, w_000_174, w_000_175, w_000_176, w_000_177, w_000_178, w_000_179, w_000_180, w_000_181, w_000_182, w_000_183, w_000_184, w_000_185, w_000_186, w_000_187, w_000_188, w_000_189, w_000_190, w_000_191, w_000_192, w_000_193, w_000_194, w_000_195, w_000_196, w_000_197, w_000_198, w_000_199, w_000_200, w_000_201, w_000_202, w_000_203, w_000_204, w_000_205, w_000_206, w_000_207, w_000_208, w_000_209, w_000_210, w_000_211, w_000_212, w_000_213, w_000_214, w_000_215, w_000_216, w_000_217, w_000_218, w_000_219, w_000_220, w_000_221, w_000_222, w_000_223, w_000_224, w_000_225, w_000_226, w_000_227, w_000_228, w_000_230, w_000_231, w_000_232, w_000_233, w_000_234, w_000_235, w_000_236, w_000_237, w_000_238, w_000_239, w_000_240, w_000_241, w_000_242, w_000_243, w_000_244, w_000_245, w_000_246, w_000_247, w_000_248, w_000_249, w_000_250, w_000_251, w_000_252, w_000_253, w_000_254, w_000_255, w_000_256, w_000_257, w_000_258, w_000_259, w_000_260, w_000_262, w_000_263, w_000_264, w_000_265, w_000_266, w_000_267, w_000_268, w_000_269, w_000_270, w_000_271, w_000_272, w_000_273, w_000_274, w_000_275, w_000_276, w_000_277, w_000_278, w_000_279, w_000_280, w_000_281, w_000_282, w_000_283, w_000_284, w_000_285, w_000_286, w_000_287, w_000_288, w_000_289, w_000_290, w_000_291, w_000_292, w_000_293, w_000_294, w_000_295, w_000_296, w_000_297, w_000_298, w_000_299, w_000_300, w_000_301, w_000_302, w_000_303, w_000_304, w_000_305, w_000_306, w_000_307, w_000_308, w_000_309, w_000_310, w_000_311, w_000_312, w_000_313, w_000_314, w_000_315, w_000_316, w_000_317, w_000_318, w_000_319, w_000_320, w_000_321, w_000_322, w_000_323, w_000_324, w_000_325, w_000_326, w_000_327, w_000_328, w_000_329, w_000_330, w_000_331, w_000_332, w_000_333, w_000_334, w_000_335, w_000_336, w_000_337, w_000_338, w_000_339, w_000_340, w_000_341, w_000_342, w_000_343, w_000_344, w_000_345, w_000_346, w_000_347, w_000_348, w_000_349, w_000_350, w_000_351, w_000_352, w_000_353, w_000_354, w_000_355, w_000_356, w_000_357, w_000_358, w_000_359, w_000_360, w_000_361, w_000_362, w_000_364, w_000_365, w_000_366, w_000_367, w_000_369, w_000_370, w_000_371, w_000_372, w_000_373, w_000_374, w_000_375, w_000_376, w_000_377, w_000_378, w_000_379, w_000_380, w_000_381, w_000_382, w_000_383, w_000_384, w_000_385, w_000_386, w_000_387, w_000_388, w_000_389, w_000_390, w_000_391, w_000_392, w_000_393, w_000_394, w_000_395, w_000_396, w_000_397, w_000_398, w_000_399, w_000_400, w_000_401, w_000_402, w_000_403, w_000_404, w_000_405, w_000_406, w_000_407, w_000_408, w_000_409, w_000_410, w_000_411, w_000_412, w_000_413, w_000_414, w_000_415, w_000_416, w_000_417, w_000_418, w_000_419, w_000_420, w_000_421, w_000_422, w_000_423, w_000_424, w_000_425, w_000_426, w_000_427, w_000_428, w_000_429, w_000_430, w_000_431, w_000_432, w_000_433, w_000_434, w_000_435, w_000_436, w_000_437, w_000_438, w_000_439, w_000_440, w_000_441, w_000_442, w_000_443, w_000_444, w_000_445, w_000_446, w_000_447, w_000_448, w_000_449, w_000_450, w_000_451, w_000_452, w_000_453, w_000_454, w_000_455, w_000_456, w_000_457, w_000_458, w_000_459, w_000_460, w_000_461, w_000_462, w_000_463, w_000_464, w_000_465, w_000_466, w_000_467, w_000_468, w_000_469, w_000_470, w_000_471, w_000_472, w_000_473, w_000_474, w_000_475, w_000_476, w_000_477, w_000_478, w_000_479, w_000_480, w_000_481, w_000_482, w_000_483, w_000_484, w_000_485, w_000_486, w_000_487, w_000_488, w_000_489, w_000_490, w_000_491, w_000_492, w_000_493, w_000_494, w_000_495, w_000_496, w_000_497, w_000_498, w_000_499, w_000_500, w_000_501, w_000_502, w_000_503, w_000_504, w_000_505, w_000_506, w_000_507, w_000_508, w_000_509, w_000_510, w_000_511, w_000_512, w_000_513, w_000_514, w_000_515, w_000_516, w_000_517, w_000_518, w_000_519, w_000_520, w_000_521, w_000_522, w_000_523, w_000_524, w_000_525, w_000_526, w_000_527, w_000_528, w_000_529, w_000_530, w_000_531, w_000_532, w_000_533, w_000_534, w_000_535, w_000_536, w_000_537, w_000_538, w_000_539, w_000_540, w_000_541, w_000_542, w_000_543, w_000_544, w_000_545, w_000_546, w_000_547, w_000_548, w_000_549, w_000_550, w_000_551, w_000_552, w_000_553, w_000_554, w_000_555, w_000_556, w_000_557, w_000_558, w_000_559, w_000_560, w_000_561, w_000_562, w_000_563, w_000_564, w_000_565, w_000_566, w_000_567, w_000_568, w_000_569, w_000_570, w_000_571, w_000_572, w_000_573, w_000_574, w_000_575, w_000_576, w_000_577, w_000_578, w_000_579, w_000_580, w_000_581, w_000_582, w_000_583, w_000_584, w_000_585, w_000_586, w_000_587, w_000_588, w_000_589, w_000_590, w_000_591, w_000_592, w_000_593, w_000_594, w_000_595, w_000_596, w_000_597, w_000_598, w_000_599, w_000_600, w_000_601, w_000_602, w_000_603, w_000_604, w_000_605, w_000_606, w_000_607, w_000_608, w_000_609, w_000_610, w_000_611, w_000_612, w_000_613, w_000_614, w_000_615, w_000_616, w_000_617, w_000_618, w_000_619, w_000_620, w_000_621, w_000_622, w_000_623, w_000_624, w_000_625, w_000_626, w_000_627, w_000_628, w_000_629, w_000_630, w_000_631, w_000_632, w_000_633, w_000_634, w_000_635, w_000_636, w_000_637, w_000_638, w_000_639, w_000_640, w_000_641, w_000_642, w_000_643, w_000_644, w_000_645, w_000_646, w_000_647, w_000_648, w_000_649, w_000_650, w_000_651, w_000_652, w_000_653, w_000_654, w_000_655, w_000_656, w_000_657, w_000_658, w_000_659, w_000_660, w_000_661, w_000_662, w_000_663, w_000_664, w_000_665, w_000_666, w_000_667, w_000_669, w_000_670, w_000_671, w_000_672, w_000_673, w_000_674, w_000_675, w_000_676, w_000_677, w_000_678, w_000_679, w_000_680, w_000_681, w_000_682, w_000_683, w_000_684, w_000_685, w_000_686, w_000_687, w_000_688, w_000_689, w_000_690, w_000_691, w_000_692, w_000_693, w_000_694, w_000_695, w_000_696, w_000_697, w_000_698, w_000_699, w_000_700, w_000_701, w_000_702, w_000_703, w_000_704, w_000_705, w_000_706, w_000_707, w_000_708, w_000_709, w_000_710, w_000_711, w_000_712, w_000_713, w_000_714, w_000_715, w_000_716, w_000_717, w_000_718, w_000_719, w_000_720, w_000_721, w_000_722, w_000_723, w_000_724, w_000_725, w_000_726, w_000_727, w_000_728, w_000_729, w_000_730, w_000_731, w_000_732, w_000_733, w_000_734, w_000_735, w_000_736, w_000_737, w_000_738, w_000_739, w_000_740, w_000_741, w_000_742, w_000_743, w_000_744, w_000_745, w_000_746, w_000_747, w_000_748, w_000_749, w_000_750, w_000_751, w_000_752, w_000_753, w_000_754, w_000_755, w_000_756, w_000_757, w_000_758, w_000_759, w_000_760, w_000_761, w_000_762, w_000_763, w_000_765, w_000_766, w_000_767, w_000_769, w_000_770, w_000_772, w_000_773, w_000_774, w_000_775, w_000_776, w_000_777, w_000_779, w_000_780, w_000_781, w_000_782, w_000_783, w_000_784, w_000_785, w_000_786, w_000_787, w_000_788, w_000_789, w_000_790, w_000_791, w_000_792, w_000_793, w_000_794, w_000_795, w_000_796, w_000_797, w_000_798, w_000_799, w_000_801, w_000_802, w_000_803, w_000_804, w_000_805, w_000_806, w_000_807, w_000_808, w_000_809, w_000_810, w_000_811, w_000_812, w_000_813, w_000_814, w_000_815, w_000_816, w_000_817, w_000_818, w_000_819, w_000_820, w_000_821, w_000_822, w_000_823, w_000_824, w_000_825, w_000_826, w_000_827, w_000_828, w_000_829, w_000_830, w_000_831, w_000_832, w_000_833, w_000_834, w_000_835, w_000_836, w_000_837, w_000_838, w_000_839, w_000_840, w_000_841, w_000_842, w_000_843, w_000_844, w_000_845, w_000_846, w_000_847, w_000_848, w_000_849, w_000_850, w_000_851, w_000_852, w_000_853, w_000_854, w_000_855, w_000_856, w_000_857, w_000_858, w_000_859, w_000_860, w_000_861, w_000_862, w_000_863, w_000_864, w_000_865, w_000_866, w_000_867, w_000_868, w_000_869, w_000_870, w_000_871, w_000_872, w_000_873, w_000_874, w_000_875, w_000_876, w_000_877, w_000_878, w_000_879, w_000_880, w_000_881, w_000_882, w_000_883, w_000_885, w_000_886, w_000_887, w_000_889, w_000_890, w_000_891, w_000_893, w_000_894, w_000_895, w_000_896, w_000_897, w_000_898, w_000_899, w_000_900, w_000_901, w_000_903, w_000_904, w_000_905, w_000_906, w_000_907, w_000_908, w_000_909, w_000_910, w_000_912, w_000_914, w_000_915, w_000_916, w_000_917, w_000_918, w_000_919, w_000_923, w_000_924, w_000_925, w_000_926, w_000_928, w_000_929, w_000_930, w_000_931, w_000_932, w_000_934, w_000_935, w_000_936, w_000_937, w_000_938, w_000_939, w_000_943, w_000_944, w_000_945, w_000_947, w_000_949, w_000_950, w_000_952, w_000_953, w_000_954, w_000_955, w_000_956, w_000_958, w_000_959, w_000_960, w_000_963, w_000_964, w_000_965, w_000_967, w_000_968, w_000_969, w_000_970, w_000_971, w_000_977, w_000_979, w_000_980, w_000_981, w_000_982, w_000_983;
  output w_1000_000, w_1000_001, w_1000_002, w_1000_003, w_1000_004, w_1000_005, w_1000_006, w_1000_007, w_1000_008, w_1000_009, w_1000_010, w_1000_011, w_1000_012, w_1000_013, w_1000_014, w_1000_015, w_1000_016, w_1000_017, w_1000_018, w_1000_019, w_1000_020, w_1000_021, w_1000_022, w_1000_023, w_1000_024, w_1000_025, w_1000_026, w_1000_027, w_1000_028, w_1000_029, w_1000_030, w_1000_031, w_1000_032, w_1000_033, w_1000_034, w_1000_035, w_1000_036, w_1000_037, w_1000_038, w_1000_039, w_1000_040, w_1000_041, w_1000_042, w_1000_043, w_1000_044, w_1000_045, w_1000_046, w_1000_047, w_1000_048, w_1000_049, w_1000_050, w_1000_051, w_1000_052, w_1000_053, w_1000_054, w_1000_055, w_1000_056, w_1000_057, w_1000_058, w_1000_059, w_1000_060, w_1000_061, w_1000_062, w_1000_063, w_1000_064, w_1000_065, w_1000_066, w_1000_067, w_1000_068, w_1000_069, w_1000_070, w_1000_071, w_1000_072, w_1000_073, w_1000_074, w_1000_075, w_1000_076, w_1000_077, w_1000_078, w_1000_079, w_1000_080, w_1000_081, w_1000_082, w_1000_083, w_1000_084, w_1000_085, w_1000_086, w_1000_087, w_1000_088, w_1000_089, w_1000_090, w_1000_091, w_1000_092, w_1000_093, w_1000_094, w_1000_095, w_1000_096, w_1000_097, w_1000_098, w_1000_099, w_1000_100, w_1000_101, w_1000_102, w_1000_103, w_1000_104, w_1000_105, w_1000_106, w_1000_107, w_1000_108, w_1000_109, w_1000_110, w_1000_111, w_1000_112, w_1000_113, w_1000_114, w_1000_115, w_1000_116, w_1000_117, w_1000_118, w_1000_119, w_1000_120, w_1000_121, w_1000_122, w_1000_123, w_1000_124, w_1000_125, w_1000_126, w_1000_127, w_1000_128, w_1000_129, w_1000_130, w_1000_131, w_1000_132, w_1000_133, w_1000_134, w_1000_135, w_1000_136, w_1000_137, w_1000_138, w_1000_139, w_1000_140, w_1000_141, w_1000_142, w_1000_143, w_1000_144, w_1000_145, w_1000_146, w_1000_147, w_1000_148, w_1000_149, w_1000_150, w_1000_151, w_1000_152, w_1000_153, w_1000_154, w_1000_155, w_1000_156, w_1000_157, w_1000_158, w_1000_159, w_1000_160, w_1000_161, w_1000_162, w_1000_163, w_1000_164, w_1000_165, w_1000_166, w_1000_167, w_1000_168, w_1000_169, w_1000_170, w_1000_171, w_1000_172, w_1000_173, w_1000_174, w_1000_175, w_1000_176, w_1000_177, w_1000_178, w_1000_179, w_1000_180, w_1000_181, w_1000_182, w_1000_183, w_1000_184, w_1000_185;
  wire w_000_000, w_000_001, w_000_002, w_000_003, w_000_004, w_000_005, w_000_006, w_000_007, w_000_008, w_000_009, w_000_010, w_000_011, w_000_012, w_000_013, w_000_014, w_000_015, w_000_016, w_000_017, w_000_018, w_000_019, w_000_020, w_000_021, w_000_022, w_000_023, w_000_024, w_000_025, w_000_026, w_000_027, w_000_028, w_000_029, w_000_030, w_000_031, w_000_032, w_000_033, w_000_034, w_000_035, w_000_036, w_000_037, w_000_038, w_000_039, w_000_040, w_000_041, w_000_042, w_000_043, w_000_044, w_000_045, w_000_046, w_000_047, w_000_048, w_000_049, w_000_050, w_000_051, w_000_052, w_000_053, w_000_054, w_000_055, w_000_056, w_000_057, w_000_058, w_000_059, w_000_060, w_000_061, w_000_062, w_000_063, w_000_064, w_000_065, w_000_066, w_000_067, w_000_068, w_000_069, w_000_070, w_000_071, w_000_072, w_000_073, w_000_074, w_000_075, w_000_076, w_000_077, w_000_078, w_000_079, w_000_080, w_000_081, w_000_082, w_000_083, w_000_084, w_000_085, w_000_086, w_000_087, w_000_088, w_000_089, w_000_090, w_000_091, w_000_092, w_000_093, w_000_094, w_000_095, w_000_096, w_000_097, w_000_098, w_000_099, w_000_100, w_000_101, w_000_102, w_000_103, w_000_104, w_000_105, w_000_106, w_000_107, w_000_108, w_000_109, w_000_110, w_000_111, w_000_112, w_000_113, w_000_114, w_000_115, w_000_116, w_000_117, w_000_118, w_000_119, w_000_120, w_000_121, w_000_122, w_000_123, w_000_124, w_000_125, w_000_126, w_000_127, w_000_128, w_000_129, w_000_130, w_000_131, w_000_132, w_000_133, w_000_134, w_000_135, w_000_136, w_000_137, w_000_138, w_000_139, w_000_140, w_000_141, w_000_142, w_000_143, w_000_144, w_000_145, w_000_146, w_000_147, w_000_148, w_000_149, w_000_150, w_000_151, w_000_152, w_000_153, w_000_154, w_000_155, w_000_156, w_000_157, w_000_158, w_000_159, w_000_160, w_000_161, w_000_162, w_000_163, w_000_164, w_000_165, w_000_166, w_000_167, w_000_168, w_000_169, w_000_170, w_000_171, w_000_172, w_000_173, w_000_174, w_000_175, w_000_176, w_000_177, w_000_178, w_000_179, w_000_180, w_000_181, w_000_182, w_000_183, w_000_184, w_000_185, w_000_186, w_000_187, w_000_188, w_000_189, w_000_190, w_000_191, w_000_192, w_000_193, w_000_194, w_000_195, w_000_196, w_000_197, w_000_198, w_000_199, w_000_200, w_000_201, w_000_202, w_000_203, w_000_204, w_000_205, w_000_206, w_000_207, w_000_208, w_000_209, w_000_210, w_000_211, w_000_212, w_000_213, w_000_214, w_000_215, w_000_216, w_000_217, w_000_218, w_000_219, w_000_220, w_000_221, w_000_222, w_000_223, w_000_224, w_000_225, w_000_226, w_000_227, w_000_228, w_000_230, w_000_231, w_000_232, w_000_233, w_000_234, w_000_235, w_000_236, w_000_237, w_000_238, w_000_239, w_000_240, w_000_241, w_000_242, w_000_243, w_000_244, w_000_245, w_000_246, w_000_247, w_000_248, w_000_249, w_000_250, w_000_251, w_000_252, w_000_253, w_000_254, w_000_255, w_000_256, w_000_257, w_000_258, w_000_259, w_000_260, w_000_262, w_000_263, w_000_264, w_000_265, w_000_266, w_000_267, w_000_268, w_000_269, w_000_270, w_000_271, w_000_272, w_000_273, w_000_274, w_000_275, w_000_276, w_000_277, w_000_278, w_000_279, w_000_280, w_000_281, w_000_282, w_000_283, w_000_284, w_000_285, w_000_286, w_000_287, w_000_288, w_000_289, w_000_290, w_000_291, w_000_292, w_000_293, w_000_294, w_000_295, w_000_296, w_000_297, w_000_298, w_000_299, w_000_300, w_000_301, w_000_302, w_000_303, w_000_304, w_000_305, w_000_306, w_000_307, w_000_308, w_000_309, w_000_310, w_000_311, w_000_312, w_000_313, w_000_314, w_000_315, w_000_316, w_000_317, w_000_318, w_000_319, w_000_320, w_000_321, w_000_322, w_000_323, w_000_324, w_000_325, w_000_326, w_000_327, w_000_328, w_000_329, w_000_330, w_000_331, w_000_332, w_000_333, w_000_334, w_000_335, w_000_336, w_000_337, w_000_338, w_000_339, w_000_340, w_000_341, w_000_342, w_000_343, w_000_344, w_000_345, w_000_346, w_000_347, w_000_348, w_000_349, w_000_350, w_000_351, w_000_352, w_000_353, w_000_354, w_000_355, w_000_356, w_000_357, w_000_358, w_000_359, w_000_360, w_000_361, w_000_362, w_000_364, w_000_365, w_000_366, w_000_367, w_000_369, w_000_370, w_000_371, w_000_372, w_000_373, w_000_374, w_000_375, w_000_376, w_000_377, w_000_378, w_000_379, w_000_380, w_000_381, w_000_382, w_000_383, w_000_384, w_000_385, w_000_386, w_000_387, w_000_388, w_000_389, w_000_390, w_000_391, w_000_392, w_000_393, w_000_394, w_000_395, w_000_396, w_000_397, w_000_398, w_000_399, w_000_400, w_000_401, w_000_402, w_000_403, w_000_404, w_000_405, w_000_406, w_000_407, w_000_408, w_000_409, w_000_410, w_000_411, w_000_412, w_000_413, w_000_414, w_000_415, w_000_416, w_000_417, w_000_418, w_000_419, w_000_420, w_000_421, w_000_422, w_000_423, w_000_424, w_000_425, w_000_426, w_000_427, w_000_428, w_000_429, w_000_430, w_000_431, w_000_432, w_000_433, w_000_434, w_000_435, w_000_436, w_000_437, w_000_438, w_000_439, w_000_440, w_000_441, w_000_442, w_000_443, w_000_444, w_000_445, w_000_446, w_000_447, w_000_448, w_000_449, w_000_450, w_000_451, w_000_452, w_000_453, w_000_454, w_000_455, w_000_456, w_000_457, w_000_458, w_000_459, w_000_460, w_000_461, w_000_462, w_000_463, w_000_464, w_000_465, w_000_466, w_000_467, w_000_468, w_000_469, w_000_470, w_000_471, w_000_472, w_000_473, w_000_474, w_000_475, w_000_476, w_000_477, w_000_478, w_000_479, w_000_480, w_000_481, w_000_482, w_000_483, w_000_484, w_000_485, w_000_486, w_000_487, w_000_488, w_000_489, w_000_490, w_000_491, w_000_492, w_000_493, w_000_494, w_000_495, w_000_496, w_000_497, w_000_498, w_000_499, w_000_500, w_000_501, w_000_502, w_000_503, w_000_504, w_000_505, w_000_506, w_000_507, w_000_508, w_000_509, w_000_510, w_000_511, w_000_512, w_000_513, w_000_514, w_000_515, w_000_516, w_000_517, w_000_518, w_000_519, w_000_520, w_000_521, w_000_522, w_000_523, w_000_524, w_000_525, w_000_526, w_000_527, w_000_528, w_000_529, w_000_530, w_000_531, w_000_532, w_000_533, w_000_534, w_000_535, w_000_536, w_000_537, w_000_538, w_000_539, w_000_540, w_000_541, w_000_542, w_000_543, w_000_544, w_000_545, w_000_546, w_000_547, w_000_548, w_000_549, w_000_550, w_000_551, w_000_552, w_000_553, w_000_554, w_000_555, w_000_556, w_000_557, w_000_558, w_000_559, w_000_560, w_000_561, w_000_562, w_000_563, w_000_564, w_000_565, w_000_566, w_000_567, w_000_568, w_000_569, w_000_570, w_000_571, w_000_572, w_000_573, w_000_574, w_000_575, w_000_576, w_000_577, w_000_578, w_000_579, w_000_580, w_000_581, w_000_582, w_000_583, w_000_584, w_000_585, w_000_586, w_000_587, w_000_588, w_000_589, w_000_590, w_000_591, w_000_592, w_000_593, w_000_594, w_000_595, w_000_596, w_000_597, w_000_598, w_000_599, w_000_600, w_000_601, w_000_602, w_000_603, w_000_604, w_000_605, w_000_606, w_000_607, w_000_608, w_000_609, w_000_610, w_000_611, w_000_612, w_000_613, w_000_614, w_000_615, w_000_616, w_000_617, w_000_618, w_000_619, w_000_620, w_000_621, w_000_622, w_000_623, w_000_624, w_000_625, w_000_626, w_000_627, w_000_628, w_000_629, w_000_630, w_000_631, w_000_632, w_000_633, w_000_634, w_000_635, w_000_636, w_000_637, w_000_638, w_000_639, w_000_640, w_000_641, w_000_642, w_000_643, w_000_644, w_000_645, w_000_646, w_000_647, w_000_648, w_000_649, w_000_650, w_000_651, w_000_652, w_000_653, w_000_654, w_000_655, w_000_656, w_000_657, w_000_658, w_000_659, w_000_660, w_000_661, w_000_662, w_000_663, w_000_664, w_000_665, w_000_666, w_000_667, w_000_669, w_000_670, w_000_671, w_000_672, w_000_673, w_000_674, w_000_675, w_000_676, w_000_677, w_000_678, w_000_679, w_000_680, w_000_681, w_000_682, w_000_683, w_000_684, w_000_685, w_000_686, w_000_687, w_000_688, w_000_689, w_000_690, w_000_691, w_000_692, w_000_693, w_000_694, w_000_695, w_000_696, w_000_697, w_000_698, w_000_699, w_000_700, w_000_701, w_000_702, w_000_703, w_000_704, w_000_705, w_000_706, w_000_707, w_000_708, w_000_709, w_000_710, w_000_711, w_000_712, w_000_713, w_000_714, w_000_715, w_000_716, w_000_717, w_000_718, w_000_719, w_000_720, w_000_721, w_000_722, w_000_723, w_000_724, w_000_725, w_000_726, w_000_727, w_000_728, w_000_729, w_000_730, w_000_731, w_000_732, w_000_733, w_000_734, w_000_735, w_000_736, w_000_737, w_000_738, w_000_739, w_000_740, w_000_741, w_000_742, w_000_743, w_000_744, w_000_745, w_000_746, w_000_747, w_000_748, w_000_749, w_000_750, w_000_751, w_000_752, w_000_753, w_000_754, w_000_755, w_000_756, w_000_757, w_000_758, w_000_759, w_000_760, w_000_761, w_000_762, w_000_763, w_000_765, w_000_766, w_000_767, w_000_769, w_000_770, w_000_772, w_000_773, w_000_774, w_000_775, w_000_776, w_000_777, w_000_779, w_000_780, w_000_781, w_000_782, w_000_783, w_000_784, w_000_785, w_000_786, w_000_787, w_000_788, w_000_789, w_000_790, w_000_791, w_000_792, w_000_793, w_000_794, w_000_795, w_000_796, w_000_797, w_000_798, w_000_799, w_000_801, w_000_802, w_000_803, w_000_804, w_000_805, w_000_806, w_000_807, w_000_808, w_000_809, w_000_810, w_000_811, w_000_812, w_000_813, w_000_814, w_000_815, w_000_816, w_000_817, w_000_818, w_000_819, w_000_820, w_000_821, w_000_822, w_000_823, w_000_824, w_000_825, w_000_826, w_000_827, w_000_828, w_000_829, w_000_830, w_000_831, w_000_832, w_000_833, w_000_834, w_000_835, w_000_836, w_000_837, w_000_838, w_000_839, w_000_840, w_000_841, w_000_842, w_000_843, w_000_844, w_000_845, w_000_846, w_000_847, w_000_848, w_000_849, w_000_850, w_000_851, w_000_852, w_000_853, w_000_854, w_000_855, w_000_856, w_000_857, w_000_858, w_000_859, w_000_860, w_000_861, w_000_862, w_000_863, w_000_864, w_000_865, w_000_866, w_000_867, w_000_868, w_000_869, w_000_870, w_000_871, w_000_872, w_000_873, w_000_874, w_000_875, w_000_876, w_000_877, w_000_878, w_000_879, w_000_880, w_000_881, w_000_882, w_000_883, w_000_885, w_000_886, w_000_887, w_000_889, w_000_890, w_000_891, w_000_893, w_000_894, w_000_895, w_000_896, w_000_897, w_000_898, w_000_899, w_000_900, w_000_901, w_000_903, w_000_904, w_000_905, w_000_906, w_000_907, w_000_908, w_000_909, w_000_910, w_000_912, w_000_914, w_000_915, w_000_916, w_000_917, w_000_918, w_000_919, w_000_923, w_000_924, w_000_925, w_000_926, w_000_928, w_000_929, w_000_930, w_000_931, w_000_932, w_000_934, w_000_935, w_000_936, w_000_937, w_000_938, w_000_939, w_000_943, w_000_944, w_000_945, w_000_947, w_000_949, w_000_950, w_000_952, w_000_953, w_000_954, w_000_955, w_000_956, w_000_958, w_000_959, w_000_960, w_000_963, w_000_964, w_000_965, w_000_967, w_000_968, w_000_969, w_000_970, w_000_971, w_000_977, w_000_979, w_000_980, w_000_981, w_000_982, w_000_983;
  wire w_001_000, w_001_001, w_001_002, w_001_003, w_001_004, w_001_005, w_001_006, w_001_007, w_001_008, w_001_009, w_001_010, w_001_011, w_001_012, w_001_013, w_001_014, w_001_015, w_001_016, w_001_017, w_001_018, w_001_019, w_001_020, w_001_021, w_001_022, w_001_023, w_001_024, w_001_026, w_001_027, w_001_028, w_001_029, w_001_030, w_001_031, w_001_032, w_001_033, w_001_034, w_001_035, w_001_036, w_001_037, w_001_038, w_001_039, w_001_040, w_001_041, w_001_042, w_001_043, w_001_044, w_001_046, w_001_047, w_001_048, w_001_050, w_001_051, w_001_052, w_001_053, w_001_054, w_001_055, w_001_056, w_001_057, w_001_058, w_001_059, w_001_060, w_001_061, w_001_062, w_001_063, w_001_064, w_001_065, w_001_066, w_001_068, w_001_069, w_001_070, w_001_071, w_001_072, w_001_073, w_001_074, w_001_075, w_001_076, w_001_077, w_001_078, w_001_079, w_001_080, w_001_081, w_001_082, w_001_083, w_001_084, w_001_085, w_001_086, w_001_087, w_001_088, w_001_089, w_001_090, w_001_091, w_001_092, w_001_093, w_001_094, w_001_095, w_001_096, w_001_097, w_001_098, w_001_099, w_001_100, w_001_101, w_001_102, w_001_103, w_001_104, w_001_107, w_001_108, w_001_109, w_001_110, w_001_111, w_001_112, w_001_114, w_001_115, w_001_118, w_001_119, w_001_120, w_001_121, w_001_122, w_001_123, w_001_124, w_001_125, w_001_126, w_001_127, w_001_128, w_001_129, w_001_130, w_001_131, w_001_132, w_001_133, w_001_134, w_001_136, w_001_138, w_001_139, w_001_140, w_001_141, w_001_142, w_001_143, w_001_144, w_001_146, w_001_147, w_001_148, w_001_149, w_001_150, w_001_151, w_001_152, w_001_154, w_001_155, w_001_156, w_001_157, w_001_158, w_001_160, w_001_163, w_001_164, w_001_165, w_001_167, w_001_168, w_001_170, w_001_171, w_001_173, w_001_174, w_001_175, w_001_176, w_001_177, w_001_178, w_001_179, w_001_180, w_001_181, w_001_182, w_001_184, w_001_186, w_001_187, w_001_188, w_001_189, w_001_190, w_001_191, w_001_192, w_001_193, w_001_194, w_001_195, w_001_196, w_001_197, w_001_198, w_001_199, w_001_201, w_001_202, w_001_203, w_001_205, w_001_206, w_001_207, w_001_210, w_001_211, w_001_213, w_001_214, w_001_215, w_001_216, w_001_217, w_001_218, w_001_219, w_001_221, w_001_222, w_001_224, w_001_225, w_001_226, w_001_228, w_001_229, w_001_230, w_001_231, w_001_233, w_001_234, w_001_235, w_001_236, w_001_237, w_001_238, w_001_239, w_001_241, w_001_243, w_001_244, w_001_245, w_001_246, w_001_247, w_001_249, w_001_250, w_001_251, w_001_253, w_001_255, w_001_256, w_001_257, w_001_259, w_001_260, w_001_261, w_001_263, w_001_264, w_001_265, w_001_266, w_001_267, w_001_268, w_001_269, w_001_270, w_001_271, w_001_274, w_001_275, w_001_276, w_001_277, w_001_278, w_001_279, w_001_280, w_001_281, w_001_282, w_001_283, w_001_284, w_001_285, w_001_286, w_001_287, w_001_288, w_001_290, w_001_291, w_001_293, w_001_295, w_001_296, w_001_297, w_001_299, w_001_300, w_001_301, w_001_303, w_001_304, w_001_305, w_001_306, w_001_307, w_001_308, w_001_310, w_001_311, w_001_312, w_001_313, w_001_314, w_001_316, w_001_317, w_001_318, w_001_319, w_001_320, w_001_321, w_001_322, w_001_323, w_001_324, w_001_325, w_001_326, w_001_327, w_001_328, w_001_329, w_001_330, w_001_332, w_001_333, w_001_334, w_001_335, w_001_339, w_001_340, w_001_341, w_001_342, w_001_343, w_001_345, w_001_346, w_001_347, w_001_348, w_001_349, w_001_350, w_001_351, w_001_352, w_001_353, w_001_354, w_001_355, w_001_356, w_001_357, w_001_358, w_001_360, w_001_361, w_001_362, w_001_363, w_001_365, w_001_366, w_001_367, w_001_368, w_001_369, w_001_370, w_001_371, w_001_374, w_001_375, w_001_376, w_001_377, w_001_378, w_001_380, w_001_381, w_001_382, w_001_385, w_001_387, w_001_388, w_001_390, w_001_391, w_001_393, w_001_394, w_001_395, w_001_396, w_001_397, w_001_398, w_001_399, w_001_400, w_001_401, w_001_402, w_001_403, w_001_405, w_001_406, w_001_407, w_001_408, w_001_409, w_001_410, w_001_411, w_001_412, w_001_414, w_001_415, w_001_416, w_001_417, w_001_418, w_001_420, w_001_422, w_001_423, w_001_425, w_001_426, w_001_427, w_001_428, w_001_429, w_001_430, w_001_432, w_001_433, w_001_435, w_001_436, w_001_437, w_001_438, w_001_439, w_001_440, w_001_441, w_001_442, w_001_443, w_001_445, w_001_446, w_001_447, w_001_448, w_001_449, w_001_451, w_001_452, w_001_453, w_001_454, w_001_455, w_001_456, w_001_457, w_001_458, w_001_459, w_001_460, w_001_462, w_001_464, w_001_465, w_001_466, w_001_467, w_001_468, w_001_469, w_001_470, w_001_471, w_001_472, w_001_473, w_001_474, w_001_475, w_001_476, w_001_477, w_001_478, w_001_479, w_001_480, w_001_481, w_001_482, w_001_483, w_001_484, w_001_485, w_001_486, w_001_487, w_001_488, w_001_489, w_001_490, w_001_491, w_001_492, w_001_493, w_001_494, w_001_495, w_001_496, w_001_497, w_001_498, w_001_500, w_001_501, w_001_502, w_001_503, w_001_504, w_001_505, w_001_506, w_001_507, w_001_508, w_001_509, w_001_510, w_001_512, w_001_513, w_001_514, w_001_515, w_001_516, w_001_518, w_001_519, w_001_521, w_001_522, w_001_523, w_001_524, w_001_525, w_001_527, w_001_528, w_001_529, w_001_531, w_001_532, w_001_533, w_001_534, w_001_537, w_001_538, w_001_539, w_001_540, w_001_542, w_001_543, w_001_544, w_001_546, w_001_547, w_001_548, w_001_549, w_001_551, w_001_553, w_001_555, w_001_557, w_001_558, w_001_559, w_001_561, w_001_562, w_001_564, w_001_565, w_001_566, w_001_567, w_001_568, w_001_569, w_001_570, w_001_571, w_001_572, w_001_573, w_001_574, w_001_575, w_001_576, w_001_577, w_001_578, w_001_579, w_001_580, w_001_581, w_001_582, w_001_584, w_001_585, w_001_586, w_001_587, w_001_589, w_001_590, w_001_591, w_001_592, w_001_593, w_001_595, w_001_597, w_001_598, w_001_599, w_001_600, w_001_601, w_001_602, w_001_603, w_001_604, w_001_605, w_001_606, w_001_607, w_001_608, w_001_609, w_001_611, w_001_612, w_001_613, w_001_614, w_001_615, w_001_616, w_001_617, w_001_618, w_001_619, w_001_620, w_001_622, w_001_623, w_001_624, w_001_625, w_001_627, w_001_629, w_001_631, w_001_632, w_001_633, w_001_634, w_001_635, w_001_636, w_001_637, w_001_638, w_001_639, w_001_640, w_001_641, w_001_642, w_001_644, w_001_645, w_001_647, w_001_650, w_001_652, w_001_653, w_001_654, w_001_655, w_001_656, w_001_657, w_001_658, w_001_659, w_001_661, w_001_662, w_001_663, w_001_665, w_001_666, w_001_667, w_001_669, w_001_670, w_001_671, w_001_672, w_001_673, w_001_674, w_001_675, w_001_677, w_001_678, w_001_679, w_001_680, w_001_681, w_001_683, w_001_684, w_001_685, w_001_686, w_001_687, w_001_688, w_001_689, w_001_690, w_001_691, w_001_692, w_001_694, w_001_695, w_001_696, w_001_697, w_001_698, w_001_700, w_001_701, w_001_702, w_001_703, w_001_704, w_001_706, w_001_707, w_001_709, w_001_710, w_001_711, w_001_712, w_001_713, w_001_714, w_001_716, w_001_717, w_001_718, w_001_719, w_001_720, w_001_721, w_001_722, w_001_723, w_001_725, w_001_726, w_001_727, w_001_728, w_001_729, w_001_730, w_001_731, w_001_732, w_001_734, w_001_737, w_001_738, w_001_742, w_001_743, w_001_744, w_001_745, w_001_746, w_001_748, w_001_750, w_001_751, w_001_752, w_001_753, w_001_755, w_001_756, w_001_757, w_001_759, w_001_760, w_001_761, w_001_762, w_001_763, w_001_764, w_001_765, w_001_766, w_001_767, w_001_768, w_001_769, w_001_770, w_001_771, w_001_772, w_001_773, w_001_774, w_001_775, w_001_777, w_001_778, w_001_779, w_001_780, w_001_782, w_001_783, w_001_784, w_001_785, w_001_786, w_001_787, w_001_788, w_001_789, w_001_790, w_001_791, w_001_792, w_001_793, w_001_794, w_001_796, w_001_797, w_001_798, w_001_799, w_001_800, w_001_801, w_001_802, w_001_803, w_001_804, w_001_805, w_001_807, w_001_809, w_001_810, w_001_811, w_001_812, w_001_813, w_001_814, w_001_816, w_001_817, w_001_818, w_001_819, w_001_820, w_001_822, w_001_824, w_001_825, w_001_826, w_001_827, w_001_828, w_001_829, w_001_832, w_001_834, w_001_835, w_001_838, w_001_839, w_001_842, w_001_843, w_001_844, w_001_845, w_001_846, w_001_847, w_001_848, w_001_850, w_001_852, w_001_853, w_001_854, w_001_856, w_001_857, w_001_858, w_001_859, w_001_860, w_001_861, w_001_864, w_001_865, w_001_866, w_001_867, w_001_868, w_001_870, w_001_871, w_001_872, w_001_874, w_001_876, w_001_878, w_001_880, w_001_881, w_001_882, w_001_883, w_001_884, w_001_885, w_001_886, w_001_888, w_001_889, w_001_890, w_001_892, w_001_893, w_001_894, w_001_895, w_001_896;
  wire w_002_000, w_002_001, w_002_002, w_002_003, w_002_004, w_002_005, w_002_007, w_002_008, w_002_009, w_002_010, w_002_011, w_002_012, w_002_013, w_002_014, w_002_015, w_002_016, w_002_017, w_002_019, w_002_020, w_002_021, w_002_022, w_002_023, w_002_024, w_002_026, w_002_027, w_002_028, w_002_029, w_002_030, w_002_031, w_002_032, w_002_033, w_002_034, w_002_035, w_002_036, w_002_038, w_002_039, w_002_040, w_002_041, w_002_042, w_002_043, w_002_044, w_002_045, w_002_046, w_002_047, w_002_048, w_002_049, w_002_051, w_002_052, w_002_053, w_002_054, w_002_055, w_002_056, w_002_057, w_002_059, w_002_060, w_002_061, w_002_062, w_002_063, w_002_064, w_002_065, w_002_066, w_002_067, w_002_068, w_002_069, w_002_070, w_002_071, w_002_072, w_002_073, w_002_074, w_002_075, w_002_076, w_002_077, w_002_078, w_002_079, w_002_080, w_002_081, w_002_082, w_002_085, w_002_086, w_002_087, w_002_088, w_002_089, w_002_090, w_002_091, w_002_092, w_002_093, w_002_094, w_002_096, w_002_097, w_002_099, w_002_100, w_002_101, w_002_102, w_002_104, w_002_105, w_002_106, w_002_107, w_002_108, w_002_110, w_002_111, w_002_112, w_002_114, w_002_115, w_002_116, w_002_117, w_002_118, w_002_119, w_002_120, w_002_121, w_002_122, w_002_123, w_002_124, w_002_125, w_002_126, w_002_127, w_002_128, w_002_129, w_002_130, w_002_131, w_002_132, w_002_133, w_002_134, w_002_135, w_002_136, w_002_137, w_002_138, w_002_139, w_002_140, w_002_141, w_002_142, w_002_143, w_002_144, w_002_145, w_002_146, w_002_147, w_002_148, w_002_149, w_002_150, w_002_151, w_002_152, w_002_153, w_002_154, w_002_156, w_002_157, w_002_158, w_002_159, w_002_160, w_002_161, w_002_162, w_002_163, w_002_164, w_002_165, w_002_166, w_002_167, w_002_168, w_002_169, w_002_170, w_002_171, w_002_172, w_002_173, w_002_174, w_002_175, w_002_176, w_002_178, w_002_179, w_002_181, w_002_182, w_002_183, w_002_184, w_002_185, w_002_186, w_002_187, w_002_188, w_002_189, w_002_190, w_002_192, w_002_193, w_002_194, w_002_195, w_002_196, w_002_198, w_002_199, w_002_200, w_002_201, w_002_202, w_002_203, w_002_204, w_002_205, w_002_206, w_002_207, w_002_208, w_002_209, w_002_210, w_002_211, w_002_212, w_002_214, w_002_215, w_002_216, w_002_217, w_002_218, w_002_219, w_002_220, w_002_221, w_002_222, w_002_223, w_002_224, w_002_225, w_002_226, w_002_227, w_002_228, w_002_229, w_002_231, w_002_232, w_002_233, w_002_234, w_002_235, w_002_236, w_002_237, w_002_238, w_002_240, w_002_242, w_002_243, w_002_244, w_002_245, w_002_246, w_002_247, w_002_248, w_002_249, w_002_250, w_002_251, w_002_253, w_002_254, w_002_255, w_002_256, w_002_257, w_002_258, w_002_259, w_002_260, w_002_261, w_002_262, w_002_263, w_002_264, w_002_265, w_002_266, w_002_267, w_002_268, w_002_269, w_002_270, w_002_271, w_002_272, w_002_273, w_002_274, w_002_275, w_002_276, w_002_277, w_002_278, w_002_279, w_002_280, w_002_281, w_002_283, w_002_284, w_002_286, w_002_288, w_002_289, w_002_290, w_002_291, w_002_292, w_002_293, w_002_294, w_002_295, w_002_296, w_002_297, w_002_298, w_002_299, w_002_300, w_002_301, w_002_302, w_002_303, w_002_304, w_002_305, w_002_306, w_002_307, w_002_308, w_002_309, w_002_310, w_002_311, w_002_312, w_002_313, w_002_314, w_002_315, w_002_316, w_002_317, w_002_318, w_002_320, w_002_321, w_002_322, w_002_323, w_002_324, w_002_325, w_002_326, w_002_327, w_002_328, w_002_329, w_002_330, w_002_331, w_002_333, w_002_334, w_002_335, w_002_336, w_002_337, w_002_338, w_002_339, w_002_340, w_002_341, w_002_342, w_002_343, w_002_344, w_002_345, w_002_346, w_002_347, w_002_348, w_002_349, w_002_350, w_002_351, w_002_352, w_002_353, w_002_354, w_002_355, w_002_356, w_002_357, w_002_358, w_002_359, w_002_360, w_002_361, w_002_362, w_002_363, w_002_364, w_002_365, w_002_367, w_002_369, w_002_370, w_002_371, w_002_372, w_002_373, w_002_374, w_002_375, w_002_376, w_002_377, w_002_378, w_002_379, w_002_380, w_002_383, w_002_384, w_002_385, w_002_386, w_002_387, w_002_388, w_002_389, w_002_390, w_002_391, w_002_392, w_002_393, w_002_394, w_002_396, w_002_397, w_002_398, w_002_400, w_002_401, w_002_402, w_002_403, w_002_404, w_002_405, w_002_406, w_002_408, w_002_409, w_002_410, w_002_411, w_002_412, w_002_413, w_002_414, w_002_415, w_002_416, w_002_417, w_002_418, w_002_419, w_002_420, w_002_421, w_002_422, w_002_423, w_002_424, w_002_425, w_002_427, w_002_428, w_002_429, w_002_430, w_002_431, w_002_432, w_002_433, w_002_434, w_002_435, w_002_437, w_002_438, w_002_439, w_002_440, w_002_441, w_002_442, w_002_443, w_002_444, w_002_445, w_002_446, w_002_447, w_002_448, w_002_449, w_002_450, w_002_451, w_002_452, w_002_453, w_002_454, w_002_455, w_002_456, w_002_457, w_002_458, w_002_459, w_002_460, w_002_461, w_002_462, w_002_463, w_002_464, w_002_465, w_002_466, w_002_467, w_002_469, w_002_470, w_002_471, w_002_472, w_002_473, w_002_474, w_002_475, w_002_476, w_002_478, w_002_479, w_002_480, w_002_482, w_002_483, w_002_484, w_002_485, w_002_486, w_002_487, w_002_488, w_002_489, w_002_490, w_002_491, w_002_492, w_002_493, w_002_494, w_002_495, w_002_496, w_002_497;
  wire w_003_000, w_003_001, w_003_002, w_003_003, w_003_004, w_003_005, w_003_006, w_003_007, w_003_008, w_003_009, w_003_010, w_003_011, w_003_012, w_003_013, w_003_014, w_003_015, w_003_016, w_003_017, w_003_018, w_003_019, w_003_020, w_003_021, w_003_022, w_003_023, w_003_024, w_003_025, w_003_026, w_003_027, w_003_028, w_003_029, w_003_030, w_003_031, w_003_032, w_003_033, w_003_034, w_003_035, w_003_036, w_003_037, w_003_038, w_003_039, w_003_040, w_003_041, w_003_042, w_003_043, w_003_044, w_003_045, w_003_046, w_003_047, w_003_048, w_003_049, w_003_050, w_003_051, w_003_052, w_003_053, w_003_054, w_003_055, w_003_056, w_003_057, w_003_058, w_003_059, w_003_060, w_003_061, w_003_062, w_003_063, w_003_064, w_003_065, w_003_066, w_003_067, w_003_068, w_003_069, w_003_070, w_003_071, w_003_072, w_003_073, w_003_074, w_003_075, w_003_076, w_003_077, w_003_078, w_003_079, w_003_080, w_003_081, w_003_082, w_003_083, w_003_084, w_003_085, w_003_086, w_003_087, w_003_088, w_003_089, w_003_090, w_003_091, w_003_092, w_003_093, w_003_094, w_003_095, w_003_096, w_003_097, w_003_098, w_003_099, w_003_100, w_003_101, w_003_102, w_003_103, w_003_104, w_003_105, w_003_106, w_003_107, w_003_108, w_003_109, w_003_110, w_003_111, w_003_112, w_003_113, w_003_114, w_003_115, w_003_116, w_003_117, w_003_118, w_003_119, w_003_120, w_003_121, w_003_122, w_003_123, w_003_124, w_003_125, w_003_126, w_003_127, w_003_128, w_003_129, w_003_130, w_003_131, w_003_132, w_003_133, w_003_134, w_003_135, w_003_136, w_003_137, w_003_138, w_003_139, w_003_140, w_003_141, w_003_142, w_003_143, w_003_144, w_003_145, w_003_146, w_003_147, w_003_148, w_003_149, w_003_150, w_003_151, w_003_152, w_003_153, w_003_154, w_003_155, w_003_156, w_003_157, w_003_158, w_003_159, w_003_160, w_003_161, w_003_162, w_003_163, w_003_164, w_003_165, w_003_166, w_003_167, w_003_168, w_003_169, w_003_170, w_003_171, w_003_172, w_003_173, w_003_174, w_003_175, w_003_176, w_003_177, w_003_178, w_003_179, w_003_180, w_003_181, w_003_182, w_003_183, w_003_184, w_003_185, w_003_186, w_003_187, w_003_188, w_003_189, w_003_190, w_003_191, w_003_192, w_003_193, w_003_194, w_003_195, w_003_196, w_003_197, w_003_198, w_003_199, w_003_200, w_003_201, w_003_202, w_003_203, w_003_204, w_003_205, w_003_206, w_003_207, w_003_208, w_003_209, w_003_210, w_003_211, w_003_212, w_003_213, w_003_214, w_003_215, w_003_216, w_003_217, w_003_218, w_003_219, w_003_220, w_003_221, w_003_222, w_003_223, w_003_224, w_003_225;
  wire w_004_000, w_004_001, w_004_002, w_004_003, w_004_004, w_004_005, w_004_006, w_004_007, w_004_008, w_004_009, w_004_010, w_004_011, w_004_012, w_004_013, w_004_014, w_004_015, w_004_016, w_004_017, w_004_018, w_004_019, w_004_020, w_004_021, w_004_022, w_004_023, w_004_024, w_004_025, w_004_026, w_004_027, w_004_028, w_004_029, w_004_030, w_004_031, w_004_032, w_004_033, w_004_034, w_004_035, w_004_036, w_004_037, w_004_038;
  wire w_005_000, w_005_001, w_005_002, w_005_003, w_005_004, w_005_005, w_005_006, w_005_007, w_005_008, w_005_009, w_005_010, w_005_011, w_005_012, w_005_013, w_005_014, w_005_015, w_005_016, w_005_017, w_005_018, w_005_019, w_005_020, w_005_023, w_005_024, w_005_026, w_005_028, w_005_029, w_005_030, w_005_031, w_005_032, w_005_033, w_005_034, w_005_035, w_005_036, w_005_037, w_005_038, w_005_039, w_005_040, w_005_042, w_005_043, w_005_045, w_005_047, w_005_048, w_005_049, w_005_050, w_005_051, w_005_053, w_005_054, w_005_055, w_005_056, w_005_057, w_005_058, w_005_059, w_005_060, w_005_061, w_005_062, w_005_063, w_005_064, w_005_065, w_005_066, w_005_067, w_005_069, w_005_070, w_005_071, w_005_072, w_005_073, w_005_074, w_005_075, w_005_076, w_005_078, w_005_080, w_005_081, w_005_082, w_005_083, w_005_084, w_005_085, w_005_086, w_005_088, w_005_089, w_005_090, w_005_091, w_005_092, w_005_093, w_005_094, w_005_095, w_005_096, w_005_097, w_005_098, w_005_099, w_005_100, w_005_101, w_005_102, w_005_103, w_005_104, w_005_105, w_005_106, w_005_107, w_005_108, w_005_109, w_005_110, w_005_112, w_005_113, w_005_114, w_005_116, w_005_117, w_005_118, w_005_119, w_005_120, w_005_121, w_005_123, w_005_124, w_005_126, w_005_128, w_005_129, w_005_131, w_005_132, w_005_133, w_005_134, w_005_135, w_005_136, w_005_137, w_005_138, w_005_139, w_005_141, w_005_142, w_005_143, w_005_144, w_005_145, w_005_147, w_005_148, w_005_149, w_005_150, w_005_151, w_005_152, w_005_153, w_005_154, w_005_155, w_005_156, w_005_157, w_005_158, w_005_159, w_005_160, w_005_161, w_005_163, w_005_164, w_005_165, w_005_166, w_005_167, w_005_168, w_005_169, w_005_170, w_005_171, w_005_172, w_005_173, w_005_174, w_005_175, w_005_176, w_005_177, w_005_178, w_005_179, w_005_180, w_005_181, w_005_184, w_005_185, w_005_186, w_005_188, w_005_189, w_005_190, w_005_191, w_005_193, w_005_194, w_005_195, w_005_196, w_005_197, w_005_199, w_005_200, w_005_201, w_005_202, w_005_203, w_005_204, w_005_205, w_005_206, w_005_207, w_005_208, w_005_210, w_005_211, w_005_212, w_005_213, w_005_214, w_005_216, w_005_217, w_005_218, w_005_219, w_005_220, w_005_221, w_005_223, w_005_224, w_005_225, w_005_226, w_005_227, w_005_228, w_005_229, w_005_230, w_005_232, w_005_233, w_005_234, w_005_235, w_005_237, w_005_238, w_005_239, w_005_240, w_005_242, w_005_243, w_005_244, w_005_245, w_005_246, w_005_247, w_005_248, w_005_249, w_005_250, w_005_251, w_005_252, w_005_253, w_005_254, w_005_256, w_005_257, w_005_258, w_005_259, w_005_260, w_005_261, w_005_262, w_005_264, w_005_265, w_005_266, w_005_268, w_005_269, w_005_270, w_005_271, w_005_272, w_005_273, w_005_274, w_005_275, w_005_276, w_005_277, w_005_278, w_005_280, w_005_281, w_005_282, w_005_283, w_005_284, w_005_285, w_005_286, w_005_287, w_005_288, w_005_289, w_005_291, w_005_292, w_005_293, w_005_294, w_005_295, w_005_296, w_005_297, w_005_298, w_005_299, w_005_300, w_005_302, w_005_303, w_005_304, w_005_305, w_005_306, w_005_307, w_005_308, w_005_309, w_005_310, w_005_311, w_005_313, w_005_314, w_005_315, w_005_316, w_005_317, w_005_319, w_005_320, w_005_322, w_005_323, w_005_324, w_005_325, w_005_327, w_005_328, w_005_329, w_005_330, w_005_331, w_005_333, w_005_334, w_005_335, w_005_336, w_005_337, w_005_338, w_005_339, w_005_342, w_005_344, w_005_346, w_005_347, w_005_349, w_005_350, w_005_351, w_005_352, w_005_353, w_005_354, w_005_355, w_005_356, w_005_357, w_005_358, w_005_359, w_005_360, w_005_361, w_005_362, w_005_363, w_005_364, w_005_365, w_005_366, w_005_367, w_005_368, w_005_369, w_005_371, w_005_373, w_005_374, w_005_375, w_005_376, w_005_377, w_005_378, w_005_379, w_005_380, w_005_381, w_005_382, w_005_384, w_005_385, w_005_386, w_005_387, w_005_388, w_005_390, w_005_391, w_005_392, w_005_394, w_005_395, w_005_396, w_005_397, w_005_399, w_005_400, w_005_401, w_005_402, w_005_403, w_005_404, w_005_405, w_005_407, w_005_408, w_005_409, w_005_410, w_005_411, w_005_412, w_005_413, w_005_414, w_005_415, w_005_416, w_005_417, w_005_418, w_005_419, w_005_420, w_005_421, w_005_422, w_005_423, w_005_424, w_005_425, w_005_427, w_005_428, w_005_429, w_005_431, w_005_433, w_005_436, w_005_440, w_005_441, w_005_443, w_005_444, w_005_445, w_005_446, w_005_448, w_005_449, w_005_450, w_005_452, w_005_453, w_005_454, w_005_455, w_005_456, w_005_459, w_005_460, w_005_461, w_005_462, w_005_463, w_005_465, w_005_466, w_005_467, w_005_470, w_005_471, w_005_472, w_005_473, w_005_474, w_005_476, w_005_477, w_005_478, w_005_480, w_005_482, w_005_483, w_005_485, w_005_486, w_005_490, w_005_493, w_005_495, w_005_496, w_005_497, w_005_499, w_005_502, w_005_503, w_005_509, w_005_511, w_005_512, w_005_515, w_005_516, w_005_517, w_005_518, w_005_521, w_005_524, w_005_525, w_005_526, w_005_531, w_005_532, w_005_537, w_005_539, w_005_542, w_005_544, w_005_545, w_005_547, w_005_548, w_005_549, w_005_551, w_005_556, w_005_559, w_005_560, w_005_561, w_005_564, w_005_565, w_005_569, w_005_570, w_005_574;
  wire w_006_000, w_006_002, w_006_003, w_006_004, w_006_005, w_006_007, w_006_008, w_006_009, w_006_010, w_006_011, w_006_012, w_006_013, w_006_014, w_006_015, w_006_016, w_006_017, w_006_018, w_006_020, w_006_021, w_006_022, w_006_023, w_006_024, w_006_025, w_006_026, w_006_027, w_006_028, w_006_029, w_006_030, w_006_031, w_006_034, w_006_035, w_006_036, w_006_038, w_006_039, w_006_040, w_006_041, w_006_042, w_006_043, w_006_044, w_006_045, w_006_046, w_006_048, w_006_050, w_006_051, w_006_052, w_006_053, w_006_054, w_006_055, w_006_056, w_006_057, w_006_058, w_006_059, w_006_060, w_006_061, w_006_062, w_006_063, w_006_064, w_006_065, w_006_066, w_006_067, w_006_068, w_006_069, w_006_071, w_006_073, w_006_074, w_006_075, w_006_076, w_006_078, w_006_079, w_006_080, w_006_082, w_006_084, w_006_085, w_006_086, w_006_087, w_006_088, w_006_089, w_006_090, w_006_091, w_006_094, w_006_095, w_006_096, w_006_097, w_006_098, w_006_099, w_006_100, w_006_101, w_006_102, w_006_103, w_006_104, w_006_105, w_006_106, w_006_107, w_006_108, w_006_109, w_006_110, w_006_111, w_006_112, w_006_113, w_006_114, w_006_115, w_006_116, w_006_117, w_006_118, w_006_119, w_006_120, w_006_121, w_006_122, w_006_123, w_006_124, w_006_125, w_006_126, w_006_127, w_006_128, w_006_129, w_006_130, w_006_131, w_006_132, w_006_133, w_006_135, w_006_136, w_006_137, w_006_138, w_006_139, w_006_140, w_006_141, w_006_142, w_006_143, w_006_144, w_006_145, w_006_147, w_006_148, w_006_149, w_006_150, w_006_153, w_006_154, w_006_155, w_006_156, w_006_157, w_006_158, w_006_159, w_006_160, w_006_161, w_006_162, w_006_163, w_006_164, w_006_165, w_006_166, w_006_167, w_006_168, w_006_169, w_006_170, w_006_171, w_006_172, w_006_173, w_006_174, w_006_175, w_006_176, w_006_177, w_006_178, w_006_179, w_006_180, w_006_181, w_006_182, w_006_183, w_006_184, w_006_185, w_006_186, w_006_187, w_006_188, w_006_189, w_006_191, w_006_192, w_006_193, w_006_195, w_006_196, w_006_197, w_006_198, w_006_201, w_006_202, w_006_203, w_006_205, w_006_206, w_006_207, w_006_208, w_006_209, w_006_210, w_006_211, w_006_212, w_006_213, w_006_214, w_006_215, w_006_216, w_006_218, w_006_220, w_006_221, w_006_222, w_006_223, w_006_224, w_006_225, w_006_226, w_006_227, w_006_228, w_006_229, w_006_230, w_006_231, w_006_232, w_006_233, w_006_234, w_006_235, w_006_236, w_006_237, w_006_238, w_006_239, w_006_240, w_006_241, w_006_242, w_006_243, w_006_244, w_006_245, w_006_246, w_006_247, w_006_248, w_006_249, w_006_250, w_006_251, w_006_252, w_006_253, w_006_254, w_006_255, w_006_256, w_006_257, w_006_258, w_006_259, w_006_260, w_006_261, w_006_262, w_006_263, w_006_264, w_006_265, w_006_266, w_006_267, w_006_268, w_006_270, w_006_271, w_006_272, w_006_273, w_006_274, w_006_275, w_006_276, w_006_277, w_006_278, w_006_279, w_006_280, w_006_281, w_006_282, w_006_283, w_006_284, w_006_285, w_006_286, w_006_287, w_006_288, w_006_289, w_006_290, w_006_291, w_006_292, w_006_293, w_006_294, w_006_295, w_006_296, w_006_297, w_006_298, w_006_299, w_006_300, w_006_302, w_006_303, w_006_304, w_006_305, w_006_306, w_006_307, w_006_308, w_006_309, w_006_310, w_006_311, w_006_312, w_006_313, w_006_314, w_006_315, w_006_316, w_006_317, w_006_318, w_006_319, w_006_320, w_006_321, w_006_322, w_006_323, w_006_324, w_006_325, w_006_326, w_006_327, w_006_328, w_006_329, w_006_330, w_006_331, w_006_332;
  wire w_007_000, w_007_001, w_007_002, w_007_004, w_007_005, w_007_007, w_007_010, w_007_011, w_007_012, w_007_013, w_007_014, w_007_015, w_007_017, w_007_018, w_007_019, w_007_020, w_007_021, w_007_023, w_007_024, w_007_026, w_007_027, w_007_029, w_007_030, w_007_031, w_007_032, w_007_033, w_007_035, w_007_038, w_007_039, w_007_040, w_007_041, w_007_042, w_007_043, w_007_044, w_007_045, w_007_046, w_007_047, w_007_048, w_007_049, w_007_050, w_007_052, w_007_053, w_007_054, w_007_055, w_007_057, w_007_058, w_007_060, w_007_062, w_007_063, w_007_064, w_007_065, w_007_067, w_007_068, w_007_069, w_007_070, w_007_072, w_007_073, w_007_074, w_007_075, w_007_076, w_007_077, w_007_078, w_007_079, w_007_080, w_007_081, w_007_082, w_007_083, w_007_085, w_007_088, w_007_089, w_007_091, w_007_092, w_007_093, w_007_094, w_007_095, w_007_097, w_007_098, w_007_099, w_007_100, w_007_101, w_007_103, w_007_105, w_007_107, w_007_108, w_007_109, w_007_110, w_007_111, w_007_113, w_007_115, w_007_116, w_007_117, w_007_119, w_007_121, w_007_122, w_007_123, w_007_127, w_007_128, w_007_129, w_007_130, w_007_131, w_007_132, w_007_134, w_007_135, w_007_136, w_007_137, w_007_138, w_007_139, w_007_140, w_007_142, w_007_143, w_007_144, w_007_145, w_007_147, w_007_148, w_007_149, w_007_150, w_007_151, w_007_152, w_007_153, w_007_155, w_007_156, w_007_157, w_007_158, w_007_159, w_007_160, w_007_161, w_007_162, w_007_163, w_007_164, w_007_165, w_007_166, w_007_167, w_007_168, w_007_169, w_007_171, w_007_173, w_007_175, w_007_177, w_007_179, w_007_182, w_007_183, w_007_185, w_007_186, w_007_187, w_007_188, w_007_189, w_007_190, w_007_192, w_007_193, w_007_194, w_007_195, w_007_196, w_007_198, w_007_199, w_007_200, w_007_201, w_007_202, w_007_203, w_007_204, w_007_205, w_007_207, w_007_208, w_007_209, w_007_210, w_007_212, w_007_213, w_007_214, w_007_215, w_007_216, w_007_217, w_007_218, w_007_219, w_007_220, w_007_221, w_007_222, w_007_223, w_007_224, w_007_228, w_007_229, w_007_230, w_007_232, w_007_233, w_007_234, w_007_235, w_007_236, w_007_237, w_007_238, w_007_239, w_007_240, w_007_243, w_007_244, w_007_245, w_007_246, w_007_247, w_007_248, w_007_249, w_007_250, w_007_251, w_007_252, w_007_253, w_007_254, w_007_255, w_007_256, w_007_257, w_007_259, w_007_260, w_007_261, w_007_262, w_007_264, w_007_265, w_007_266, w_007_267, w_007_268, w_007_269, w_007_272, w_007_273, w_007_275, w_007_276, w_007_277, w_007_278, w_007_280, w_007_281, w_007_282, w_007_283, w_007_284, w_007_286, w_007_287, w_007_288, w_007_293, w_007_294, w_007_295, w_007_296, w_007_297, w_007_298, w_007_299, w_007_301, w_007_302, w_007_303, w_007_304, w_007_306, w_007_307, w_007_308, w_007_309, w_007_310, w_007_311, w_007_313, w_007_314, w_007_315, w_007_316, w_007_317, w_007_318, w_007_319, w_007_321, w_007_322, w_007_324, w_007_327, w_007_328, w_007_329, w_007_331, w_007_332, w_007_333, w_007_335, w_007_336, w_007_337, w_007_338, w_007_340, w_007_341, w_007_342, w_007_343, w_007_345, w_007_346, w_007_347, w_007_348, w_007_349, w_007_350, w_007_351, w_007_352, w_007_353, w_007_356, w_007_357, w_007_358, w_007_359, w_007_360, w_007_361, w_007_362, w_007_363, w_007_364, w_007_365, w_007_366, w_007_367, w_007_369, w_007_371, w_007_373, w_007_374, w_007_375, w_007_376, w_007_377, w_007_378, w_007_381, w_007_383, w_007_384, w_007_385, w_007_386, w_007_387, w_007_388, w_007_390, w_007_391, w_007_392, w_007_393, w_007_394, w_007_395, w_007_398, w_007_399, w_007_400, w_007_401, w_007_402, w_007_403, w_007_404, w_007_405, w_007_406, w_007_407, w_007_408, w_007_409, w_007_411, w_007_413, w_007_414, w_007_415, w_007_416, w_007_417, w_007_418, w_007_419, w_007_420, w_007_421, w_007_422, w_007_423, w_007_425, w_007_426, w_007_427, w_007_428, w_007_430, w_007_431, w_007_432, w_007_433, w_007_435, w_007_436, w_007_437, w_007_438, w_007_446, w_007_447, w_007_448, w_007_450, w_007_451, w_007_454, w_007_456, w_007_459, w_007_460, w_007_463, w_007_464, w_007_472, w_007_475, w_007_476, w_007_484, w_007_485, w_007_487, w_007_488, w_007_489, w_007_491, w_007_495, w_007_497, w_007_499, w_007_500, w_007_501, w_007_504, w_007_507, w_007_509, w_007_511, w_007_512, w_007_513, w_007_515, w_007_517, w_007_524, w_007_526, w_007_532, w_007_535, w_007_537, w_007_538, w_007_539, w_007_540, w_007_543, w_007_546, w_007_549, w_007_551, w_007_552, w_007_553, w_007_554, w_007_556, w_007_558, w_007_559;
  wire w_008_001, w_008_002, w_008_004, w_008_006, w_008_007, w_008_010, w_008_012, w_008_013, w_008_015, w_008_016, w_008_017, w_008_018, w_008_021, w_008_022, w_008_023, w_008_024, w_008_025, w_008_026, w_008_028, w_008_030, w_008_033, w_008_034, w_008_035, w_008_036, w_008_037, w_008_038, w_008_043, w_008_044, w_008_046, w_008_049, w_008_050, w_008_051, w_008_053, w_008_054, w_008_056, w_008_061, w_008_064, w_008_067, w_008_069, w_008_071, w_008_072, w_008_073, w_008_074, w_008_077, w_008_078, w_008_079, w_008_084, w_008_086, w_008_088, w_008_090, w_008_092, w_008_096, w_008_097, w_008_100, w_008_102, w_008_104, w_008_107, w_008_108, w_008_109, w_008_116, w_008_118, w_008_122, w_008_126, w_008_129, w_008_130, w_008_131, w_008_133, w_008_134, w_008_135, w_008_138, w_008_142, w_008_143, w_008_145, w_008_147, w_008_149, w_008_154, w_008_155, w_008_156, w_008_158, w_008_161, w_008_163, w_008_167, w_008_168, w_008_169, w_008_170, w_008_172, w_008_174, w_008_176, w_008_178, w_008_179, w_008_182, w_008_184, w_008_186, w_008_187, w_008_188, w_008_191, w_008_192, w_008_194, w_008_200, w_008_202, w_008_209, w_008_210, w_008_211, w_008_213, w_008_215, w_008_216, w_008_217, w_008_218, w_008_220, w_008_222, w_008_225, w_008_226, w_008_227, w_008_230, w_008_231, w_008_232, w_008_234, w_008_235, w_008_236, w_008_237, w_008_241, w_008_242, w_008_244, w_008_246, w_008_247, w_008_251, w_008_252, w_008_253, w_008_254, w_008_257, w_008_259, w_008_260, w_008_261, w_008_263, w_008_264, w_008_267, w_008_268, w_008_269, w_008_271, w_008_272, w_008_275, w_008_276, w_008_277, w_008_278, w_008_279, w_008_280, w_008_281, w_008_282, w_008_283, w_008_285, w_008_288, w_008_289, w_008_294, w_008_297, w_008_299, w_008_300, w_008_302, w_008_303, w_008_304, w_008_305, w_008_306, w_008_310, w_008_314, w_008_318, w_008_319, w_008_325, w_008_326, w_008_327, w_008_328, w_008_331, w_008_332, w_008_333, w_008_335, w_008_340, w_008_343, w_008_344, w_008_346, w_008_347, w_008_348, w_008_349, w_008_354, w_008_355, w_008_356, w_008_358, w_008_361, w_008_365, w_008_373, w_008_374, w_008_377, w_008_379, w_008_383, w_008_384, w_008_386, w_008_387, w_008_388, w_008_389, w_008_392, w_008_396, w_008_397, w_008_398, w_008_400, w_008_401, w_008_405, w_008_406, w_008_407, w_008_408, w_008_409, w_008_411, w_008_414, w_008_423, w_008_425, w_008_428, w_008_432, w_008_434, w_008_435, w_008_437, w_008_442, w_008_446, w_008_447, w_008_448, w_008_450, w_008_458, w_008_459, w_008_461, w_008_462, w_008_466, w_008_473, w_008_474, w_008_477, w_008_478, w_008_480, w_008_482, w_008_484, w_008_485, w_008_486, w_008_487, w_008_488, w_008_490, w_008_491, w_008_494, w_008_496, w_008_497, w_008_499, w_008_501, w_008_503, w_008_505, w_008_510, w_008_514, w_008_515, w_008_517, w_008_520, w_008_527, w_008_528, w_008_529, w_008_534, w_008_542, w_008_545, w_008_548, w_008_553, w_008_555, w_008_557, w_008_559, w_008_560, w_008_562, w_008_565, w_008_566, w_008_567, w_008_568, w_008_574, w_008_575, w_008_578, w_008_581, w_008_582, w_008_585, w_008_586, w_008_588, w_008_591, w_008_595, w_008_596, w_008_597, w_008_598, w_008_599, w_008_600, w_008_601, w_008_604, w_008_608, w_008_609, w_008_610, w_008_611, w_008_613, w_008_615, w_008_616, w_008_619, w_008_620, w_008_621, w_008_629, w_008_631, w_008_632, w_008_633, w_008_636, w_008_638, w_008_642, w_008_645, w_008_646, w_008_647, w_008_651, w_008_652, w_008_654, w_008_655, w_008_656, w_008_658, w_008_661, w_008_662, w_008_665, w_008_666, w_008_668, w_008_669, w_008_670, w_008_671, w_008_672, w_008_674, w_008_675, w_008_676, w_008_677, w_008_678, w_008_679, w_008_680, w_008_681, w_008_682, w_008_684, w_008_685, w_008_689, w_008_690, w_008_692, w_008_694, w_008_702, w_008_703, w_008_704, w_008_706, w_008_707, w_008_708, w_008_712, w_008_714, w_008_717, w_008_718, w_008_720, w_008_722, w_008_727, w_008_734, w_008_735, w_008_737, w_008_739, w_008_746, w_008_747, w_008_748, w_008_749, w_008_750, w_008_756, w_008_758, w_008_759, w_008_760, w_008_761, w_008_764, w_008_765, w_008_768, w_008_769, w_008_770, w_008_771, w_008_772, w_008_773, w_008_779, w_008_780, w_008_785, w_008_790, w_008_792, w_008_793, w_008_794, w_008_795, w_008_803, w_008_804, w_008_806, w_008_808, w_008_810, w_008_813, w_008_814, w_008_815, w_008_820, w_008_822, w_008_824, w_008_826, w_008_827, w_008_828, w_008_829, w_008_830, w_008_832, w_008_835, w_008_836, w_008_837, w_008_840, w_008_848, w_008_850, w_008_853, w_008_857, w_008_861, w_008_862, w_008_863, w_008_864, w_008_866, w_008_874, w_008_877, w_008_878, w_008_879, w_008_880, w_008_881, w_008_882, w_008_884, w_008_885, w_008_886, w_008_888, w_008_889, w_008_890, w_008_891, w_008_892, w_008_893, w_008_894, w_008_896, w_008_897, w_008_898, w_008_899, w_008_900, w_008_906, w_008_908, w_008_910, w_008_912, w_008_914, w_008_917, w_008_918, w_008_919, w_008_920, w_008_921, w_008_922, w_008_923, w_008_925, w_008_926, w_008_927, w_008_930, w_008_931, w_008_933, w_008_935, w_008_936, w_008_939, w_008_941, w_008_943, w_008_947, w_008_949, w_008_951, w_008_952, w_008_953, w_008_955, w_008_959;
  wire w_009_000, w_009_001, w_009_002, w_009_003, w_009_004, w_009_005, w_009_006, w_009_007, w_009_008, w_009_009, w_009_010, w_009_011, w_009_012, w_009_013, w_009_014, w_009_015, w_009_016, w_009_017, w_009_018, w_009_019, w_009_020, w_009_021, w_009_022, w_009_023, w_009_024, w_009_025, w_009_026, w_009_027, w_009_028, w_009_029, w_009_030, w_009_031, w_009_032, w_009_033, w_009_034, w_009_035, w_009_036, w_009_037, w_009_038, w_009_039, w_009_040, w_009_041, w_009_042, w_009_043, w_009_044, w_009_045, w_009_046, w_009_047, w_009_048, w_009_049, w_009_050, w_009_051, w_009_052, w_009_053, w_009_054, w_009_055, w_009_056, w_009_057, w_009_058, w_009_059, w_009_060, w_009_061, w_009_062, w_009_063, w_009_064, w_009_065, w_009_066, w_009_067, w_009_068;
  wire w_010_002, w_010_003, w_010_004, w_010_005, w_010_006, w_010_007, w_010_008, w_010_009, w_010_010, w_010_011, w_010_012, w_010_013, w_010_014, w_010_015, w_010_016, w_010_017, w_010_018, w_010_020, w_010_021, w_010_023, w_010_025, w_010_027, w_010_029, w_010_031, w_010_033, w_010_034, w_010_035, w_010_037, w_010_039, w_010_040, w_010_042, w_010_043, w_010_044, w_010_047, w_010_049, w_010_050, w_010_052, w_010_053, w_010_054, w_010_057, w_010_058, w_010_059, w_010_060, w_010_061, w_010_063, w_010_065, w_010_067, w_010_070, w_010_072, w_010_073, w_010_074, w_010_077, w_010_078, w_010_079, w_010_080, w_010_081, w_010_082, w_010_084, w_010_085, w_010_086, w_010_087, w_010_088, w_010_090, w_010_091, w_010_092, w_010_094, w_010_095, w_010_097, w_010_099, w_010_103, w_010_107, w_010_109, w_010_110, w_010_111, w_010_113, w_010_114, w_010_115, w_010_116, w_010_117, w_010_118, w_010_120, w_010_121, w_010_122, w_010_123, w_010_125, w_010_127, w_010_128, w_010_130, w_010_132, w_010_134, w_010_136, w_010_137, w_010_139, w_010_140, w_010_141, w_010_143, w_010_144, w_010_145, w_010_146, w_010_147, w_010_148, w_010_152, w_010_155, w_010_156, w_010_157, w_010_158, w_010_159, w_010_160, w_010_161, w_010_162, w_010_163, w_010_164, w_010_165, w_010_166, w_010_170, w_010_171, w_010_176, w_010_177, w_010_178, w_010_181, w_010_184, w_010_190, w_010_192, w_010_193, w_010_196, w_010_197, w_010_198, w_010_200, w_010_204, w_010_205, w_010_208, w_010_210, w_010_211, w_010_212, w_010_218, w_010_220, w_010_222, w_010_223, w_010_225, w_010_226, w_010_229, w_010_232, w_010_234, w_010_236, w_010_240, w_010_246, w_010_247, w_010_249, w_010_251, w_010_253, w_010_255, w_010_256, w_010_257, w_010_259, w_010_260, w_010_261, w_010_264, w_010_265, w_010_267, w_010_269, w_010_272, w_010_278, w_010_279, w_010_280, w_010_281, w_010_294, w_010_295, w_010_296, w_010_297, w_010_298, w_010_302, w_010_304, w_010_307, w_010_310, w_010_311, w_010_312, w_010_313, w_010_315, w_010_316, w_010_321, w_010_323, w_010_326, w_010_329, w_010_330, w_010_332, w_010_334, w_010_335, w_010_338, w_010_339, w_010_340, w_010_344, w_010_346, w_010_349, w_010_353, w_010_358, w_010_359, w_010_365, w_010_366, w_010_367, w_010_370, w_010_374, w_010_376, w_010_377, w_010_378, w_010_379, w_010_381, w_010_385, w_010_387, w_010_388, w_010_389, w_010_391, w_010_392, w_010_396, w_010_397, w_010_401, w_010_403, w_010_404, w_010_406, w_010_407, w_010_409, w_010_413, w_010_414, w_010_415, w_010_416, w_010_417, w_010_420, w_010_424, w_010_426, w_010_430, w_010_432, w_010_436, w_010_438, w_010_440, w_010_445, w_010_446, w_010_448, w_010_449, w_010_450, w_010_452, w_010_453, w_010_456, w_010_459, w_010_461, w_010_463, w_010_465, w_010_466, w_010_467, w_010_468, w_010_473, w_010_474, w_010_475, w_010_479, w_010_480, w_010_484, w_010_486, w_010_488, w_010_491, w_010_492, w_010_494, w_010_499, w_010_501, w_010_504, w_010_506, w_010_507, w_010_511, w_010_514, w_010_518, w_010_519, w_010_520, w_010_522, w_010_523, w_010_525, w_010_526, w_010_528, w_010_530, w_010_531, w_010_536, w_010_539, w_010_540, w_010_542, w_010_543, w_010_547, w_010_548, w_010_549, w_010_550, w_010_551, w_010_557, w_010_562, w_010_565, w_010_567, w_010_570, w_010_571, w_010_573, w_010_575, w_010_576, w_010_579, w_010_580, w_010_583, w_010_586, w_010_588, w_010_590, w_010_591, w_010_592, w_010_595, w_010_596, w_010_597, w_010_598, w_010_599, w_010_601, w_010_606, w_010_607, w_010_609, w_010_612, w_010_613, w_010_614, w_010_615, w_010_618, w_010_622, w_010_623, w_010_624, w_010_626, w_010_627, w_010_628, w_010_632, w_010_633, w_010_637, w_010_640, w_010_641, w_010_642, w_010_643, w_010_645, w_010_646, w_010_649, w_010_650, w_010_652, w_010_653, w_010_654, w_010_657, w_010_659, w_010_665, w_010_667, w_010_670, w_010_680, w_010_683, w_010_685, w_010_688, w_010_689, w_010_693, w_010_694, w_010_697, w_010_698, w_010_699, w_010_703, w_010_706, w_010_707, w_010_708, w_010_712, w_010_714, w_010_715, w_010_716, w_010_717, w_010_718, w_010_719, w_010_729, w_010_730, w_010_734, w_010_736, w_010_738, w_010_740, w_010_741, w_010_744, w_010_746, w_010_747, w_010_749, w_010_751, w_010_754, w_010_756, w_010_757, w_010_760, w_010_766, w_010_767, w_010_768, w_010_771, w_010_772, w_010_773, w_010_776, w_010_777, w_010_779, w_010_780, w_010_781, w_010_785, w_010_790, w_010_793, w_010_795, w_010_798, w_010_802, w_010_804, w_010_805, w_010_806, w_010_807, w_010_809, w_010_810, w_010_812, w_010_813, w_010_815, w_010_817, w_010_819, w_010_820, w_010_821, w_010_822, w_010_825, w_010_827, w_010_831, w_010_833, w_010_834;
  wire w_011_000, w_011_001, w_011_003, w_011_004, w_011_006, w_011_007, w_011_008, w_011_009, w_011_010, w_011_011, w_011_013, w_011_014, w_011_016, w_011_017, w_011_018, w_011_020, w_011_022, w_011_023, w_011_025, w_011_026, w_011_029, w_011_030, w_011_031, w_011_032, w_011_033, w_011_034, w_011_037, w_011_039, w_011_040, w_011_041, w_011_042, w_011_043, w_011_044, w_011_045, w_011_046, w_011_047, w_011_049, w_011_050, w_011_053, w_011_056, w_011_057, w_011_058, w_011_059, w_011_062, w_011_063, w_011_064, w_011_065, w_011_066, w_011_067, w_011_068, w_011_069, w_011_071, w_011_072, w_011_075, w_011_078, w_011_079, w_011_082, w_011_084, w_011_087, w_011_088, w_011_090, w_011_091, w_011_092, w_011_093, w_011_094, w_011_096, w_011_097, w_011_101, w_011_102, w_011_103, w_011_106, w_011_107, w_011_109, w_011_110, w_011_111, w_011_112, w_011_114, w_011_118, w_011_120, w_011_121, w_011_122, w_011_125, w_011_126, w_011_127, w_011_129, w_011_130, w_011_131, w_011_133, w_011_135, w_011_136, w_011_137, w_011_138, w_011_140, w_011_141, w_011_142, w_011_143, w_011_144, w_011_146, w_011_150, w_011_153, w_011_154, w_011_155, w_011_156, w_011_157, w_011_158, w_011_159, w_011_160, w_011_161, w_011_162, w_011_163, w_011_164, w_011_167, w_011_168, w_011_170, w_011_171, w_011_172, w_011_173, w_011_175, w_011_176, w_011_177, w_011_178, w_011_180, w_011_182, w_011_183, w_011_186, w_011_187, w_011_190, w_011_191, w_011_192, w_011_193, w_011_195, w_011_198, w_011_200, w_011_201, w_011_203, w_011_205, w_011_206, w_011_209, w_011_211, w_011_212, w_011_213, w_011_216, w_011_217, w_011_221, w_011_222, w_011_223, w_011_224, w_011_225, w_011_226, w_011_227, w_011_229, w_011_231, w_011_232, w_011_233, w_011_236, w_011_239, w_011_240, w_011_241, w_011_242, w_011_243, w_011_245, w_011_246, w_011_247, w_011_250, w_011_251, w_011_253, w_011_254, w_011_257, w_011_258, w_011_259, w_011_260, w_011_261, w_011_262, w_011_263, w_011_264, w_011_265, w_011_266, w_011_267, w_011_268, w_011_269, w_011_271, w_011_272, w_011_273, w_011_274, w_011_276, w_011_277, w_011_278, w_011_280, w_011_281, w_011_282, w_011_283, w_011_287, w_011_288, w_011_291, w_011_292, w_011_295, w_011_297, w_011_299, w_011_304, w_011_305, w_011_306, w_011_308, w_011_309, w_011_310, w_011_312, w_011_314, w_011_315, w_011_317, w_011_318, w_011_322, w_011_327, w_011_335, w_011_336, w_011_337, w_011_339, w_011_340, w_011_343, w_011_347, w_011_349, w_011_351, w_011_353, w_011_355, w_011_356, w_011_359, w_011_360, w_011_361, w_011_367, w_011_369, w_011_370, w_011_371, w_011_372, w_011_373, w_011_374, w_011_376, w_011_380, w_011_387, w_011_394, w_011_395, w_011_396, w_011_398, w_011_399, w_011_402, w_011_403, w_011_406, w_011_407, w_011_409, w_011_412, w_011_415, w_011_419, w_011_420, w_011_422, w_011_423, w_011_426, w_011_430, w_011_433, w_011_434, w_011_437, w_011_449, w_011_456, w_011_457, w_011_458, w_011_459, w_011_460, w_011_463, w_011_464, w_011_467, w_011_474, w_011_476, w_011_477, w_011_478, w_011_485, w_011_486, w_011_492, w_011_495, w_011_496, w_011_500, w_011_501, w_011_502, w_011_503, w_011_504, w_011_505, w_011_510, w_011_511, w_011_513, w_011_514, w_011_520, w_011_523, w_011_525, w_011_526, w_011_530, w_011_534, w_011_535, w_011_537, w_011_540, w_011_543, w_011_546, w_011_548, w_011_553, w_011_556, w_011_558, w_011_560, w_011_564, w_011_565, w_011_566, w_011_568, w_011_569, w_011_577, w_011_578, w_011_581, w_011_583, w_011_584, w_011_587, w_011_596, w_011_601, w_011_603, w_011_604, w_011_606, w_011_607, w_011_608, w_011_610, w_011_615, w_011_618, w_011_619, w_011_622, w_011_624, w_011_628, w_011_631, w_011_635, w_011_637, w_011_644, w_011_645, w_011_646, w_011_648, w_011_649, w_011_650, w_011_652, w_011_655, w_011_656, w_011_657, w_011_659, w_011_661, w_011_662, w_011_666, w_011_667, w_011_669, w_011_673, w_011_675, w_011_678, w_011_679;
  wire w_012_002, w_012_003, w_012_006, w_012_007, w_012_008, w_012_010, w_012_011, w_012_012, w_012_017, w_012_018, w_012_022, w_012_023, w_012_025, w_012_026, w_012_027, w_012_028, w_012_030, w_012_037, w_012_038, w_012_039, w_012_040, w_012_042, w_012_043, w_012_044, w_012_045, w_012_048, w_012_050, w_012_054, w_012_055, w_012_056, w_012_057, w_012_058, w_012_061, w_012_062, w_012_063, w_012_066, w_012_068, w_012_069, w_012_070, w_012_071, w_012_072, w_012_076, w_012_077, w_012_080, w_012_083, w_012_084, w_012_085, w_012_086, w_012_088, w_012_089, w_012_091, w_012_092, w_012_093, w_012_096, w_012_098, w_012_099, w_012_101, w_012_102, w_012_104, w_012_105, w_012_106, w_012_107, w_012_108, w_012_109, w_012_110, w_012_112, w_012_113, w_012_114, w_012_115, w_012_116, w_012_117, w_012_121, w_012_124, w_012_126, w_012_127, w_012_128, w_012_130, w_012_133, w_012_134, w_012_136, w_012_137, w_012_138, w_012_139, w_012_142, w_012_143, w_012_149, w_012_151, w_012_154, w_012_155, w_012_157, w_012_158, w_012_159, w_012_161, w_012_162, w_012_163, w_012_165, w_012_166, w_012_167, w_012_169, w_012_170, w_012_171, w_012_172, w_012_173, w_012_174, w_012_177, w_012_178, w_012_179, w_012_182, w_012_183, w_012_184, w_012_185, w_012_186, w_012_188, w_012_190, w_012_191, w_012_192, w_012_193, w_012_195, w_012_197, w_012_199, w_012_203, w_012_204, w_012_206, w_012_207, w_012_209, w_012_211, w_012_212, w_012_216, w_012_217, w_012_218, w_012_220, w_012_221, w_012_223, w_012_224, w_012_226, w_012_231, w_012_236, w_012_237, w_012_238, w_012_242, w_012_244, w_012_245, w_012_246, w_012_248, w_012_249, w_012_252, w_012_253, w_012_256, w_012_257, w_012_260, w_012_262, w_012_263, w_012_265, w_012_266, w_012_268, w_012_269, w_012_270, w_012_271, w_012_272, w_012_273, w_012_275, w_012_276, w_012_279, w_012_280, w_012_281, w_012_284, w_012_287, w_012_288, w_012_289, w_012_290, w_012_297, w_012_299, w_012_300, w_012_301, w_012_303, w_012_304, w_012_306, w_012_307, w_012_308, w_012_312, w_012_314, w_012_316, w_012_317, w_012_318, w_012_321, w_012_322, w_012_323, w_012_324, w_012_325, w_012_327, w_012_329, w_012_330, w_012_331, w_012_332, w_012_336, w_012_337, w_012_338, w_012_339, w_012_341, w_012_343, w_012_344, w_012_345, w_012_349, w_012_350, w_012_352, w_012_357, w_012_359, w_012_361, w_012_365, w_012_367, w_012_369, w_012_371, w_012_373, w_012_374, w_012_375, w_012_378, w_012_382, w_012_383, w_012_384, w_012_385, w_012_387, w_012_388, w_012_389, w_012_392, w_012_395, w_012_396, w_012_397, w_012_399, w_012_400, w_012_403, w_012_405, w_012_406, w_012_409, w_012_410, w_012_411, w_012_413, w_012_414, w_012_415, w_012_416, w_012_419, w_012_420, w_012_422, w_012_423, w_012_424, w_012_425, w_012_426, w_012_427, w_012_428, w_012_429, w_012_431, w_012_432, w_012_434, w_012_435, w_012_436, w_012_437, w_012_438, w_012_439, w_012_441, w_012_442, w_012_446, w_012_447, w_012_451, w_012_453, w_012_456, w_012_458, w_012_459, w_012_460, w_012_462, w_012_463, w_012_465, w_012_469, w_012_470, w_012_471, w_012_472, w_012_474, w_012_477, w_012_478, w_012_488, w_012_491, w_012_493, w_012_494, w_012_500, w_012_504, w_012_511, w_012_516, w_012_519, w_012_523, w_012_524, w_012_525, w_012_531, w_012_533, w_012_535, w_012_538, w_012_539, w_012_543, w_012_544, w_012_551;
  wire w_013_002, w_013_003, w_013_004, w_013_005, w_013_006, w_013_009, w_013_010, w_013_011, w_013_012, w_013_013, w_013_014, w_013_016, w_013_017, w_013_019, w_013_020, w_013_022, w_013_025, w_013_026, w_013_028, w_013_029, w_013_030, w_013_031, w_013_032, w_013_033, w_013_034, w_013_035, w_013_037, w_013_039, w_013_042, w_013_044, w_013_045, w_013_047, w_013_048, w_013_050, w_013_052, w_013_054, w_013_057, w_013_058, w_013_060, w_013_064, w_013_065, w_013_067, w_013_073, w_013_074, w_013_075, w_013_077, w_013_078, w_013_079, w_013_080, w_013_081, w_013_086, w_013_090, w_013_096, w_013_097, w_013_098, w_013_099, w_013_100, w_013_102, w_013_104, w_013_105, w_013_106, w_013_107, w_013_108, w_013_112, w_013_114, w_013_116, w_013_119, w_013_120, w_013_121, w_013_123, w_013_126, w_013_127, w_013_128, w_013_129, w_013_133, w_013_136, w_013_139, w_013_140, w_013_142, w_013_143, w_013_146, w_013_147, w_013_148, w_013_150, w_013_152, w_013_154, w_013_157, w_013_158, w_013_159, w_013_160, w_013_161, w_013_164, w_013_165, w_013_167, w_013_170, w_013_171, w_013_172, w_013_174, w_013_175, w_013_176, w_013_177, w_013_178, w_013_180, w_013_181, w_013_184, w_013_186, w_013_187, w_013_188, w_013_189, w_013_191, w_013_192, w_013_194, w_013_197, w_013_198, w_013_202, w_013_203, w_013_204, w_013_207, w_013_208, w_013_209, w_013_210, w_013_213, w_013_219, w_013_220, w_013_223, w_013_224, w_013_228, w_013_233, w_013_235, w_013_237, w_013_238, w_013_239, w_013_240, w_013_241, w_013_242, w_013_243, w_013_244, w_013_249, w_013_251, w_013_252, w_013_253, w_013_254, w_013_258, w_013_259, w_013_260, w_013_261, w_013_263, w_013_264, w_013_265, w_013_267, w_013_268, w_013_271, w_013_272, w_013_273, w_013_274, w_013_276, w_013_277, w_013_278, w_013_279, w_013_280, w_013_281, w_013_282, w_013_285, w_013_286, w_013_288, w_013_290, w_013_291, w_013_292, w_013_297, w_013_298, w_013_299, w_013_300, w_013_301, w_013_302, w_013_303, w_013_305, w_013_307, w_013_308, w_013_309, w_013_310, w_013_311, w_013_312, w_013_313, w_013_315, w_013_316, w_013_317, w_013_319, w_013_320, w_013_321, w_013_324, w_013_325, w_013_326, w_013_327, w_013_328, w_013_329, w_013_330, w_013_333, w_013_335, w_013_338, w_013_339, w_013_350, w_013_353, w_013_355, w_013_357, w_013_362, w_013_363, w_013_365, w_013_368, w_013_370, w_013_372, w_013_373, w_013_375, w_013_376, w_013_377, w_013_379, w_013_381, w_013_382, w_013_384, w_013_386, w_013_387, w_013_389, w_013_391, w_013_392, w_013_396, w_013_399, w_013_404, w_013_405, w_013_406, w_013_407, w_013_409, w_013_412, w_013_415, w_013_416, w_013_417, w_013_418, w_013_419, w_013_420, w_013_421, w_013_422, w_013_423, w_013_424, w_013_426, w_013_428, w_013_430, w_013_431, w_013_433, w_013_434, w_013_437, w_013_441, w_013_442, w_013_444, w_013_445, w_013_446, w_013_448, w_013_449, w_013_450, w_013_451, w_013_452, w_013_453, w_013_455, w_013_457, w_013_458, w_013_459, w_013_462, w_013_463, w_013_465, w_013_466, w_013_469, w_013_470, w_013_471, w_013_475, w_013_477, w_013_478, w_013_479, w_013_480, w_013_481, w_013_485, w_013_486, w_013_487, w_013_488;
  wire w_014_000, w_014_006, w_014_008, w_014_010, w_014_013, w_014_017, w_014_020, w_014_021, w_014_024, w_014_025, w_014_026, w_014_030, w_014_031, w_014_032, w_014_033, w_014_034, w_014_035, w_014_036, w_014_039, w_014_040, w_014_042, w_014_043, w_014_046, w_014_051, w_014_052, w_014_053, w_014_054, w_014_055, w_014_056, w_014_057, w_014_058, w_014_060, w_014_061, w_014_063, w_014_064, w_014_069, w_014_070, w_014_071, w_014_072, w_014_073, w_014_076, w_014_078, w_014_080, w_014_085, w_014_086, w_014_087, w_014_088, w_014_091, w_014_092, w_014_093, w_014_095, w_014_097, w_014_098, w_014_099, w_014_101, w_014_104, w_014_109, w_014_111, w_014_115, w_014_116, w_014_119, w_014_123, w_014_124, w_014_125, w_014_127, w_014_128, w_014_130, w_014_131, w_014_135, w_014_136, w_014_137, w_014_139, w_014_140, w_014_141, w_014_142, w_014_143, w_014_145, w_014_147, w_014_150, w_014_152, w_014_155, w_014_157, w_014_158, w_014_159, w_014_160, w_014_161, w_014_162, w_014_163, w_014_164, w_014_165, w_014_167, w_014_168, w_014_169, w_014_179, w_014_180, w_014_181, w_014_183, w_014_184, w_014_186, w_014_188, w_014_190, w_014_191, w_014_192, w_014_198, w_014_201, w_014_210, w_014_213, w_014_217, w_014_218, w_014_219, w_014_220, w_014_221, w_014_222, w_014_223, w_014_225, w_014_226, w_014_228, w_014_230, w_014_235, w_014_236, w_014_237, w_014_240, w_014_241, w_014_243, w_014_245, w_014_247, w_014_248, w_014_250, w_014_251, w_014_252, w_014_253, w_014_254, w_014_255, w_014_256, w_014_259, w_014_260, w_014_263, w_014_264, w_014_267, w_014_268, w_014_269, w_014_270, w_014_271, w_014_275, w_014_276, w_014_277, w_014_279, w_014_281, w_014_282, w_014_283, w_014_285, w_014_286, w_014_287, w_014_289, w_014_291, w_014_292, w_014_293, w_014_298, w_014_300, w_014_303, w_014_305, w_014_306, w_014_307, w_014_308, w_014_310, w_014_311, w_014_314, w_014_315, w_014_320, w_014_322, w_014_323, w_014_324, w_014_325, w_014_329, w_014_330, w_014_331, w_014_333, w_014_337, w_014_340, w_014_341, w_014_344, w_014_345, w_014_346, w_014_348, w_014_349, w_014_351, w_014_353, w_014_354, w_014_356, w_014_357, w_014_359, w_014_360, w_014_362, w_014_363, w_014_365, w_014_367, w_014_375, w_014_380, w_014_383, w_014_389, w_014_392, w_014_399, w_014_401, w_014_403, w_014_405, w_014_409, w_014_411, w_014_415, w_014_417, w_014_420, w_014_424, w_014_426, w_014_434, w_014_435, w_014_437, w_014_442, w_014_443, w_014_444, w_014_446, w_014_449, w_014_451, w_014_453, w_014_457, w_014_464, w_014_465, w_014_469, w_014_470, w_014_472, w_014_474, w_014_479, w_014_482, w_014_485, w_014_487, w_014_500, w_014_503, w_014_504, w_014_507, w_014_509, w_014_515, w_014_516, w_014_518, w_014_520, w_014_524, w_014_527, w_014_529, w_014_533, w_014_534, w_014_538, w_014_540, w_014_542, w_014_543, w_014_545, w_014_546, w_014_549, w_014_554, w_014_557, w_014_559, w_014_560, w_014_564, w_014_566, w_014_568, w_014_571, w_014_573, w_014_574, w_014_576, w_014_577, w_014_582, w_014_584, w_014_586, w_014_594, w_014_595, w_014_598, w_014_602, w_014_603, w_014_608, w_014_609, w_014_613, w_014_626, w_014_629, w_014_632, w_014_634, w_014_635, w_014_636, w_014_637;
  wire w_015_000, w_015_001, w_015_002, w_015_003, w_015_004, w_015_008, w_015_010, w_015_011, w_015_012, w_015_013, w_015_015, w_015_018, w_015_019, w_015_021, w_015_024, w_015_025, w_015_026, w_015_027, w_015_029, w_015_031, w_015_032, w_015_035, w_015_036, w_015_037, w_015_041, w_015_042, w_015_043, w_015_044, w_015_045, w_015_047, w_015_048, w_015_049, w_015_051, w_015_052, w_015_053, w_015_057, w_015_058, w_015_059, w_015_061, w_015_062, w_015_064, w_015_067, w_015_071, w_015_072, w_015_078, w_015_079, w_015_080, w_015_081, w_015_083, w_015_084, w_015_088, w_015_089, w_015_090, w_015_092, w_015_093, w_015_094, w_015_095, w_015_096, w_015_098, w_015_099, w_015_101, w_015_103, w_015_106, w_015_108, w_015_112, w_015_114, w_015_117, w_015_118, w_015_122, w_015_124, w_015_126, w_015_127, w_015_128, w_015_129, w_015_130, w_015_131, w_015_134, w_015_135, w_015_136, w_015_138, w_015_139, w_015_140, w_015_141, w_015_142, w_015_143, w_015_146, w_015_150, w_015_151, w_015_154, w_015_155, w_015_156, w_015_157, w_015_158, w_015_159, w_015_160, w_015_164, w_015_165, w_015_166, w_015_168, w_015_170, w_015_171, w_015_172, w_015_173, w_015_175, w_015_178, w_015_180, w_015_187, w_015_190, w_015_191, w_015_193, w_015_196, w_015_197, w_015_199, w_015_201, w_015_205, w_015_206, w_015_207, w_015_209, w_015_210, w_015_211, w_015_214, w_015_216, w_015_221, w_015_226, w_015_227, w_015_233, w_015_235, w_015_238, w_015_254, w_015_255, w_015_258, w_015_264, w_015_265, w_015_275, w_015_277, w_015_278, w_015_280, w_015_282, w_015_284, w_015_304, w_015_314, w_015_315, w_015_316, w_015_319, w_015_322, w_015_323, w_015_324, w_015_328, w_015_330, w_015_333, w_015_339, w_015_341, w_015_345, w_015_346, w_015_348, w_015_349, w_015_350, w_015_359, w_015_363, w_015_365, w_015_367, w_015_368, w_015_369, w_015_373, w_015_394, w_015_395, w_015_397, w_015_404, w_015_406, w_015_412, w_015_418, w_015_424, w_015_426, w_015_427, w_015_429, w_015_434, w_015_438, w_015_440, w_015_442, w_015_443, w_015_444, w_015_445, w_015_447, w_015_450, w_015_453, w_015_457, w_015_458, w_015_459, w_015_462, w_015_465, w_015_470, w_015_474, w_015_476, w_015_479, w_015_482, w_015_490, w_015_492, w_015_493, w_015_494, w_015_496, w_015_499, w_015_504, w_015_510, w_015_512, w_015_517, w_015_519, w_015_521, w_015_522, w_015_525, w_015_529, w_015_532, w_015_535, w_015_538, w_015_541, w_015_547, w_015_554, w_015_559, w_015_583, w_015_585, w_015_592, w_015_594, w_015_595, w_015_597, w_015_600, w_015_603, w_015_604, w_015_605, w_015_608, w_015_611, w_015_618, w_015_619, w_015_621, w_015_624, w_015_625, w_015_629, w_015_631, w_015_635, w_015_636, w_015_643, w_015_644, w_015_648, w_015_652, w_015_654, w_015_655, w_015_657, w_015_659, w_015_661, w_015_669, w_015_676, w_015_689, w_015_691, w_015_692, w_015_693, w_015_695, w_015_696, w_015_699, w_015_703, w_015_704, w_015_706, w_015_707, w_015_713, w_015_714, w_015_716, w_015_718, w_015_722, w_015_730, w_015_733, w_015_734, w_015_737, w_015_738, w_015_742, w_015_743, w_015_744, w_015_755, w_015_758, w_015_759, w_015_760, w_015_761, w_015_763, w_015_766, w_015_773, w_015_774, w_015_776, w_015_778, w_015_779, w_015_780, w_015_782, w_015_793;
  wire w_016_001, w_016_002, w_016_003, w_016_004, w_016_006, w_016_007, w_016_010, w_016_012, w_016_013, w_016_016, w_016_021, w_016_022, w_016_024, w_016_025, w_016_026, w_016_027, w_016_028, w_016_029, w_016_034, w_016_035, w_016_036, w_016_037, w_016_038, w_016_039, w_016_040, w_016_042, w_016_043, w_016_047, w_016_048, w_016_049, w_016_050, w_016_052, w_016_053, w_016_054, w_016_057, w_016_059, w_016_060, w_016_062, w_016_063, w_016_064, w_016_065, w_016_067, w_016_070, w_016_072, w_016_074, w_016_075, w_016_076, w_016_077, w_016_079, w_016_081, w_016_083, w_016_084, w_016_085, w_016_089, w_016_090, w_016_093, w_016_096, w_016_099, w_016_100, w_016_101, w_016_102, w_016_104, w_016_105, w_016_106, w_016_108, w_016_110, w_016_111, w_016_112, w_016_113, w_016_114, w_016_116, w_016_122, w_016_124, w_016_125, w_016_127, w_016_128, w_016_129, w_016_135, w_016_136, w_016_137, w_016_138, w_016_141, w_016_142, w_016_143, w_016_144, w_016_146, w_016_148, w_016_155, w_016_156, w_016_161, w_016_162, w_016_170, w_016_171, w_016_172, w_016_173, w_016_174, w_016_175, w_016_178, w_016_179, w_016_181, w_016_182, w_016_184, w_016_185, w_016_186, w_016_188, w_016_190, w_016_191, w_016_194, w_016_195, w_016_197, w_016_198, w_016_204, w_016_206, w_016_207, w_016_208, w_016_209, w_016_210, w_016_211, w_016_213, w_016_214, w_016_215, w_016_217, w_016_218, w_016_219, w_016_220, w_016_221, w_016_224, w_016_225, w_016_226, w_016_228, w_016_232, w_016_235, w_016_239, w_016_240, w_016_243, w_016_247, w_016_251, w_016_252, w_016_253, w_016_255, w_016_257, w_016_259, w_016_260, w_016_270, w_016_271, w_016_272, w_016_273, w_016_274, w_016_275, w_016_276, w_016_278, w_016_281, w_016_282, w_016_285, w_016_289, w_016_290, w_016_295, w_016_297, w_016_298, w_016_299, w_016_300, w_016_301, w_016_302, w_016_303, w_016_305, w_016_306, w_016_307, w_016_313, w_016_315, w_016_316, w_016_317, w_016_318, w_016_319, w_016_320, w_016_322, w_016_323, w_016_326, w_016_327, w_016_328, w_016_329, w_016_330, w_016_333, w_016_337, w_016_338, w_016_345, w_016_347, w_016_348, w_016_349, w_016_351, w_016_353, w_016_354, w_016_356, w_016_358, w_016_359, w_016_362, w_016_363, w_016_364, w_016_367, w_016_368, w_016_370, w_016_371, w_016_372, w_016_374, w_016_376, w_016_378, w_016_380, w_016_381, w_016_387, w_016_390, w_016_393, w_016_394, w_016_397, w_016_398, w_016_400, w_016_404, w_016_405, w_016_406, w_016_407, w_016_411, w_016_416, w_016_418, w_016_420, w_016_422, w_016_423, w_016_424, w_016_425, w_016_428, w_016_429, w_016_435, w_016_436, w_016_437, w_016_438, w_016_439, w_016_440, w_016_442, w_016_445, w_016_448, w_016_450, w_016_452, w_016_453, w_016_455, w_016_459, w_016_461, w_016_465, w_016_466, w_016_467, w_016_471, w_016_472, w_016_473, w_016_474, w_016_475, w_016_476, w_016_477, w_016_481, w_016_484, w_016_485, w_016_487, w_016_492, w_016_494, w_016_495, w_016_496, w_016_500, w_016_501;
  wire w_017_000, w_017_001, w_017_002, w_017_003, w_017_004, w_017_005, w_017_006, w_017_007, w_017_008, w_017_009, w_017_010, w_017_011, w_017_012, w_017_013, w_017_014, w_017_015, w_017_016, w_017_017, w_017_018, w_017_019, w_017_020, w_017_021, w_017_022, w_017_023, w_017_024, w_017_025, w_017_026, w_017_027;
  wire w_018_000, w_018_002, w_018_003, w_018_006, w_018_008, w_018_010, w_018_013, w_018_014, w_018_015, w_018_016, w_018_017, w_018_019, w_018_020, w_018_021, w_018_023, w_018_024, w_018_025, w_018_026, w_018_027, w_018_030, w_018_031, w_018_032, w_018_033, w_018_034, w_018_035, w_018_036, w_018_038, w_018_039, w_018_040, w_018_041, w_018_043, w_018_046, w_018_047, w_018_048, w_018_049, w_018_051, w_018_052, w_018_053, w_018_054, w_018_056, w_018_057, w_018_058, w_018_059, w_018_060, w_018_062, w_018_064, w_018_066, w_018_067, w_018_068, w_018_069, w_018_070, w_018_072, w_018_073, w_018_074, w_018_075, w_018_076, w_018_077, w_018_079, w_018_081, w_018_082, w_018_084, w_018_086, w_018_088, w_018_089, w_018_090, w_018_091, w_018_092, w_018_093, w_018_096, w_018_097, w_018_098, w_018_101, w_018_102, w_018_103, w_018_104, w_018_106, w_018_107, w_018_108, w_018_109, w_018_110, w_018_111, w_018_112, w_018_113, w_018_114, w_018_115, w_018_116, w_018_117, w_018_118, w_018_119, w_018_120, w_018_121, w_018_122, w_018_123, w_018_124, w_018_125, w_018_126, w_018_129, w_018_130, w_018_131, w_018_132, w_018_133, w_018_134, w_018_135, w_018_136, w_018_139, w_018_141, w_018_143, w_018_144, w_018_145, w_018_146, w_018_150, w_018_151, w_018_153, w_018_155, w_018_156, w_018_157, w_018_158, w_018_159, w_018_163, w_018_164, w_018_165, w_018_166, w_018_167, w_018_168, w_018_170, w_018_171, w_018_172, w_018_174, w_018_175, w_018_176, w_018_177, w_018_180, w_018_181, w_018_182, w_018_183, w_018_184, w_018_186, w_018_188, w_018_190, w_018_191, w_018_192, w_018_193, w_018_194, w_018_196, w_018_197, w_018_198;
  wire w_019_002, w_019_004, w_019_005, w_019_008, w_019_010, w_019_011, w_019_012, w_019_014, w_019_015, w_019_019, w_019_020, w_019_021, w_019_024, w_019_025, w_019_026, w_019_027, w_019_032, w_019_037, w_019_039, w_019_040, w_019_042, w_019_043, w_019_044, w_019_046, w_019_048, w_019_049, w_019_050, w_019_051, w_019_055, w_019_056, w_019_057, w_019_060, w_019_064, w_019_065, w_019_067, w_019_068, w_019_069, w_019_070, w_019_072, w_019_073, w_019_074, w_019_077, w_019_078, w_019_082, w_019_084, w_019_085, w_019_088, w_019_089, w_019_092, w_019_093, w_019_094, w_019_096, w_019_097, w_019_099, w_019_100, w_019_101, w_019_102, w_019_103, w_019_111, w_019_116, w_019_118, w_019_121, w_019_124, w_019_125, w_019_126, w_019_128, w_019_129, w_019_130, w_019_133, w_019_135, w_019_138, w_019_144, w_019_145, w_019_146, w_019_147, w_019_148, w_019_149, w_019_152, w_019_153, w_019_154, w_019_155, w_019_157, w_019_160, w_019_163, w_019_165, w_019_168, w_019_169, w_019_170, w_019_171, w_019_173, w_019_174, w_019_179, w_019_182, w_019_184, w_019_185, w_019_186, w_019_187, w_019_191, w_019_192, w_019_197, w_019_200, w_019_205, w_019_207, w_019_209, w_019_213, w_019_214, w_019_215, w_019_219, w_019_228, w_019_229, w_019_230, w_019_233, w_019_234, w_019_235, w_019_241, w_019_242, w_019_243, w_019_245, w_019_246, w_019_248, w_019_249, w_019_255, w_019_258, w_019_259, w_019_260, w_019_261, w_019_265, w_019_269, w_019_274, w_019_275, w_019_277, w_019_279, w_019_286, w_019_288, w_019_291, w_019_294, w_019_295, w_019_296, w_019_297, w_019_299, w_019_300, w_019_303, w_019_305, w_019_306, w_019_307, w_019_308, w_019_310, w_019_314, w_019_317, w_019_318, w_019_319, w_019_320, w_019_321, w_019_322, w_019_327, w_019_329, w_019_332, w_019_335, w_019_339, w_019_340, w_019_342, w_019_344, w_019_345, w_019_347, w_019_352, w_019_353, w_019_357, w_019_359, w_019_360, w_019_362, w_019_363, w_019_364, w_019_371, w_019_374, w_019_377, w_019_378, w_019_384, w_019_386, w_019_389, w_019_396, w_019_402, w_019_403, w_019_404, w_019_406, w_019_407, w_019_413, w_019_416, w_019_417, w_019_421;
  wire w_020_000, w_020_001, w_020_002, w_020_003, w_020_004, w_020_005, w_020_006, w_020_007, w_020_008, w_020_009, w_020_010, w_020_011, w_020_012, w_020_013, w_020_014, w_020_015, w_020_016, w_020_017, w_020_019, w_020_020, w_020_021, w_020_022, w_020_023, w_020_024, w_020_025, w_020_026, w_020_027, w_020_028, w_020_029, w_020_030, w_020_032, w_020_033, w_020_034, w_020_035, w_020_036, w_020_037, w_020_038, w_020_039, w_020_040, w_020_041, w_020_042, w_020_043, w_020_044, w_020_045, w_020_046, w_020_047, w_020_048, w_020_049, w_020_050, w_020_052, w_020_053, w_020_054, w_020_057, w_020_058, w_020_060, w_020_061, w_020_062, w_020_063, w_020_064, w_020_066, w_020_067, w_020_068, w_020_069, w_020_070, w_020_071, w_020_072, w_020_073, w_020_074, w_020_075, w_020_077, w_020_078, w_020_080, w_020_081, w_020_082, w_020_083, w_020_084, w_020_085, w_020_086, w_020_087, w_020_088, w_020_089, w_020_090, w_020_091, w_020_092, w_020_093, w_020_095, w_020_096, w_020_098, w_020_099, w_020_100, w_020_102, w_020_103, w_020_104, w_020_105, w_020_106, w_020_107, w_020_108, w_020_111, w_020_112, w_020_114, w_020_115, w_020_116, w_020_117, w_020_118, w_020_119, w_020_120, w_020_121, w_020_122, w_020_123, w_020_124, w_020_126, w_020_127, w_020_128, w_020_129, w_020_130, w_020_131, w_020_132, w_020_133, w_020_134, w_020_135, w_020_136, w_020_137;
  wire w_021_000, w_021_001, w_021_003, w_021_006, w_021_007, w_021_008, w_021_009, w_021_010, w_021_012, w_021_013, w_021_014, w_021_016, w_021_018, w_021_019, w_021_020, w_021_024, w_021_025, w_021_026, w_021_027, w_021_028, w_021_029, w_021_030, w_021_033, w_021_035, w_021_036, w_021_037, w_021_039, w_021_040, w_021_041, w_021_042, w_021_044, w_021_045, w_021_046, w_021_047, w_021_048, w_021_049, w_021_050, w_021_051, w_021_052, w_021_053, w_021_055, w_021_058, w_021_059, w_021_060, w_021_061, w_021_063, w_021_064, w_021_065, w_021_066, w_021_070, w_021_071, w_021_075, w_021_076, w_021_079, w_021_082, w_021_083, w_021_084, w_021_086, w_021_088, w_021_089, w_021_091, w_021_093, w_021_095, w_021_099, w_021_101, w_021_105, w_021_106, w_021_107, w_021_108, w_021_111, w_021_119, w_021_120, w_021_122, w_021_123, w_021_126, w_021_127, w_021_128, w_021_129, w_021_130, w_021_131, w_021_133, w_021_136, w_021_137, w_021_138, w_021_139, w_021_141, w_021_142, w_021_143, w_021_145, w_021_149, w_021_151, w_021_152, w_021_154, w_021_155, w_021_156, w_021_157, w_021_158, w_021_159, w_021_161, w_021_162, w_021_163, w_021_164, w_021_166, w_021_169, w_021_170, w_021_171, w_021_172, w_021_178, w_021_179, w_021_181, w_021_183, w_021_184, w_021_185, w_021_186, w_021_187, w_021_190, w_021_191, w_021_192, w_021_194, w_021_195, w_021_198, w_021_199, w_021_201, w_021_204, w_021_209, w_021_210, w_021_211, w_021_215, w_021_218, w_021_219, w_021_220, w_021_221, w_021_222, w_021_224, w_021_228, w_021_229, w_021_230, w_021_234, w_021_236, w_021_237, w_021_239, w_021_240, w_021_243, w_021_244, w_021_245, w_021_247, w_021_248, w_021_252, w_021_256, w_021_257, w_021_259, w_021_261, w_021_264, w_021_266, w_021_270, w_021_272, w_021_273, w_021_275, w_021_277, w_021_281, w_021_283, w_021_284, w_021_289, w_021_290, w_021_294, w_021_298, w_021_303, w_021_305, w_021_306, w_021_307, w_021_310, w_021_313, w_021_314, w_021_317, w_021_319, w_021_320, w_021_322, w_021_324, w_021_326, w_021_328, w_021_329, w_021_330, w_021_335, w_021_337, w_021_340, w_021_341, w_021_342, w_021_343, w_021_348, w_021_352, w_021_353, w_021_360;
  wire w_022_002, w_022_003, w_022_006, w_022_008, w_022_010, w_022_020, w_022_021, w_022_025, w_022_026, w_022_031, w_022_032, w_022_033, w_022_034, w_022_039, w_022_043, w_022_046, w_022_049, w_022_052, w_022_054, w_022_055, w_022_057, w_022_061, w_022_065, w_022_066, w_022_067, w_022_068, w_022_072, w_022_073, w_022_076, w_022_081, w_022_084, w_022_087, w_022_088, w_022_090, w_022_097, w_022_099, w_022_100, w_022_101, w_022_103, w_022_105, w_022_109, w_022_110, w_022_113, w_022_117, w_022_118, w_022_119, w_022_124, w_022_126, w_022_128, w_022_129, w_022_139, w_022_143, w_022_144, w_022_146, w_022_149, w_022_151, w_022_152, w_022_155, w_022_159, w_022_160, w_022_161, w_022_162, w_022_163, w_022_165, w_022_168, w_022_169, w_022_174, w_022_175, w_022_177, w_022_181, w_022_183, w_022_185, w_022_187, w_022_193, w_022_197, w_022_198, w_022_202, w_022_205, w_022_206, w_022_209, w_022_210, w_022_213, w_022_222, w_022_225, w_022_226, w_022_229, w_022_234, w_022_236, w_022_239, w_022_242, w_022_243, w_022_244, w_022_246, w_022_256, w_022_258, w_022_259, w_022_260, w_022_262, w_022_267, w_022_268, w_022_269, w_022_270, w_022_271, w_022_274, w_022_275, w_022_276, w_022_277, w_022_278, w_022_280, w_022_281, w_022_282, w_022_286, w_022_290, w_022_291, w_022_293, w_022_294, w_022_297, w_022_301, w_022_304, w_022_305, w_022_307, w_022_310, w_022_311, w_022_314, w_022_315, w_022_316, w_022_318, w_022_319, w_022_320, w_022_321, w_022_322, w_022_323, w_022_325, w_022_326, w_022_328, w_022_335, w_022_336, w_022_337, w_022_339, w_022_341, w_022_343, w_022_344, w_022_345, w_022_349, w_022_352, w_022_353, w_022_358, w_022_360, w_022_361, w_022_364, w_022_370, w_022_372, w_022_375, w_022_376, w_022_383, w_022_385, w_022_388, w_022_391, w_022_392, w_022_395, w_022_398, w_022_400, w_022_401, w_022_402, w_022_405, w_022_406, w_022_412, w_022_414, w_022_415, w_022_416, w_022_418, w_022_421, w_022_426, w_022_427, w_022_428, w_022_429, w_022_430, w_022_431, w_022_432, w_022_433, w_022_436, w_022_439, w_022_446, w_022_453, w_022_455, w_022_457, w_022_464, w_022_469, w_022_472, w_022_479, w_022_482, w_022_486, w_022_489, w_022_495, w_022_498, w_022_503, w_022_506, w_022_508, w_022_511, w_022_512, w_022_516, w_022_517, w_022_519, w_022_524, w_022_527, w_022_537, w_022_540, w_022_543;
  wire w_023_002, w_023_012, w_023_013, w_023_015, w_023_020, w_023_024, w_023_037, w_023_038, w_023_040, w_023_041, w_023_047, w_023_049, w_023_051, w_023_053, w_023_054, w_023_058, w_023_059, w_023_064, w_023_065, w_023_068, w_023_071, w_023_073, w_023_078, w_023_079, w_023_086, w_023_088, w_023_089, w_023_092, w_023_093, w_023_099, w_023_100, w_023_104, w_023_106, w_023_108, w_023_109, w_023_110, w_023_111, w_023_112, w_023_118, w_023_120, w_023_127, w_023_132, w_023_134, w_023_136, w_023_137, w_023_138, w_023_139, w_023_140, w_023_143, w_023_148, w_023_153, w_023_154, w_023_157, w_023_158, w_023_161, w_023_166, w_023_170, w_023_172, w_023_174, w_023_175, w_023_177, w_023_178, w_023_181, w_023_184, w_023_186, w_023_188, w_023_190, w_023_193, w_023_196, w_023_197, w_023_200, w_023_206, w_023_211, w_023_212, w_023_215, w_023_216, w_023_226, w_023_228, w_023_230, w_023_231, w_023_232, w_023_234, w_023_239, w_023_240, w_023_241, w_023_242, w_023_248, w_023_249, w_023_250, w_023_251, w_023_252, w_023_253, w_023_255, w_023_267, w_023_269, w_023_271, w_023_274, w_023_277, w_023_278, w_023_291, w_023_293, w_023_295, w_023_297, w_023_302, w_023_305, w_023_306, w_023_307, w_023_309, w_023_311, w_023_316, w_023_321, w_023_325, w_023_326, w_023_333, w_023_334, w_023_348, w_023_351, w_023_352, w_023_358, w_023_359, w_023_369, w_023_383, w_023_387, w_023_400, w_023_403, w_023_405, w_023_413, w_023_416, w_023_423, w_023_427, w_023_429, w_023_432, w_023_435, w_023_444, w_023_445, w_023_448, w_023_451, w_023_455, w_023_457, w_023_459, w_023_462, w_023_468, w_023_470, w_023_472, w_023_477, w_023_489, w_023_493, w_023_499, w_023_500, w_023_502, w_023_503, w_023_507, w_023_513, w_023_518, w_023_520, w_023_522, w_023_528, w_023_529, w_023_530, w_023_531, w_023_547, w_023_548, w_023_551, w_023_553, w_023_558, w_023_559, w_023_569, w_023_572, w_023_576, w_023_578, w_023_584, w_023_588, w_023_594, w_023_601, w_023_603, w_023_604, w_023_611, w_023_614, w_023_621, w_023_622, w_023_624, w_023_628, w_023_633, w_023_656, w_023_659, w_023_660, w_023_664, w_023_666, w_023_668, w_023_670, w_023_679;
  wire w_024_000, w_024_008, w_024_012, w_024_014, w_024_019, w_024_020, w_024_024, w_024_029, w_024_034, w_024_037, w_024_040, w_024_041, w_024_042, w_024_050, w_024_051, w_024_052, w_024_053, w_024_056, w_024_057, w_024_068, w_024_069, w_024_070, w_024_072, w_024_076, w_024_079, w_024_080, w_024_082, w_024_083, w_024_084, w_024_089, w_024_090, w_024_093, w_024_094, w_024_096, w_024_103, w_024_104, w_024_105, w_024_108, w_024_112, w_024_122, w_024_128, w_024_129, w_024_130, w_024_131, w_024_133, w_024_136, w_024_138, w_024_141, w_024_142, w_024_145, w_024_146, w_024_158, w_024_159, w_024_161, w_024_162, w_024_164, w_024_166, w_024_170, w_024_171, w_024_174, w_024_176, w_024_180, w_024_182, w_024_183, w_024_189, w_024_191, w_024_192, w_024_194, w_024_196, w_024_200, w_024_207, w_024_209, w_024_217, w_024_218, w_024_220, w_024_225, w_024_228, w_024_229, w_024_231, w_024_236, w_024_238, w_024_244, w_024_247, w_024_249, w_024_251, w_024_255, w_024_257, w_024_259, w_024_263, w_024_264, w_024_265, w_024_266, w_024_267, w_024_268, w_024_270, w_024_276, w_024_283, w_024_284, w_024_285, w_024_287, w_024_289, w_024_291, w_024_292, w_024_293, w_024_297, w_024_298, w_024_302, w_024_307, w_024_309, w_024_316, w_024_319, w_024_321, w_024_322, w_024_323, w_024_326, w_024_331, w_024_333, w_024_334, w_024_335, w_024_336, w_024_339, w_024_341, w_024_342, w_024_343, w_024_344, w_024_345, w_024_347, w_024_351, w_024_353, w_024_357, w_024_361, w_024_364, w_024_366, w_024_367, w_024_377, w_024_380, w_024_381, w_024_382, w_024_388, w_024_391, w_024_393, w_024_394, w_024_397, w_024_398, w_024_399, w_024_400, w_024_401, w_024_402, w_024_404, w_024_407, w_024_416, w_024_426, w_024_429, w_024_435, w_024_437, w_024_446, w_024_452, w_024_455, w_024_473, w_024_476, w_024_486, w_024_491, w_024_495, w_024_496, w_024_497, w_024_501, w_024_507, w_024_511, w_024_515, w_024_522, w_024_523, w_024_529, w_024_537, w_024_539, w_024_540, w_024_546, w_024_549, w_024_555, w_024_556, w_024_557, w_024_560, w_024_570, w_024_574, w_024_577, w_024_588, w_024_590, w_024_592;
  wire w_025_003, w_025_005, w_025_008, w_025_009, w_025_011, w_025_012, w_025_014, w_025_015, w_025_018, w_025_020, w_025_022, w_025_025, w_025_026, w_025_032, w_025_033, w_025_036, w_025_039, w_025_041, w_025_042, w_025_047, w_025_050, w_025_056, w_025_057, w_025_060, w_025_061, w_025_066, w_025_067, w_025_068, w_025_071, w_025_075, w_025_077, w_025_079, w_025_083, w_025_087, w_025_090, w_025_093, w_025_094, w_025_100, w_025_103, w_025_105, w_025_107, w_025_108, w_025_115, w_025_125, w_025_126, w_025_131, w_025_132, w_025_136, w_025_144, w_025_145, w_025_146, w_025_147, w_025_153, w_025_154, w_025_155, w_025_156, w_025_157, w_025_158, w_025_159, w_025_160, w_025_163, w_025_169, w_025_171, w_025_177, w_025_180, w_025_181, w_025_183, w_025_187, w_025_188, w_025_189, w_025_195, w_025_199, w_025_202, w_025_203, w_025_206, w_025_208, w_025_215, w_025_221, w_025_223, w_025_225, w_025_226, w_025_228, w_025_232, w_025_233, w_025_238, w_025_239, w_025_246, w_025_247, w_025_250, w_025_251, w_025_262, w_025_269, w_025_272, w_025_274, w_025_275, w_025_280, w_025_281, w_025_282, w_025_286, w_025_290, w_025_292, w_025_294, w_025_295, w_025_297, w_025_306, w_025_307, w_025_308, w_025_314, w_025_317, w_025_339, w_025_342, w_025_346, w_025_347, w_025_348, w_025_358, w_025_362, w_025_373, w_025_378, w_025_382, w_025_396, w_025_405, w_025_406, w_025_412, w_025_419, w_025_428, w_025_429, w_025_437, w_025_454, w_025_465, w_025_468, w_025_473, w_025_477, w_025_478, w_025_480, w_025_488, w_025_497, w_025_498, w_025_506, w_025_510, w_025_514, w_025_516, w_025_519, w_025_530, w_025_531, w_025_532, w_025_535, w_025_539, w_025_542, w_025_552, w_025_553, w_025_554, w_025_555, w_025_556, w_025_557, w_025_571, w_025_572, w_025_576, w_025_585, w_025_591, w_025_595, w_025_606, w_025_613, w_025_614, w_025_625, w_025_626, w_025_630, w_025_635, w_025_640, w_025_648, w_025_654, w_025_656, w_025_657, w_025_658, w_025_660, w_025_663, w_025_665, w_025_668, w_025_678;
  wire w_026_001, w_026_003, w_026_007, w_026_008, w_026_009, w_026_011, w_026_012, w_026_014, w_026_017, w_026_023, w_026_024, w_026_025, w_026_026, w_026_028, w_026_029, w_026_030, w_026_031, w_026_032, w_026_034, w_026_035, w_026_037, w_026_038, w_026_039, w_026_040, w_026_045, w_026_046, w_026_047, w_026_048, w_026_049, w_026_051, w_026_054, w_026_055, w_026_056, w_026_058, w_026_061, w_026_062, w_026_063, w_026_064, w_026_065, w_026_068, w_026_073, w_026_075, w_026_078, w_026_079, w_026_080, w_026_088, w_026_089, w_026_091, w_026_092, w_026_094, w_026_095, w_026_096, w_026_097, w_026_098, w_026_100, w_026_103, w_026_106, w_026_108, w_026_110, w_026_116, w_026_124, w_026_125, w_026_131, w_026_139, w_026_142, w_026_149, w_026_155, w_026_156, w_026_158, w_026_161, w_026_170, w_026_172, w_026_174, w_026_175, w_026_176, w_026_180, w_026_181, w_026_183, w_026_189, w_026_194, w_026_195, w_026_200, w_026_206, w_026_209, w_026_210, w_026_215, w_026_216, w_026_217, w_026_218, w_026_219, w_026_224, w_026_226, w_026_228, w_026_231, w_026_232, w_026_235, w_026_236, w_026_239, w_026_243, w_026_246, w_026_247, w_026_249, w_026_252, w_026_253, w_026_257, w_026_264, w_026_265, w_026_266, w_026_269, w_026_272, w_026_273, w_026_274, w_026_275, w_026_277, w_026_279, w_026_280, w_026_282, w_026_283, w_026_294, w_026_295, w_026_296, w_026_297, w_026_298, w_026_301, w_026_303, w_026_305, w_026_307, w_026_308, w_026_309, w_026_310, w_026_311, w_026_317, w_026_321, w_026_323, w_026_325, w_026_326, w_026_328, w_026_331, w_026_332, w_026_333, w_026_338, w_026_340, w_026_341, w_026_349, w_026_351, w_026_353, w_026_355, w_026_356, w_026_358, w_026_361, w_026_364, w_026_365, w_026_368, w_026_370, w_026_374, w_026_375, w_026_376, w_026_377, w_026_379, w_026_381, w_026_382, w_026_383, w_026_387, w_026_388, w_026_390, w_026_392, w_026_393, w_026_395, w_026_396, w_026_399, w_026_400, w_026_401, w_026_407, w_026_408, w_026_410, w_026_419, w_026_421, w_026_424, w_026_430, w_026_431, w_026_435, w_026_436, w_026_438;
  wire w_027_006, w_027_007, w_027_011, w_027_014, w_027_016, w_027_027, w_027_035, w_027_040, w_027_041, w_027_042, w_027_050, w_027_054, w_027_055, w_027_063, w_027_067, w_027_069, w_027_075, w_027_077, w_027_080, w_027_083, w_027_085, w_027_087, w_027_091, w_027_095, w_027_101, w_027_108, w_027_111, w_027_114, w_027_115, w_027_118, w_027_124, w_027_127, w_027_128, w_027_130, w_027_134, w_027_141, w_027_143, w_027_144, w_027_145, w_027_154, w_027_162, w_027_164, w_027_165, w_027_168, w_027_171, w_027_172, w_027_173, w_027_177, w_027_189, w_027_195, w_027_198, w_027_207, w_027_208, w_027_222, w_027_225, w_027_227, w_027_234, w_027_236, w_027_250, w_027_257, w_027_259, w_027_267, w_027_272, w_027_280, w_027_285, w_027_294, w_027_299, w_027_300, w_027_307, w_027_311, w_027_320, w_027_324, w_027_336, w_027_339, w_027_343, w_027_344, w_027_348, w_027_353, w_027_373, w_027_383, w_027_400, w_027_401, w_027_412, w_027_413, w_027_414, w_027_419, w_027_426, w_027_429, w_027_431, w_027_433, w_027_434, w_027_437, w_027_440, w_027_445, w_027_459, w_027_460, w_027_466, w_027_470, w_027_478, w_027_486, w_027_497, w_027_522, w_027_525, w_027_526, w_027_535, w_027_537, w_027_543, w_027_546, w_027_548, w_027_564, w_027_565, w_027_568, w_027_573, w_027_576, w_027_584, w_027_600, w_027_602, w_027_606, w_027_614, w_027_619, w_027_622, w_027_624, w_027_625, w_027_628, w_027_629, w_027_635, w_027_647, w_027_656, w_027_658, w_027_659, w_027_663, w_027_668, w_027_671, w_027_672, w_027_676, w_027_678, w_027_681, w_027_683, w_027_690, w_027_696, w_027_699, w_027_707, w_027_712, w_027_717, w_027_725, w_027_736, w_027_742, w_027_757, w_027_762, w_027_768, w_027_776, w_027_779, w_027_791, w_027_794, w_027_796, w_027_797, w_027_811, w_027_813, w_027_816, w_027_819, w_027_826;
  wire w_028_004, w_028_012, w_028_013, w_028_015, w_028_017, w_028_020, w_028_024, w_028_025, w_028_027, w_028_028, w_028_029, w_028_030, w_028_033, w_028_036, w_028_042, w_028_043, w_028_049, w_028_052, w_028_062, w_028_065, w_028_066, w_028_067, w_028_070, w_028_073, w_028_076, w_028_078, w_028_079, w_028_081, w_028_087, w_028_088, w_028_092, w_028_102, w_028_107, w_028_108, w_028_109, w_028_112, w_028_119, w_028_125, w_028_128, w_028_131, w_028_132, w_028_135, w_028_143, w_028_144, w_028_146, w_028_156, w_028_161, w_028_162, w_028_167, w_028_171, w_028_180, w_028_186, w_028_201, w_028_202, w_028_206, w_028_210, w_028_211, w_028_216, w_028_218, w_028_219, w_028_220, w_028_222, w_028_234, w_028_235, w_028_237, w_028_241, w_028_246, w_028_258, w_028_276, w_028_277, w_028_281, w_028_289, w_028_294, w_028_296, w_028_302, w_028_311, w_028_313, w_028_318, w_028_323, w_028_326, w_028_328, w_028_345, w_028_349, w_028_358, w_028_359, w_028_360, w_028_366, w_028_368, w_028_369, w_028_371, w_028_376, w_028_397, w_028_403, w_028_404, w_028_406, w_028_411, w_028_424, w_028_427, w_028_429, w_028_432, w_028_436, w_028_439, w_028_440, w_028_442, w_028_456, w_028_462, w_028_468, w_028_470, w_028_472, w_028_475, w_028_482, w_028_487, w_028_492, w_028_494, w_028_496, w_028_506, w_028_509, w_028_511, w_028_527, w_028_535, w_028_544, w_028_546, w_028_566, w_028_567, w_028_573, w_028_574, w_028_577, w_028_581, w_028_590, w_028_595, w_028_599, w_028_613, w_028_615, w_028_625, w_028_626, w_028_629, w_028_630, w_028_631, w_028_638, w_028_647, w_028_648, w_028_652, w_028_664, w_028_682, w_028_693, w_028_709, w_028_715, w_028_728, w_028_729, w_028_735, w_028_739, w_028_745, w_028_762, w_028_764, w_028_767, w_028_768, w_028_777, w_028_783, w_028_785, w_028_793, w_028_799, w_028_811, w_028_817, w_028_827, w_028_848, w_028_854, w_028_855, w_028_862, w_028_875, w_028_876, w_028_877, w_028_882, w_028_885, w_028_886, w_028_890, w_028_895, w_028_899, w_028_900;
  wire w_029_004, w_029_007, w_029_008, w_029_009, w_029_010, w_029_011, w_029_016, w_029_020, w_029_021, w_029_024, w_029_026, w_029_027, w_029_029, w_029_030, w_029_031, w_029_034, w_029_035, w_029_036, w_029_038, w_029_039, w_029_040, w_029_041, w_029_042, w_029_044, w_029_046, w_029_047, w_029_050, w_029_051, w_029_054, w_029_056, w_029_061, w_029_062, w_029_063, w_029_064, w_029_067, w_029_070, w_029_071, w_029_072, w_029_073, w_029_075, w_029_077, w_029_080, w_029_082, w_029_084, w_029_086, w_029_087, w_029_089, w_029_092, w_029_093, w_029_094, w_029_096, w_029_099, w_029_101, w_029_103, w_029_106, w_029_110, w_029_111, w_029_113, w_029_114, w_029_115, w_029_116, w_029_117, w_029_118, w_029_119, w_029_120, w_029_123, w_029_124, w_029_125, w_029_126, w_029_129, w_029_130, w_029_131, w_029_133, w_029_134, w_029_135, w_029_136, w_029_138, w_029_139, w_029_140, w_029_148, w_029_149, w_029_151, w_029_154, w_029_157, w_029_158, w_029_160, w_029_162, w_029_163, w_029_166, w_029_171, w_029_173, w_029_174, w_029_178, w_029_183, w_029_186, w_029_187, w_029_188, w_029_189, w_029_190, w_029_191, w_029_192, w_029_193, w_029_196, w_029_199, w_029_202, w_029_207, w_029_209, w_029_211, w_029_214, w_029_215, w_029_216, w_029_217, w_029_218;
  wire w_030_001, w_030_002, w_030_003, w_030_004, w_030_005, w_030_010, w_030_011, w_030_012, w_030_016, w_030_019, w_030_028, w_030_030, w_030_031, w_030_033, w_030_035, w_030_038, w_030_041, w_030_044, w_030_045, w_030_046, w_030_049, w_030_050, w_030_052, w_030_053, w_030_064, w_030_071, w_030_072, w_030_073, w_030_075, w_030_076, w_030_080, w_030_082, w_030_089, w_030_105, w_030_109, w_030_123, w_030_133, w_030_145, w_030_149, w_030_151, w_030_152, w_030_158, w_030_160, w_030_163, w_030_166, w_030_174, w_030_176, w_030_177, w_030_178, w_030_182, w_030_184, w_030_186, w_030_189, w_030_193, w_030_194, w_030_196, w_030_198, w_030_201, w_030_202, w_030_203, w_030_205, w_030_206, w_030_210, w_030_216, w_030_217, w_030_230, w_030_231, w_030_234, w_030_239, w_030_240, w_030_242, w_030_244, w_030_246, w_030_247, w_030_248, w_030_252, w_030_253, w_030_255, w_030_258, w_030_265, w_030_269, w_030_271, w_030_274, w_030_275, w_030_281, w_030_282, w_030_287, w_030_288, w_030_294, w_030_305, w_030_308, w_030_311, w_030_312, w_030_314, w_030_318, w_030_324, w_030_335, w_030_340, w_030_341, w_030_342, w_030_347, w_030_353, w_030_357, w_030_358, w_030_360, w_030_362, w_030_364, w_030_367, w_030_371, w_030_380, w_030_385, w_030_386, w_030_387, w_030_390, w_030_391, w_030_399, w_030_401, w_030_405, w_030_408, w_030_409, w_030_410, w_030_412, w_030_415, w_030_418, w_030_420, w_030_423, w_030_424, w_030_433, w_030_435, w_030_438, w_030_444, w_030_445, w_030_450, w_030_461, w_030_462, w_030_463, w_030_468, w_030_473, w_030_477, w_030_478, w_030_480, w_030_481, w_030_483, w_030_484, w_030_487, w_030_490, w_030_491, w_030_495;
  wire w_031_002, w_031_003, w_031_004, w_031_010, w_031_011, w_031_015, w_031_016, w_031_017, w_031_019, w_031_023, w_031_025, w_031_027, w_031_030, w_031_031, w_031_035, w_031_043, w_031_045, w_031_050, w_031_055, w_031_057, w_031_071, w_031_078, w_031_082, w_031_085, w_031_087, w_031_089, w_031_090, w_031_091, w_031_094, w_031_095, w_031_103, w_031_118, w_031_121, w_031_123, w_031_130, w_031_135, w_031_150, w_031_154, w_031_161, w_031_167, w_031_171, w_031_178, w_031_183, w_031_187, w_031_194, w_031_196, w_031_198, w_031_199, w_031_204, w_031_210, w_031_211, w_031_212, w_031_215, w_031_216, w_031_219, w_031_224, w_031_227, w_031_229, w_031_232, w_031_234, w_031_235, w_031_240, w_031_241, w_031_243, w_031_244, w_031_246, w_031_247, w_031_251, w_031_261, w_031_270, w_031_277, w_031_280, w_031_288, w_031_293, w_031_294, w_031_296, w_031_297, w_031_298, w_031_299, w_031_302, w_031_303, w_031_306, w_031_308, w_031_310, w_031_312, w_031_314, w_031_319, w_031_324, w_031_329, w_031_332, w_031_333, w_031_340, w_031_345, w_031_347, w_031_355, w_031_362, w_031_364, w_031_365, w_031_367, w_031_368, w_031_373, w_031_374, w_031_382, w_031_391, w_031_399, w_031_406, w_031_409, w_031_410, w_031_413, w_031_420, w_031_421, w_031_438, w_031_442, w_031_443, w_031_446, w_031_454;
  wire w_032_003, w_032_007, w_032_010, w_032_012, w_032_014, w_032_020, w_032_023, w_032_031, w_032_033, w_032_047, w_032_051, w_032_057, w_032_060, w_032_064, w_032_074, w_032_092, w_032_095, w_032_096, w_032_098, w_032_100, w_032_107, w_032_113, w_032_116, w_032_119, w_032_121, w_032_124, w_032_126, w_032_127, w_032_130, w_032_144, w_032_146, w_032_148, w_032_151, w_032_161, w_032_162, w_032_169, w_032_170, w_032_175, w_032_178, w_032_179, w_032_180, w_032_187, w_032_188, w_032_204, w_032_210, w_032_212, w_032_225, w_032_227, w_032_232, w_032_233, w_032_234, w_032_237, w_032_238, w_032_259, w_032_267, w_032_268, w_032_289, w_032_292, w_032_297, w_032_298, w_032_307, w_032_308, w_032_315, w_032_322, w_032_332, w_032_336, w_032_347, w_032_354, w_032_362, w_032_365, w_032_370, w_032_372, w_032_376, w_032_378, w_032_380, w_032_383, w_032_397, w_032_406, w_032_416, w_032_421, w_032_424, w_032_449, w_032_454, w_032_455, w_032_466, w_032_477, w_032_498, w_032_499, w_032_523, w_032_546, w_032_548, w_032_554, w_032_556, w_032_570, w_032_585, w_032_588, w_032_591, w_032_593, w_032_594, w_032_596, w_032_602, w_032_603, w_032_636, w_032_649, w_032_654, w_032_655, w_032_658, w_032_668, w_032_692, w_032_705, w_032_707, w_032_715, w_032_716, w_032_732, w_032_738, w_032_753, w_032_759, w_032_762, w_032_765, w_032_777, w_032_778, w_032_790, w_032_803, w_032_804, w_032_807, w_032_810;
  wire w_033_004, w_033_006, w_033_007, w_033_011, w_033_015, w_033_016, w_033_030, w_033_031, w_033_037, w_033_038, w_033_040, w_033_041, w_033_042, w_033_043, w_033_045, w_033_049, w_033_050, w_033_052, w_033_053, w_033_067, w_033_071, w_033_074, w_033_084, w_033_099, w_033_116, w_033_124, w_033_135, w_033_145, w_033_174, w_033_182, w_033_190, w_033_192, w_033_193, w_033_195, w_033_196, w_033_202, w_033_208, w_033_210, w_033_218, w_033_221, w_033_232, w_033_247, w_033_254, w_033_257, w_033_267, w_033_268, w_033_283, w_033_294, w_033_296, w_033_301, w_033_307, w_033_311, w_033_314, w_033_315, w_033_319, w_033_325, w_033_326, w_033_339, w_033_345, w_033_352, w_033_354, w_033_358, w_033_361, w_033_372, w_033_384, w_033_386, w_033_391, w_033_397, w_033_402, w_033_405, w_033_406, w_033_407, w_033_414, w_033_416, w_033_420, w_033_428, w_033_435, w_033_437, w_033_454, w_033_467, w_033_471, w_033_493, w_033_497, w_033_499, w_033_511, w_033_525, w_033_535, w_033_546, w_033_547, w_033_548, w_033_549, w_033_568, w_033_569, w_033_571, w_033_594, w_033_597, w_033_598, w_033_601, w_033_610, w_033_613, w_033_629, w_033_630, w_033_645, w_033_675, w_033_679, w_033_691, w_033_692, w_033_699, w_033_700, w_033_709, w_033_718, w_033_721, w_033_723, w_033_726, w_033_736, w_033_739, w_033_751, w_033_763, w_033_771, w_033_773, w_033_778, w_033_788, w_033_805, w_033_815, w_033_834, w_033_849, w_033_856, w_033_862, w_033_878, w_033_897, w_033_902, w_033_905, w_033_909;
  wire w_034_001, w_034_005, w_034_012, w_034_013, w_034_018, w_034_022, w_034_023, w_034_028, w_034_031, w_034_032, w_034_033, w_034_034, w_034_041, w_034_042, w_034_043, w_034_044, w_034_045, w_034_054, w_034_060, w_034_063, w_034_068, w_034_076, w_034_087, w_034_088, w_034_089, w_034_091, w_034_092, w_034_093, w_034_096, w_034_099, w_034_100, w_034_101, w_034_103, w_034_104, w_034_113, w_034_115, w_034_116, w_034_122, w_034_123, w_034_124, w_034_127, w_034_130, w_034_136, w_034_137, w_034_138, w_034_145, w_034_149, w_034_154, w_034_160, w_034_164, w_034_177, w_034_184, w_034_194, w_034_197, w_034_206, w_034_210, w_034_211, w_034_214, w_034_217, w_034_220, w_034_227, w_034_234, w_034_235, w_034_241, w_034_242, w_034_250, w_034_260, w_034_266, w_034_270, w_034_296, w_034_317, w_034_334, w_034_344, w_034_351, w_034_414, w_034_422, w_034_429, w_034_431, w_034_433, w_034_435, w_034_446, w_034_451, w_034_458, w_034_478, w_034_483, w_034_495, w_034_501, w_034_527, w_034_534, w_034_539, w_034_554, w_034_555, w_034_567, w_034_573, w_034_579, w_034_583, w_034_588, w_034_596, w_034_618, w_034_640, w_034_666, w_034_672, w_034_681, w_034_684, w_034_691, w_034_693, w_034_721, w_034_725, w_034_729, w_034_775, w_034_785, w_034_792, w_034_798, w_034_801, w_034_805, w_034_806;
  wire w_035_003, w_035_006, w_035_009, w_035_015, w_035_024, w_035_025, w_035_032, w_035_041, w_035_051, w_035_054, w_035_072, w_035_074, w_035_078, w_035_081, w_035_083, w_035_089, w_035_092, w_035_102, w_035_114, w_035_120, w_035_121, w_035_127, w_035_129, w_035_132, w_035_134, w_035_135, w_035_142, w_035_145, w_035_150, w_035_152, w_035_156, w_035_160, w_035_163, w_035_167, w_035_169, w_035_170, w_035_179, w_035_184, w_035_191, w_035_192, w_035_195, w_035_199, w_035_212, w_035_214, w_035_220, w_035_225, w_035_230, w_035_245, w_035_258, w_035_261, w_035_265, w_035_268, w_035_274, w_035_277, w_035_286, w_035_292, w_035_297, w_035_304, w_035_307, w_035_313, w_035_323, w_035_324, w_035_326, w_035_335, w_035_346, w_035_351, w_035_370, w_035_374, w_035_382, w_035_397, w_035_400, w_035_415, w_035_429, w_035_460, w_035_467, w_035_473, w_035_479, w_035_480, w_035_487, w_035_492, w_035_518, w_035_524, w_035_527, w_035_532, w_035_535, w_035_539, w_035_540, w_035_554, w_035_563, w_035_574, w_035_578, w_035_588, w_035_592, w_035_598, w_035_607, w_035_612, w_035_616, w_035_622, w_035_629, w_035_631, w_035_633, w_035_651, w_035_652, w_035_653, w_035_654, w_035_655, w_035_656, w_035_657, w_035_658, w_035_659, w_035_660;
  wire w_036_005, w_036_008, w_036_009, w_036_013, w_036_016, w_036_018, w_036_019, w_036_021, w_036_023, w_036_031, w_036_036, w_036_040, w_036_042, w_036_043, w_036_046, w_036_052, w_036_056, w_036_061, w_036_066, w_036_068, w_036_069, w_036_070, w_036_071, w_036_073, w_036_080, w_036_082, w_036_084, w_036_085, w_036_089, w_036_090, w_036_092, w_036_093, w_036_095, w_036_097, w_036_102, w_036_103, w_036_105, w_036_111, w_036_112, w_036_113, w_036_115, w_036_122, w_036_123, w_036_125, w_036_131, w_036_132, w_036_134, w_036_138, w_036_143, w_036_145, w_036_146, w_036_147, w_036_149, w_036_151, w_036_153, w_036_154, w_036_156, w_036_158, w_036_166, w_036_171, w_036_175, w_036_177, w_036_185, w_036_193, w_036_197, w_036_199, w_036_201, w_036_205, w_036_209, w_036_217, w_036_222, w_036_228, w_036_233, w_036_234, w_036_237, w_036_238, w_036_239, w_036_247, w_036_249, w_036_260, w_036_262, w_036_266, w_036_271, w_036_273, w_036_276, w_036_277, w_036_278, w_036_282, w_036_283, w_036_285, w_036_286, w_036_287, w_036_288, w_036_289, w_036_290;
  wire w_037_000, w_037_001, w_037_004, w_037_005, w_037_006, w_037_008, w_037_009, w_037_011, w_037_012, w_037_013, w_037_014, w_037_016, w_037_017, w_037_019, w_037_020, w_037_022, w_037_024, w_037_025, w_037_026, w_037_027, w_037_032, w_037_036, w_037_039, w_037_040, w_037_041, w_037_043, w_037_047, w_037_049, w_037_051, w_037_052, w_037_055, w_037_061, w_037_063, w_037_064, w_037_066, w_037_067, w_037_070, w_037_073, w_037_074, w_037_076, w_037_077, w_037_079, w_037_081, w_037_085, w_037_090, w_037_091, w_037_095, w_037_096, w_037_097, w_037_098, w_037_099, w_037_103, w_037_105, w_037_106, w_037_107, w_037_109, w_037_111, w_037_112, w_037_113, w_037_114, w_037_115, w_037_116, w_037_119, w_037_122, w_037_124, w_037_127, w_037_128, w_037_130, w_037_131, w_037_133, w_037_140, w_037_141, w_037_142, w_037_145, w_037_147, w_037_148, w_037_149, w_037_152, w_037_154, w_037_162, w_037_163, w_037_164, w_037_165, w_037_171, w_037_176, w_037_180, w_037_183, w_037_187, w_037_189, w_037_190;
  wire w_038_009, w_038_012, w_038_015, w_038_028, w_038_031, w_038_035, w_038_037, w_038_038, w_038_041, w_038_046, w_038_047, w_038_049, w_038_050, w_038_057, w_038_094, w_038_101, w_038_114, w_038_117, w_038_118, w_038_119, w_038_122, w_038_123, w_038_135, w_038_148, w_038_149, w_038_156, w_038_157, w_038_168, w_038_172, w_038_173, w_038_177, w_038_180, w_038_186, w_038_188, w_038_190, w_038_194, w_038_202, w_038_206, w_038_224, w_038_227, w_038_235, w_038_238, w_038_277, w_038_303, w_038_305, w_038_324, w_038_335, w_038_345, w_038_388, w_038_413, w_038_432, w_038_447, w_038_448, w_038_459, w_038_469, w_038_489, w_038_521, w_038_526, w_038_543, w_038_548, w_038_559, w_038_560, w_038_562, w_038_565, w_038_573, w_038_591, w_038_612, w_038_621, w_038_625, w_038_637, w_038_640, w_038_644, w_038_648, w_038_665, w_038_689, w_038_694, w_038_696, w_038_701, w_038_709, w_038_713, w_038_735, w_038_747, w_038_748, w_038_762, w_038_764;
  wire w_039_002, w_039_003, w_039_005, w_039_007, w_039_008, w_039_010, w_039_013, w_039_017, w_039_023, w_039_031, w_039_033, w_039_036, w_039_037, w_039_040, w_039_047, w_039_049, w_039_051, w_039_056, w_039_057, w_039_062, w_039_066, w_039_067, w_039_074, w_039_089, w_039_096, w_039_103, w_039_116, w_039_119, w_039_122, w_039_125, w_039_128, w_039_129, w_039_136, w_039_144, w_039_145, w_039_146, w_039_149, w_039_153, w_039_162, w_039_164, w_039_170, w_039_175, w_039_180, w_039_183, w_039_184, w_039_187, w_039_188, w_039_189, w_039_190, w_039_197, w_039_201, w_039_204, w_039_228, w_039_232, w_039_234, w_039_235, w_039_243, w_039_250, w_039_253, w_039_259, w_039_265, w_039_268, w_039_277, w_039_284, w_039_288, w_039_289, w_039_299, w_039_303, w_039_305, w_039_309, w_039_310, w_039_312, w_039_332, w_039_333, w_039_336, w_039_340, w_039_349, w_039_362, w_039_371, w_039_375, w_039_377, w_039_381, w_039_382, w_039_385, w_039_392, w_039_395, w_039_400, w_039_405, w_039_413, w_039_417, w_039_427, w_039_431, w_039_443, w_039_444, w_039_450, w_039_456, w_039_459, w_039_460, w_039_461;
  wire w_040_003, w_040_008, w_040_016, w_040_017, w_040_025, w_040_026, w_040_027, w_040_029, w_040_033, w_040_037, w_040_043, w_040_048, w_040_057, w_040_058, w_040_060, w_040_066, w_040_068, w_040_071, w_040_075, w_040_083, w_040_084, w_040_089, w_040_095, w_040_098, w_040_102, w_040_103, w_040_104, w_040_105, w_040_110, w_040_111, w_040_112, w_040_113, w_040_115, w_040_116, w_040_117, w_040_122, w_040_126, w_040_127, w_040_128, w_040_131, w_040_132, w_040_140, w_040_141, w_040_142, w_040_148, w_040_149, w_040_151, w_040_152, w_040_155, w_040_156, w_040_158, w_040_159, w_040_167, w_040_168, w_040_169, w_040_170, w_040_173, w_040_175, w_040_176, w_040_178, w_040_182, w_040_186, w_040_194, w_040_201, w_040_204, w_040_207, w_040_210, w_040_215, w_040_217, w_040_219, w_040_224, w_040_230, w_040_235, w_040_237, w_040_243, w_040_245, w_040_248, w_040_250, w_040_252, w_040_254, w_040_257, w_040_259, w_040_264, w_040_272, w_040_274, w_040_294, w_040_298, w_040_302, w_040_305, w_040_306, w_040_308, w_040_314, w_040_316, w_040_320, w_040_321, w_040_322, w_040_323, w_040_325, w_040_327, w_040_331, w_040_338, w_040_340, w_040_347, w_040_355, w_040_357, w_040_361;
  wire w_041_000, w_041_001, w_041_002, w_041_003, w_041_005, w_041_007, w_041_008, w_041_009, w_041_010, w_041_011, w_041_012, w_041_014, w_041_015, w_041_016, w_041_017, w_041_018, w_041_019, w_041_020, w_041_022, w_041_023, w_041_026, w_041_027, w_041_028, w_041_031, w_041_032, w_041_033, w_041_035, w_041_036, w_041_037, w_041_039, w_041_043, w_041_044, w_041_045, w_041_047, w_041_048, w_041_049, w_041_050, w_041_052, w_041_054, w_041_055, w_041_057, w_041_058, w_041_060, w_041_061, w_041_062, w_041_068, w_041_070, w_041_071, w_041_073, w_041_075, w_041_076, w_041_077, w_041_078, w_041_079, w_041_082, w_041_083, w_041_084, w_041_085, w_041_086, w_041_089, w_041_091, w_041_094, w_041_096, w_041_097, w_041_098, w_041_099, w_041_100, w_041_101, w_041_102, w_041_104, w_041_106, w_041_107, w_041_111, w_041_112, w_041_113, w_041_114, w_041_115, w_041_116, w_041_117, w_041_118, w_041_119, w_041_120, w_041_121, w_041_122;
  wire w_042_001, w_042_002, w_042_003, w_042_004, w_042_005, w_042_006, w_042_011, w_042_012, w_042_013, w_042_014, w_042_016, w_042_017, w_042_018, w_042_021, w_042_024, w_042_026, w_042_028, w_042_031, w_042_033, w_042_041, w_042_042, w_042_043, w_042_045, w_042_046, w_042_050, w_042_052, w_042_055, w_042_056, w_042_057, w_042_059, w_042_064, w_042_065, w_042_066, w_042_067, w_042_068, w_042_069, w_042_070, w_042_074, w_042_077, w_042_078, w_042_081, w_042_083, w_042_084, w_042_094, w_042_097, w_042_098, w_042_099, w_042_103, w_042_108, w_042_110, w_042_114;
  wire w_043_000, w_043_001, w_043_002, w_043_003, w_043_004, w_043_005, w_043_006, w_043_007, w_043_009, w_043_010, w_043_011, w_043_013, w_043_014, w_043_015, w_043_016, w_043_017, w_043_018, w_043_019, w_043_020, w_043_021, w_043_022, w_043_023, w_043_024, w_043_025, w_043_027, w_043_028, w_043_029, w_043_031, w_043_032, w_043_035, w_043_036, w_043_038, w_043_039, w_043_040, w_043_041, w_043_042, w_043_043, w_043_044, w_043_045, w_043_046, w_043_047, w_043_048, w_043_049, w_043_051, w_043_052, w_043_053, w_043_054, w_043_055, w_043_057, w_043_058, w_043_059, w_043_060, w_043_061, w_043_062, w_043_063, w_043_064, w_043_065;
  wire w_044_007, w_044_012, w_044_014, w_044_015, w_044_017, w_044_024, w_044_031, w_044_033, w_044_036, w_044_037, w_044_038, w_044_039, w_044_040, w_044_043, w_044_047, w_044_048, w_044_049, w_044_051, w_044_055, w_044_058, w_044_061, w_044_063, w_044_067, w_044_070, w_044_075, w_044_083, w_044_093, w_044_105, w_044_107, w_044_110, w_044_114, w_044_118, w_044_120, w_044_128, w_044_133, w_044_139, w_044_140, w_044_142, w_044_145, w_044_155, w_044_156, w_044_159, w_044_162, w_044_166, w_044_172, w_044_174, w_044_175, w_044_181, w_044_183, w_044_184, w_044_188, w_044_193, w_044_194, w_044_198, w_044_199, w_044_203, w_044_216, w_044_219, w_044_220, w_044_223, w_044_227, w_044_231, w_044_232, w_044_234, w_044_261, w_044_263, w_044_273, w_044_274, w_044_276, w_044_278, w_044_292, w_044_296, w_044_304, w_044_310, w_044_312, w_044_314, w_044_315, w_044_323, w_044_338, w_044_341, w_044_343, w_044_347, w_044_348, w_044_356, w_044_360, w_044_365, w_044_371, w_044_378, w_044_384, w_044_386, w_044_391, w_044_392;
  wire w_045_001, w_045_004, w_045_005, w_045_006, w_045_013, w_045_016, w_045_018, w_045_021, w_045_029, w_045_043, w_045_053, w_045_067, w_045_074, w_045_076, w_045_079, w_045_092, w_045_093, w_045_102, w_045_105, w_045_106, w_045_108, w_045_110, w_045_111, w_045_123, w_045_127, w_045_128, w_045_141, w_045_142, w_045_145, w_045_149, w_045_151, w_045_153, w_045_160, w_045_165, w_045_170, w_045_175, w_045_179, w_045_192, w_045_193, w_045_203, w_045_206, w_045_214, w_045_223, w_045_226, w_045_227, w_045_229, w_045_243, w_045_252, w_045_253, w_045_255, w_045_258, w_045_271, w_045_277, w_045_281, w_045_294, w_045_296, w_045_315, w_045_323, w_045_324, w_045_328, w_045_339, w_045_340, w_045_341, w_045_348, w_045_353, w_045_382, w_045_411, w_045_415, w_045_421, w_045_440, w_045_443, w_045_467, w_045_474, w_045_500, w_045_503, w_045_505, w_045_506, w_045_511, w_045_531, w_045_534, w_045_548, w_045_549, w_045_560, w_045_563, w_045_564, w_045_567, w_045_593, w_045_629, w_045_633, w_045_662, w_045_667, w_045_692;
  wire w_046_000, w_046_006, w_046_012, w_046_029, w_046_035, w_046_048, w_046_052, w_046_059, w_046_062, w_046_067, w_046_070, w_046_076, w_046_091, w_046_097, w_046_098, w_046_115, w_046_120, w_046_122, w_046_141, w_046_143, w_046_148, w_046_156, w_046_157, w_046_158, w_046_171, w_046_176, w_046_178, w_046_179, w_046_181, w_046_182, w_046_184, w_046_185, w_046_194, w_046_195, w_046_212, w_046_294, w_046_300, w_046_305, w_046_310, w_046_324, w_046_327, w_046_328, w_046_333, w_046_342, w_046_367, w_046_386, w_046_393, w_046_414, w_046_420, w_046_421, w_046_422, w_046_461, w_046_467, w_046_479, w_046_488, w_046_497, w_046_501, w_046_504, w_046_510, w_046_525, w_046_539, w_046_540, w_046_545, w_046_546, w_046_559, w_046_572, w_046_614, w_046_627, w_046_642, w_046_660, w_046_664, w_046_669, w_046_673, w_046_674, w_046_689, w_046_697, w_046_733, w_046_734, w_046_767;
  wire w_047_001, w_047_006, w_047_033, w_047_056, w_047_062, w_047_066, w_047_067, w_047_082, w_047_095, w_047_096, w_047_098, w_047_105, w_047_107, w_047_118, w_047_124, w_047_146, w_047_157, w_047_158, w_047_164, w_047_171, w_047_176, w_047_178, w_047_183, w_047_187, w_047_188, w_047_190, w_047_203, w_047_208, w_047_212, w_047_226, w_047_229, w_047_230, w_047_232, w_047_238, w_047_244, w_047_245, w_047_247, w_047_257, w_047_262, w_047_272, w_047_278, w_047_279, w_047_281, w_047_288, w_047_289, w_047_295, w_047_327, w_047_332, w_047_339, w_047_348, w_047_357, w_047_364, w_047_379, w_047_385, w_047_386, w_047_396, w_047_401, w_047_404, w_047_427, w_047_436, w_047_443, w_047_448, w_047_450, w_047_460, w_047_464, w_047_470, w_047_472, w_047_474, w_047_475, w_047_481, w_047_485, w_047_492;
  wire w_048_018, w_048_023, w_048_029, w_048_034, w_048_050, w_048_068, w_048_070, w_048_078, w_048_089, w_048_090, w_048_095, w_048_097, w_048_101, w_048_111, w_048_114, w_048_116, w_048_118, w_048_121, w_048_133, w_048_136, w_048_139, w_048_158, w_048_161, w_048_188, w_048_189, w_048_198, w_048_201, w_048_203, w_048_205, w_048_218, w_048_227, w_048_276, w_048_285, w_048_296, w_048_308, w_048_313, w_048_320, w_048_335, w_048_348, w_048_368, w_048_380, w_048_384, w_048_385, w_048_410, w_048_412, w_048_418, w_048_427, w_048_445, w_048_448, w_048_450, w_048_458, w_048_479, w_048_490, w_048_493, w_048_517, w_048_519, w_048_525, w_048_542, w_048_552, w_048_559, w_048_575, w_048_591, w_048_595, w_048_599, w_048_605, w_048_606, w_048_620, w_048_673, w_048_679, w_048_694, w_048_706, w_048_732, w_048_734, w_048_738, w_048_748, w_048_780, w_048_801, w_048_803, w_048_816;
  wire w_049_003, w_049_018, w_049_041, w_049_044, w_049_069, w_049_071, w_049_075, w_049_078, w_049_147, w_049_190, w_049_192, w_049_194, w_049_210, w_049_217, w_049_218, w_049_220, w_049_245, w_049_246, w_049_247, w_049_250, w_049_259, w_049_270, w_049_298, w_049_307, w_049_309, w_049_321, w_049_327, w_049_329, w_049_334, w_049_338, w_049_341, w_049_343, w_049_358, w_049_363, w_049_383, w_049_397, w_049_412, w_049_414, w_049_445, w_049_454, w_049_459, w_049_470, w_049_478, w_049_516, w_049_521, w_049_525, w_049_534, w_049_541, w_049_548, w_049_587, w_049_602, w_049_607, w_049_619, w_049_623, w_049_629, w_049_633, w_049_649, w_049_651, w_049_654, w_049_657, w_049_690, w_049_691, w_049_706, w_049_739, w_049_742, w_049_750, w_049_786, w_049_797, w_049_828, w_049_835, w_049_855, w_049_879, w_049_883, w_049_886, w_049_913, w_049_925, w_049_930, w_049_936, w_049_943, w_049_944, w_049_965;
  wire w_050_002, w_050_003, w_050_005, w_050_035, w_050_037, w_050_038, w_050_039, w_050_044, w_050_058, w_050_059, w_050_068, w_050_083, w_050_086, w_050_088, w_050_100, w_050_102, w_050_111, w_050_141, w_050_147, w_050_152, w_050_159, w_050_166, w_050_186, w_050_192, w_050_195, w_050_198, w_050_200, w_050_215, w_050_229, w_050_231, w_050_237, w_050_244, w_050_247, w_050_248, w_050_250, w_050_255, w_050_264, w_050_282, w_050_289, w_050_294, w_050_299, w_050_301, w_050_311, w_050_322, w_050_323, w_050_344, w_050_353, w_050_361, w_050_365, w_050_366, w_050_369, w_050_370, w_050_371, w_050_376, w_050_386, w_050_389, w_050_395, w_050_396, w_050_401, w_050_407, w_050_409, w_050_413, w_050_423, w_050_438, w_050_469;
  wire w_051_002, w_051_023, w_051_031, w_051_037, w_051_046, w_051_047, w_051_050, w_051_060, w_051_066, w_051_069, w_051_071, w_051_075, w_051_094, w_051_102, w_051_108, w_051_114, w_051_115, w_051_118, w_051_123, w_051_129, w_051_134, w_051_138, w_051_142, w_051_161, w_051_165, w_051_167, w_051_178, w_051_179, w_051_184, w_051_196, w_051_204, w_051_223, w_051_240, w_051_249, w_051_255, w_051_286, w_051_288, w_051_290, w_051_299, w_051_306, w_051_307, w_051_308, w_051_313, w_051_314, w_051_317, w_051_318, w_051_320, w_051_327, w_051_336, w_051_339, w_051_342, w_051_356, w_051_360, w_051_370, w_051_372, w_051_381, w_051_382, w_051_384, w_051_392, w_051_404, w_051_409, w_051_413, w_051_417, w_051_420, w_051_438, w_051_439, w_051_457, w_051_517, w_051_527, w_051_540;
  wire w_052_002, w_052_004, w_052_006, w_052_007, w_052_008, w_052_009, w_052_012, w_052_013, w_052_015, w_052_016, w_052_017, w_052_022, w_052_023, w_052_026, w_052_029, w_052_030, w_052_031, w_052_034, w_052_035, w_052_036, w_052_037, w_052_041, w_052_046, w_052_049, w_052_051, w_052_053, w_052_058, w_052_059, w_052_060, w_052_062, w_052_064, w_052_067, w_052_068, w_052_071, w_052_073, w_052_078, w_052_080, w_052_082, w_052_099, w_052_100, w_052_101, w_052_102, w_052_106, w_052_108, w_052_109, w_052_115, w_052_117, w_052_120, w_052_121, w_052_125, w_052_126, w_052_128, w_052_129, w_052_132, w_052_133, w_052_135, w_052_137, w_052_143, w_052_144, w_052_145, w_052_147, w_052_148, w_052_150, w_052_152, w_052_153, w_052_160, w_052_162, w_052_164, w_052_165;
  wire w_053_002, w_053_005, w_053_012, w_053_019, w_053_022, w_053_030, w_053_036, w_053_042, w_053_053, w_053_055, w_053_058, w_053_069, w_053_070, w_053_081, w_053_089, w_053_092, w_053_102, w_053_109, w_053_112, w_053_145, w_053_151, w_053_175, w_053_181, w_053_193, w_053_230, w_053_236, w_053_238, w_053_289, w_053_292, w_053_297, w_053_300, w_053_310, w_053_341, w_053_346, w_053_364, w_053_377, w_053_388, w_053_391, w_053_400, w_053_404, w_053_425, w_053_437, w_053_456, w_053_492, w_053_515, w_053_526, w_053_528, w_053_533, w_053_551, w_053_562, w_053_575, w_053_582, w_053_587, w_053_592, w_053_616, w_053_645, w_053_647, w_053_654, w_053_655, w_053_676, w_053_677, w_053_707, w_053_729, w_053_733, w_053_735, w_053_760, w_053_763, w_053_816, w_053_824, w_053_835, w_053_837;
  wire w_054_008, w_054_009, w_054_014, w_054_015, w_054_016, w_054_017, w_054_020, w_054_023, w_054_029, w_054_034, w_054_035, w_054_041, w_054_054, w_054_058, w_054_060, w_054_077, w_054_079, w_054_080, w_054_081, w_054_084, w_054_085, w_054_086, w_054_089, w_054_102, w_054_110, w_054_112, w_054_116, w_054_126, w_054_128, w_054_134, w_054_141, w_054_147, w_054_152, w_054_160, w_054_163, w_054_165, w_054_167, w_054_170, w_054_179, w_054_180, w_054_185, w_054_191, w_054_195, w_054_196, w_054_200, w_054_201, w_054_203, w_054_209, w_054_210, w_054_214, w_054_215, w_054_216, w_054_217, w_054_218, w_054_221, w_054_227, w_054_234, w_054_240, w_054_246, w_054_249, w_054_251, w_054_253, w_054_255;
  wire w_055_000, w_055_001, w_055_010, w_055_011, w_055_017, w_055_022, w_055_033, w_055_035, w_055_055, w_055_065, w_055_071, w_055_080, w_055_081, w_055_105, w_055_129, w_055_138, w_055_159, w_055_163, w_055_174, w_055_176, w_055_183, w_055_192, w_055_194, w_055_210, w_055_223, w_055_233, w_055_245, w_055_250, w_055_261, w_055_311, w_055_319, w_055_336, w_055_358, w_055_375, w_055_398, w_055_474, w_055_500, w_055_503, w_055_529, w_055_548, w_055_574, w_055_593, w_055_594, w_055_596, w_055_603, w_055_607, w_055_611, w_055_615, w_055_664, w_055_688, w_055_723, w_055_731, w_055_732, w_055_744, w_055_762;
  wire w_056_003, w_056_004, w_056_007, w_056_010, w_056_012, w_056_022, w_056_034, w_056_039, w_056_045, w_056_048, w_056_065, w_056_077, w_056_081, w_056_086, w_056_088, w_056_092, w_056_096, w_056_099, w_056_112, w_056_125, w_056_128, w_056_166, w_056_170, w_056_175, w_056_177, w_056_187, w_056_188, w_056_190, w_056_193, w_056_196, w_056_212, w_056_219, w_056_227, w_056_228, w_056_231, w_056_235, w_056_236, w_056_255, w_056_256, w_056_275, w_056_279, w_056_280, w_056_284, w_056_285, w_056_299, w_056_311;
  wire w_057_002, w_057_008, w_057_010, w_057_017, w_057_021, w_057_023, w_057_024, w_057_031, w_057_039, w_057_041, w_057_043, w_057_050, w_057_051, w_057_063, w_057_067, w_057_091, w_057_092, w_057_102, w_057_113, w_057_121, w_057_122, w_057_145, w_057_154, w_057_157, w_057_167, w_057_169, w_057_190, w_057_198, w_057_200, w_057_202, w_057_209, w_057_210, w_057_233, w_057_252, w_057_253, w_057_256, w_057_262, w_057_275, w_057_305, w_057_311, w_057_316, w_057_322, w_057_323, w_057_325, w_057_336, w_057_337, w_057_350, w_057_353, w_057_357, w_057_385, w_057_393, w_057_397, w_057_403, w_057_415, w_057_417, w_057_425, w_057_435, w_057_443, w_057_445, w_057_467;
  wire w_058_002, w_058_006, w_058_009, w_058_010, w_058_015, w_058_040, w_058_050, w_058_058, w_058_064, w_058_065, w_058_070, w_058_071, w_058_072, w_058_080, w_058_085, w_058_086, w_058_094, w_058_097, w_058_108, w_058_112, w_058_115, w_058_123, w_058_128, w_058_139, w_058_140, w_058_151, w_058_154, w_058_155, w_058_167, w_058_172, w_058_176, w_058_177, w_058_179, w_058_182, w_058_190, w_058_191, w_058_196, w_058_197, w_058_199, w_058_205, w_058_215, w_058_220, w_058_221, w_058_225, w_058_227, w_058_233, w_058_238, w_058_239, w_058_247, w_058_250, w_058_281, w_058_292, w_058_302, w_058_317, w_058_320, w_058_324, w_058_335, w_058_341, w_058_347, w_058_360;
  wire w_059_018, w_059_028, w_059_030, w_059_032, w_059_044, w_059_047, w_059_058, w_059_068, w_059_076, w_059_090, w_059_092, w_059_094, w_059_097, w_059_105, w_059_116, w_059_121, w_059_123, w_059_134, w_059_135, w_059_138, w_059_142, w_059_143, w_059_145, w_059_146, w_059_147, w_059_149, w_059_151, w_059_152, w_059_154, w_059_164, w_059_169, w_059_177, w_059_179, w_059_180, w_059_192, w_059_193, w_059_209, w_059_213, w_059_214, w_059_224, w_059_230, w_059_235, w_059_237, w_059_245, w_059_247, w_059_258, w_059_263, w_059_264, w_059_272, w_059_277, w_059_278, w_059_279, w_059_282, w_059_308, w_059_317, w_059_318, w_059_333;
  wire w_060_012, w_060_018, w_060_024, w_060_035, w_060_057, w_060_071, w_060_095, w_060_101, w_060_105, w_060_120, w_060_134, w_060_142, w_060_153, w_060_155, w_060_165, w_060_171, w_060_173, w_060_178, w_060_183, w_060_185, w_060_189, w_060_212, w_060_213, w_060_215, w_060_229, w_060_240, w_060_241, w_060_242, w_060_246, w_060_247, w_060_249, w_060_257, w_060_260, w_060_263, w_060_269, w_060_288, w_060_297, w_060_301, w_060_305, w_060_307, w_060_311, w_060_313, w_060_316, w_060_320, w_060_323, w_060_331, w_060_341;
  wire w_061_009, w_061_017, w_061_023, w_061_033, w_061_034, w_061_045, w_061_052, w_061_055, w_061_063, w_061_069, w_061_070, w_061_071, w_061_078, w_061_095, w_061_123, w_061_132, w_061_147, w_061_168, w_061_172, w_061_174, w_061_216, w_061_221, w_061_222, w_061_235, w_061_238, w_061_241, w_061_245, w_061_247, w_061_250, w_061_254, w_061_255, w_061_257, w_061_267, w_061_283, w_061_286, w_061_298, w_061_300, w_061_331, w_061_333, w_061_355, w_061_360, w_061_377, w_061_379, w_061_380, w_061_394, w_061_403, w_061_410, w_061_414, w_061_432, w_061_433, w_061_461, w_061_478, w_061_490, w_061_497, w_061_502, w_061_528, w_061_560;
  wire w_062_021, w_062_022, w_062_029, w_062_031, w_062_032, w_062_037, w_062_069, w_062_100, w_062_121, w_062_124, w_062_140, w_062_149, w_062_165, w_062_166, w_062_167, w_062_174, w_062_228, w_062_240, w_062_251, w_062_252, w_062_253, w_062_272, w_062_280, w_062_292, w_062_300, w_062_312, w_062_314, w_062_353, w_062_371, w_062_373, w_062_374, w_062_386, w_062_428, w_062_432, w_062_436, w_062_440, w_062_469, w_062_471, w_062_474, w_062_478, w_062_479;
  wire w_063_027, w_063_037, w_063_038, w_063_053, w_063_054, w_063_059, w_063_064, w_063_071, w_063_081, w_063_083, w_063_084, w_063_085, w_063_098, w_063_099, w_063_103, w_063_104, w_063_107, w_063_110, w_063_119, w_063_130, w_063_133, w_063_135, w_063_138, w_063_146, w_063_162, w_063_181, w_063_193, w_063_195, w_063_198, w_063_200, w_063_201, w_063_204, w_063_205, w_063_210, w_063_212, w_063_215, w_063_216, w_063_217, w_063_225, w_063_226, w_063_231, w_063_242, w_063_258, w_063_260, w_063_266, w_063_274, w_063_286, w_063_287, w_063_290, w_063_293, w_063_303, w_063_315, w_063_322, w_063_353, w_063_357, w_063_360;
  wire w_064_002, w_064_003, w_064_021, w_064_032, w_064_036, w_064_041, w_064_070, w_064_076, w_064_086, w_064_091, w_064_102, w_064_131, w_064_138, w_064_142, w_064_146, w_064_157, w_064_169, w_064_188, w_064_247, w_064_264, w_064_271, w_064_277, w_064_311, w_064_338, w_064_340, w_064_347, w_064_355, w_064_375, w_064_411, w_064_433, w_064_448, w_064_453, w_064_477, w_064_482, w_064_493, w_064_503, w_064_515, w_064_526, w_064_534, w_064_537, w_064_554, w_064_574, w_064_606, w_064_610, w_064_630, w_064_637, w_064_665, w_064_668, w_064_679, w_064_690, w_064_692, w_064_695, w_064_727, w_064_741, w_064_749, w_064_750, w_064_789, w_064_804, w_064_806, w_064_832;
  wire w_065_006, w_065_013, w_065_017, w_065_051, w_065_091, w_065_094, w_065_095, w_065_160, w_065_204, w_065_223, w_065_251, w_065_279, w_065_305, w_065_312, w_065_333, w_065_363, w_065_373, w_065_380, w_065_422, w_065_423, w_065_433, w_065_509, w_065_527, w_065_537, w_065_551, w_065_556, w_065_585, w_065_613, w_065_631, w_065_652, w_065_665, w_065_686, w_065_697, w_065_711, w_065_732, w_065_740, w_065_742, w_065_750, w_065_850, w_065_855, w_065_861, w_065_883, w_065_895, w_065_914, w_065_920, w_065_941, w_065_944, w_065_950, w_065_951, w_065_972, w_065_978;
  wire w_066_014, w_066_017, w_066_023, w_066_024, w_066_037, w_066_039, w_066_051, w_066_054, w_066_058, w_066_072, w_066_082, w_066_107, w_066_114, w_066_115, w_066_119, w_066_124, w_066_141, w_066_146, w_066_187, w_066_202, w_066_209, w_066_210, w_066_213, w_066_224, w_066_249, w_066_282, w_066_285, w_066_295, w_066_317, w_066_345, w_066_355, w_066_359, w_066_368, w_066_371, w_066_376, w_066_392, w_066_399, w_066_400, w_066_414, w_066_465, w_066_475, w_066_476, w_066_485, w_066_493, w_066_511;
  wire w_067_029, w_067_075, w_067_077, w_067_085, w_067_121, w_067_148, w_067_151, w_067_168, w_067_178, w_067_200, w_067_216, w_067_218, w_067_224, w_067_226, w_067_229, w_067_242, w_067_245, w_067_251, w_067_263, w_067_265, w_067_283, w_067_294, w_067_334, w_067_343, w_067_363, w_067_444, w_067_508, w_067_516, w_067_615, w_067_649, w_067_711, w_067_724, w_067_728, w_067_746, w_067_754, w_067_785, w_067_786, w_067_804, w_067_816, w_067_866, w_067_880, w_067_905, w_067_920, w_067_921, w_067_939, w_067_945;
  wire w_068_005, w_068_010, w_068_011, w_068_013, w_068_018, w_068_024, w_068_025, w_068_039, w_068_049, w_068_056, w_068_068, w_068_069, w_068_081, w_068_091, w_068_093, w_068_108, w_068_128, w_068_138, w_068_141, w_068_145, w_068_150, w_068_157, w_068_171, w_068_175, w_068_178, w_068_187, w_068_191, w_068_194, w_068_198, w_068_203, w_068_212, w_068_219, w_068_234, w_068_256, w_068_258, w_068_275, w_068_283, w_068_302, w_068_303, w_068_306, w_068_307, w_068_309, w_068_313, w_068_315, w_068_327, w_068_329;
  wire w_069_000, w_069_004, w_069_005, w_069_014, w_069_017, w_069_018, w_069_022, w_069_024, w_069_029, w_069_033, w_069_058, w_069_067, w_069_070, w_069_081, w_069_084, w_069_107, w_069_108, w_069_114, w_069_125, w_069_126, w_069_137, w_069_139, w_069_143, w_069_144, w_069_145, w_069_146, w_069_149, w_069_151, w_069_159, w_069_163;
  wire w_070_026, w_070_027, w_070_053, w_070_117, w_070_147, w_070_154, w_070_204, w_070_234, w_070_256, w_070_261, w_070_289, w_070_346, w_070_356, w_070_381, w_070_388, w_070_403, w_070_446, w_070_464, w_070_484, w_070_488, w_070_493, w_070_528, w_070_530, w_070_551, w_070_552, w_070_595, w_070_629, w_070_647, w_070_659, w_070_699, w_070_702, w_070_712, w_070_730, w_070_748, w_070_752, w_070_784, w_070_792, w_070_823, w_070_829, w_070_847, w_070_864, w_070_888, w_070_915, w_070_926, w_070_935;
  wire w_071_003, w_071_007, w_071_011, w_071_016, w_071_040, w_071_041, w_071_046, w_071_057, w_071_058, w_071_060, w_071_071, w_071_076, w_071_079, w_071_095, w_071_112, w_071_115, w_071_116, w_071_125, w_071_129, w_071_134, w_071_137, w_071_147, w_071_151, w_071_158, w_071_166, w_071_174, w_071_206, w_071_207, w_071_225, w_071_230, w_071_233, w_071_239, w_071_246, w_071_249, w_071_250, w_071_253, w_071_276, w_071_281, w_071_284, w_071_286, w_071_306, w_071_312, w_071_329, w_071_337, w_071_351, w_071_363, w_071_366, w_071_400, w_071_428, w_071_431, w_071_434, w_071_436, w_071_447;
  wire w_072_000, w_072_002, w_072_003, w_072_004, w_072_006, w_072_007, w_072_008, w_072_010, w_072_011, w_072_013, w_072_014, w_072_015, w_072_016, w_072_017, w_072_019, w_072_020, w_072_021, w_072_022, w_072_023, w_072_024, w_072_026, w_072_029, w_072_030, w_072_031, w_072_032, w_072_033, w_072_034, w_072_037, w_072_038, w_072_040, w_072_041, w_072_042, w_072_046, w_072_048, w_072_049, w_072_052, w_072_054, w_072_055, w_072_057, w_072_060, w_072_063, w_072_065, w_072_067;
  wire w_073_005, w_073_012, w_073_021, w_073_030, w_073_034, w_073_059, w_073_073, w_073_090, w_073_092, w_073_095, w_073_114, w_073_117, w_073_123, w_073_156, w_073_160, w_073_214, w_073_292, w_073_322, w_073_323, w_073_331, w_073_339, w_073_409, w_073_411, w_073_413, w_073_416, w_073_430, w_073_452, w_073_479, w_073_490, w_073_506, w_073_540, w_073_550, w_073_643, w_073_645, w_073_655, w_073_663, w_073_704, w_073_705, w_073_747, w_073_766, w_073_804, w_073_818;
  wire w_074_003, w_074_048, w_074_061, w_074_067, w_074_156, w_074_214, w_074_254, w_074_258, w_074_261, w_074_273, w_074_294, w_074_297, w_074_316, w_074_328, w_074_342, w_074_358, w_074_366, w_074_378, w_074_383, w_074_463, w_074_467, w_074_479, w_074_488, w_074_531, w_074_532, w_074_588, w_074_607, w_074_633, w_074_681, w_074_691, w_074_692, w_074_751, w_074_754, w_074_787, w_074_846, w_074_847, w_074_909, w_074_915, w_074_931, w_074_944, w_074_963;
  wire w_075_008, w_075_016, w_075_024, w_075_029, w_075_036, w_075_043, w_075_051, w_075_052, w_075_069, w_075_082, w_075_089, w_075_100, w_075_101, w_075_103, w_075_108, w_075_111, w_075_114, w_075_144, w_075_179, w_075_180, w_075_188, w_075_189, w_075_192, w_075_199, w_075_229, w_075_258, w_075_260, w_075_284, w_075_285;
  wire w_076_006, w_076_008, w_076_012, w_076_044, w_076_053, w_076_056, w_076_102, w_076_107, w_076_136, w_076_142, w_076_166, w_076_175, w_076_192, w_076_220, w_076_227, w_076_236, w_076_245, w_076_269, w_076_273, w_076_310, w_076_324, w_076_330, w_076_336, w_076_342, w_076_352, w_076_356, w_076_360, w_076_363, w_076_388, w_076_393, w_076_417, w_076_422, w_076_433, w_076_437, w_076_449, w_076_582, w_076_591, w_076_616, w_076_617;
  wire w_077_012, w_077_016, w_077_018, w_077_028, w_077_041, w_077_047, w_077_069, w_077_074, w_077_083, w_077_098, w_077_100, w_077_101, w_077_104, w_077_107, w_077_108, w_077_112, w_077_121, w_077_191, w_077_193, w_077_194, w_077_197, w_077_219, w_077_240, w_077_266, w_077_281, w_077_301, w_077_317, w_077_321, w_077_323, w_077_347, w_077_381, w_077_385, w_077_400, w_077_410, w_077_419, w_077_430, w_077_443, w_077_449, w_077_472, w_077_491;
  wire w_078_007, w_078_009, w_078_017, w_078_020, w_078_028, w_078_034, w_078_042, w_078_044, w_078_049, w_078_051, w_078_053, w_078_055, w_078_073, w_078_077, w_078_087, w_078_090, w_078_102, w_078_121, w_078_132, w_078_151, w_078_161, w_078_189, w_078_199, w_078_201, w_078_203, w_078_209, w_078_211, w_078_212, w_078_221, w_078_228, w_078_233, w_078_240, w_078_251, w_078_265, w_078_271, w_078_287, w_078_288, w_078_292, w_078_297, w_078_302;
  wire w_079_000, w_079_004, w_079_015, w_079_021, w_079_046, w_079_051, w_079_068, w_079_074, w_079_078, w_079_084, w_079_086, w_079_112, w_079_114, w_079_121, w_079_129, w_079_130, w_079_136, w_079_146, w_079_150, w_079_162, w_079_163, w_079_172, w_079_182, w_079_199, w_079_218, w_079_219, w_079_228, w_079_231, w_079_234, w_079_244, w_079_247;
  wire w_080_008, w_080_009, w_080_010, w_080_011, w_080_016, w_080_022, w_080_026, w_080_028, w_080_030, w_080_031, w_080_032, w_080_038, w_080_043, w_080_046, w_080_056, w_080_058, w_080_059, w_080_061, w_080_063, w_080_064, w_080_071, w_080_075, w_080_080, w_080_086, w_080_092, w_080_093, w_080_099, w_080_102, w_080_103, w_080_104, w_080_107, w_080_108, w_080_112, w_080_114;
  wire w_081_016, w_081_017, w_081_026, w_081_041, w_081_060, w_081_083, w_081_084, w_081_090, w_081_119, w_081_122, w_081_134, w_081_139, w_081_170, w_081_212, w_081_237, w_081_240, w_081_252, w_081_270, w_081_294, w_081_360, w_081_374, w_081_383, w_081_384, w_081_458, w_081_478, w_081_527, w_081_538, w_081_563, w_081_567, w_081_582, w_081_590;
  wire w_082_004, w_082_013, w_082_015, w_082_027, w_082_028, w_082_029, w_082_033, w_082_061, w_082_063, w_082_097, w_082_146, w_082_158, w_082_163, w_082_194, w_082_197, w_082_206, w_082_212, w_082_217, w_082_218, w_082_222, w_082_228, w_082_231, w_082_232, w_082_240, w_082_248, w_082_253, w_082_257, w_082_258, w_082_266, w_082_285, w_082_301, w_082_321, w_082_323, w_082_330, w_082_334, w_082_342, w_082_344;
  wire w_083_000, w_083_021, w_083_022, w_083_023, w_083_030, w_083_068, w_083_079, w_083_087, w_083_095, w_083_109, w_083_111, w_083_137, w_083_138, w_083_147, w_083_153, w_083_158, w_083_164, w_083_173, w_083_220, w_083_224, w_083_238, w_083_240, w_083_242, w_083_249, w_083_253, w_083_259, w_083_266, w_083_274, w_083_291, w_083_302, w_083_310, w_083_435, w_083_439, w_083_441, w_083_453, w_083_596, w_083_597, w_083_618, w_083_619, w_083_649, w_083_651, w_083_653;
  wire w_084_012, w_084_029, w_084_033, w_084_035, w_084_039, w_084_050, w_084_062, w_084_074, w_084_114, w_084_122, w_084_125, w_084_128, w_084_131, w_084_148, w_084_169, w_084_190, w_084_208, w_084_231, w_084_234, w_084_240, w_084_257, w_084_268, w_084_294, w_084_299, w_084_329, w_084_428, w_084_494, w_084_526, w_084_535, w_084_567, w_084_610;
  wire w_085_000, w_085_003, w_085_004, w_085_006, w_085_008, w_085_010, w_085_011, w_085_013, w_085_016, w_085_017, w_085_019, w_085_020, w_085_021, w_085_022, w_085_023, w_085_024, w_085_026, w_085_027, w_085_037, w_085_039, w_085_041, w_085_043, w_085_044, w_085_050, w_085_051, w_085_054, w_085_055, w_085_056, w_085_057, w_085_058, w_085_059, w_085_060, w_085_070, w_085_071;
  wire w_086_001, w_086_006, w_086_012, w_086_017, w_086_026, w_086_059, w_086_060, w_086_077, w_086_090, w_086_099, w_086_106, w_086_116, w_086_143, w_086_167, w_086_182, w_086_202, w_086_215, w_086_222, w_086_242, w_086_358, w_086_364, w_086_395, w_086_408, w_086_415, w_086_427, w_086_428, w_086_482, w_086_577, w_086_590, w_086_596, w_086_642, w_086_652, w_086_659, w_086_666, w_086_668, w_086_701, w_086_705, w_086_709, w_086_720, w_086_721, w_086_725, w_086_745, w_086_750, w_086_776;
  wire w_087_024, w_087_039, w_087_040, w_087_044, w_087_049, w_087_052, w_087_053, w_087_059, w_087_069, w_087_080, w_087_109, w_087_135, w_087_144, w_087_145, w_087_147, w_087_177, w_087_195, w_087_220, w_087_226, w_087_256, w_087_263, w_087_304, w_087_313, w_087_329, w_087_348;
  wire w_088_030, w_088_037, w_088_063, w_088_077, w_088_098, w_088_108, w_088_151, w_088_163, w_088_179, w_088_189, w_088_193, w_088_207, w_088_214, w_088_230, w_088_285, w_088_379, w_088_404, w_088_458, w_088_500, w_088_533, w_088_534, w_088_618, w_088_619, w_088_655, w_088_695;
  wire w_089_006, w_089_009, w_089_015, w_089_018, w_089_019, w_089_022, w_089_024, w_089_031, w_089_056, w_089_068, w_089_074, w_089_078, w_089_079, w_089_082, w_089_088, w_089_090, w_089_091, w_089_095, w_089_098, w_089_107, w_089_113, w_089_127, w_089_135;
  wire w_090_003, w_090_019, w_090_026, w_090_038, w_090_048, w_090_066, w_090_079, w_090_086, w_090_121, w_090_127, w_090_139, w_090_160, w_090_200, w_090_205, w_090_209, w_090_212, w_090_220, w_090_224, w_090_238, w_090_244, w_090_250, w_090_252, w_090_268, w_090_270, w_090_271, w_090_281, w_090_283, w_090_295, w_090_297, w_090_328, w_090_332, w_090_335, w_090_336, w_090_337, w_090_384, w_090_393;
  wire w_091_000, w_091_002, w_091_031, w_091_036, w_091_048, w_091_068, w_091_082, w_091_125, w_091_127, w_091_145, w_091_150, w_091_170, w_091_173, w_091_179, w_091_182, w_091_186, w_091_190, w_091_206, w_091_214, w_091_232, w_091_233, w_091_279, w_091_316, w_091_347, w_091_403, w_091_408, w_091_507, w_091_552, w_091_555;
  wire w_092_011, w_092_033, w_092_034, w_092_037, w_092_038, w_092_043, w_092_083, w_092_092, w_092_122, w_092_129, w_092_130, w_092_138, w_092_210, w_092_239, w_092_282, w_092_461, w_092_503, w_092_524, w_092_546, w_092_644, w_092_680, w_092_706, w_092_747;
  wire w_093_015, w_093_107, w_093_111, w_093_130, w_093_137, w_093_169, w_093_200, w_093_203, w_093_227, w_093_241, w_093_258, w_093_279, w_093_320, w_093_346, w_093_353, w_093_374, w_093_423, w_093_484, w_093_600, w_093_720, w_093_734, w_093_769, w_093_791, w_093_825, w_093_858, w_093_878, w_093_911, w_093_915, w_093_919;
  wire w_094_011, w_094_028, w_094_055, w_094_078, w_094_113, w_094_115, w_094_124, w_094_134, w_094_150, w_094_169, w_094_208, w_094_217, w_094_292, w_094_313, w_094_415, w_094_506, w_094_671, w_094_710, w_094_726, w_094_763, w_094_781, w_094_794, w_094_817, w_094_869, w_094_884;
  wire w_095_000, w_095_002, w_095_008, w_095_009, w_095_017, w_095_019, w_095_022, w_095_028, w_095_030, w_095_040, w_095_054, w_095_074, w_095_081, w_095_094, w_095_101, w_095_108, w_095_112, w_095_115, w_095_128, w_095_131, w_095_149, w_095_150, w_095_153, w_095_163, w_095_164, w_095_165, w_095_181, w_095_182;
  wire w_096_028, w_096_075, w_096_086, w_096_097, w_096_100, w_096_108, w_096_114, w_096_118, w_096_120, w_096_124, w_096_130, w_096_131, w_096_139, w_096_160, w_096_168, w_096_185, w_096_218, w_096_229, w_096_248, w_096_254, w_096_255, w_096_293, w_096_299, w_096_346, w_096_348, w_096_380, w_096_381, w_096_419, w_096_475, w_096_566, w_096_581, w_096_628, w_096_629, w_096_630, w_096_631, w_096_632, w_096_633, w_096_634, w_096_635, w_096_636, w_096_637, w_096_638, w_096_642, w_096_643, w_096_644, w_096_645, w_096_646, w_096_647, w_096_648, w_096_649, w_096_650, w_096_651, w_096_653;
  wire w_097_001, w_097_030, w_097_038, w_097_041, w_097_045, w_097_054, w_097_057, w_097_058, w_097_069, w_097_073, w_097_077, w_097_141, w_097_171, w_097_183, w_097_192, w_097_228, w_097_231, w_097_260, w_097_329, w_097_441, w_097_495, w_097_501, w_097_502, w_097_513, w_097_583, w_097_595, w_097_602, w_097_634, w_097_636;
  wire w_098_025, w_098_035, w_098_036, w_098_048, w_098_079, w_098_095, w_098_189, w_098_222, w_098_231, w_098_257, w_098_278, w_098_310, w_098_315, w_098_329, w_098_341, w_098_410, w_098_422, w_098_450, w_098_451, w_098_465;
  wire w_099_006, w_099_020, w_099_035, w_099_036, w_099_038, w_099_059, w_099_070, w_099_077, w_099_082, w_099_085, w_099_102, w_099_105, w_099_114, w_099_120, w_099_128, w_099_130, w_099_157, w_099_158, w_099_171, w_099_181, w_099_182, w_099_183, w_099_187, w_099_194, w_099_196, w_099_205, w_099_210, w_099_230, w_099_231, w_099_234;
  wire w_100_045, w_100_104, w_100_160, w_100_171, w_100_172, w_100_174, w_100_201, w_100_202, w_100_225, w_100_257, w_100_283, w_100_305, w_100_313, w_100_335, w_100_368, w_100_392, w_100_414, w_100_429, w_100_533, w_100_556, w_100_565, w_100_608, w_100_626, w_100_642, w_100_657, w_100_754, w_100_756, w_100_819, w_100_847, w_100_914, w_100_926;
  wire w_101_002, w_101_012, w_101_016, w_101_043, w_101_047, w_101_055, w_101_066, w_101_081, w_101_083, w_101_094, w_101_106, w_101_120, w_101_122, w_101_128, w_101_130, w_101_133, w_101_141, w_101_143, w_101_144, w_101_148, w_101_152, w_101_153, w_101_159, w_101_176, w_101_185;
  wire w_102_004, w_102_031, w_102_070, w_102_094, w_102_124, w_102_155, w_102_159, w_102_160, w_102_162, w_102_195, w_102_215, w_102_233, w_102_298, w_102_381, w_102_400, w_102_450, w_102_563, w_102_571, w_102_610, w_102_611, w_102_676, w_102_678, w_102_721, w_102_750, w_102_754, w_102_779;
  wire w_103_011, w_103_040, w_103_049, w_103_057, w_103_063, w_103_160, w_103_236, w_103_246, w_103_271, w_103_302, w_103_306, w_103_361, w_103_444, w_103_447, w_103_498, w_103_582, w_103_640, w_103_649, w_103_658, w_103_663, w_103_765, w_103_791, w_103_812, w_103_825, w_103_843, w_103_848, w_103_894;
  wire w_104_012, w_104_013, w_104_019, w_104_024, w_104_035, w_104_036, w_104_038, w_104_042, w_104_062, w_104_091, w_104_108, w_104_116, w_104_122, w_104_140, w_104_159, w_104_169, w_104_176, w_104_180, w_104_225, w_104_233, w_104_246, w_104_250;
  wire w_105_017, w_105_029, w_105_038, w_105_044, w_105_117, w_105_189, w_105_190, w_105_198, w_105_219, w_105_249, w_105_255, w_105_342, w_105_346, w_105_380, w_105_397, w_105_467, w_105_486, w_105_498, w_105_533, w_105_626, w_105_701, w_105_718, w_105_787, w_105_827, w_105_852, w_105_855, w_105_891;
  wire w_106_008, w_106_016, w_106_018, w_106_049, w_106_103, w_106_115, w_106_137, w_106_141, w_106_167, w_106_205, w_106_224, w_106_237, w_106_253, w_106_291, w_106_299, w_106_302, w_106_334, w_106_418, w_106_438, w_106_512, w_106_622, w_106_642;
  wire w_107_013, w_107_014, w_107_016, w_107_018, w_107_019, w_107_021, w_107_022, w_107_025, w_107_027, w_107_030, w_107_038, w_107_046, w_107_050, w_107_072, w_107_077, w_107_082, w_107_088, w_107_100, w_107_110, w_107_115, w_107_126, w_107_127, w_107_128, w_107_141, w_107_145, w_107_147, w_107_165, w_107_169, w_107_180, w_107_181, w_107_182, w_107_190, w_107_197, w_107_203, w_107_206;
  wire w_108_000, w_108_001, w_108_002, w_108_003, w_108_005, w_108_006, w_108_007, w_108_008, w_108_009, w_108_011;
  wire w_109_005, w_109_019, w_109_040, w_109_048, w_109_049, w_109_058, w_109_068, w_109_083, w_109_130, w_109_133, w_109_142, w_109_145, w_109_147, w_109_150, w_109_153, w_109_167, w_109_169, w_109_178, w_109_232, w_109_257, w_109_259, w_109_268, w_109_275, w_109_283;
  wire w_110_005, w_110_010, w_110_041, w_110_051, w_110_053, w_110_090, w_110_095, w_110_123, w_110_143, w_110_179, w_110_195, w_110_232, w_110_303, w_110_347, w_110_350, w_110_404, w_110_414, w_110_455, w_110_486, w_110_581, w_110_647, w_110_663, w_110_664;
  wire w_111_018, w_111_028, w_111_031, w_111_044, w_111_048, w_111_062, w_111_071, w_111_082, w_111_092, w_111_101, w_111_140, w_111_146, w_111_162, w_111_183, w_111_196, w_111_202, w_111_206, w_111_238, w_111_291, w_111_312, w_111_339;
  wire w_112_013, w_112_029, w_112_048, w_112_049, w_112_060, w_112_063, w_112_067, w_112_071, w_112_082, w_112_086, w_112_087, w_112_088, w_112_089, w_112_092, w_112_095;
  wire w_113_019, w_113_041, w_113_070, w_113_080, w_113_155, w_113_167, w_113_185, w_113_210, w_113_220, w_113_223, w_113_239, w_113_248, w_113_299, w_113_304, w_113_305, w_113_322, w_113_331, w_113_351, w_113_372, w_113_423, w_113_428, w_113_453, w_113_455, w_113_515, w_113_524, w_113_548, w_113_629;
  wire w_114_006, w_114_010, w_114_024, w_114_025, w_114_048, w_114_058, w_114_059, w_114_113, w_114_132, w_114_136, w_114_187, w_114_190, w_114_231, w_114_283, w_114_286, w_114_295, w_114_302, w_114_303, w_114_318, w_114_356, w_114_366;
  wire w_115_003, w_115_019, w_115_021, w_115_025, w_115_030, w_115_031, w_115_034, w_115_036, w_115_037, w_115_045, w_115_046, w_115_057, w_115_062, w_115_069, w_115_071, w_115_073, w_115_075, w_115_079, w_115_084, w_115_086, w_115_089;
  wire w_116_007, w_116_011, w_116_013, w_116_014, w_116_018, w_116_023, w_116_027, w_116_032, w_116_034, w_116_035, w_116_037, w_116_038, w_116_040, w_116_041;
  wire w_117_015, w_117_080, w_117_081, w_117_082, w_117_087, w_117_100, w_117_105, w_117_112, w_117_135, w_117_148, w_117_156, w_117_184, w_117_185, w_117_193, w_117_196, w_117_240, w_117_247, w_117_263, w_117_283, w_117_287, w_117_290, w_117_313, w_117_315, w_117_324;
  wire w_118_035, w_118_085, w_118_091, w_118_102, w_118_112, w_118_142, w_118_160, w_118_180, w_118_181, w_118_184, w_118_190, w_118_192, w_118_211, w_118_217, w_118_234, w_118_245, w_118_258, w_118_288, w_118_291, w_118_295, w_118_325, w_118_347, w_118_350, w_118_360, w_118_384, w_118_447, w_118_580;
  wire w_119_046, w_119_051, w_119_080, w_119_117, w_119_119, w_119_121, w_119_140, w_119_148, w_119_189, w_119_190, w_119_202, w_119_221, w_119_238, w_119_285, w_119_297, w_119_299, w_119_361, w_119_363, w_119_368, w_119_406, w_119_408, w_119_419, w_119_517, w_119_561, w_119_575;
  wire w_120_005, w_120_013, w_120_016, w_120_018, w_120_021, w_120_032, w_120_035, w_120_045, w_120_055, w_120_066, w_120_068, w_120_078, w_120_087, w_120_097, w_120_102, w_120_110, w_120_111;
  wire w_121_003, w_121_077, w_121_081, w_121_124, w_121_174, w_121_175, w_121_178, w_121_182, w_121_260, w_121_301, w_121_331, w_121_354, w_121_384, w_121_470, w_121_484, w_121_485, w_121_557, w_121_590, w_121_610, w_121_637;
  wire w_122_066, w_122_069, w_122_088, w_122_135, w_122_137, w_122_208, w_122_256, w_122_268, w_122_270, w_122_278, w_122_281, w_122_302, w_122_309, w_122_348, w_122_366, w_122_385, w_122_399, w_122_436, w_122_447, w_122_458, w_122_472;
  wire w_123_011, w_123_025, w_123_027, w_123_048, w_123_062, w_123_066, w_123_073, w_123_080, w_123_090, w_123_129, w_123_160, w_123_168, w_123_191;
  wire w_124_071, w_124_091, w_124_128, w_124_134, w_124_142, w_124_157, w_124_235, w_124_283, w_124_305, w_124_470, w_124_649, w_124_697, w_124_701;
  wire w_125_007, w_125_019, w_125_022, w_125_032, w_125_054, w_125_089, w_125_092, w_125_101, w_125_124, w_125_129, w_125_181, w_125_186, w_125_190, w_125_199, w_125_207, w_125_213;
  wire w_126_034, w_126_053, w_126_112, w_126_118, w_126_141, w_126_166, w_126_241, w_126_251, w_126_280, w_126_304, w_126_385, w_126_398, w_126_461, w_126_484, w_126_517;
  wire w_127_023, w_127_029, w_127_065, w_127_068, w_127_071, w_127_076, w_127_077, w_127_085, w_127_095, w_127_109, w_127_116, w_127_130, w_127_141;
  wire w_128_003, w_128_004, w_128_005, w_128_024, w_128_027, w_128_075, w_128_081, w_128_094, w_128_103, w_128_116, w_128_125, w_128_133, w_128_146, w_128_149, w_128_162, w_128_179, w_128_199, w_128_201, w_128_202, w_128_203, w_128_208, w_128_216, w_128_217, w_128_220, w_128_239, w_128_240, w_128_243;
  wire w_129_000, w_129_001, w_129_004, w_129_006, w_129_008, w_129_011, w_129_016, w_129_022, w_129_024;
  wire w_130_002, w_130_104, w_130_213, w_130_262, w_130_269, w_130_271, w_130_291, w_130_340, w_130_422, w_130_545, w_130_620, w_130_661, w_130_726, w_130_747, w_130_767, w_130_860, w_130_866, w_130_882, w_130_917, w_130_922, w_130_925;
  wire w_131_028, w_131_070, w_131_081, w_131_082, w_131_094, w_131_100, w_131_116, w_131_120, w_131_121, w_131_181, w_131_185, w_131_578, w_131_617, w_131_632, w_131_634, w_131_682, w_131_685;
  wire w_132_033, w_132_145, w_132_160, w_132_166, w_132_192, w_132_288, w_132_300, w_132_338, w_132_353, w_132_367, w_132_383, w_132_529;
  wire w_133_010, w_133_016, w_133_024, w_133_057, w_133_086, w_133_097, w_133_158, w_133_177, w_133_236, w_133_252, w_133_266, w_133_298, w_133_327, w_133_374, w_133_416, w_133_430, w_133_516, w_133_521, w_133_559, w_133_790;
  wire w_134_003, w_134_010, w_134_097, w_134_127, w_134_203, w_134_205, w_134_252, w_134_267, w_134_285, w_134_291, w_134_326;
  wire w_135_006, w_135_009, w_135_020, w_135_047, w_135_054, w_135_064, w_135_072, w_135_074, w_135_083, w_135_105, w_135_123, w_135_139, w_135_203, w_135_204, w_135_207, w_135_219, w_135_221, w_135_226;
  wire w_136_012, w_136_037, w_136_049, w_136_050, w_136_052, w_136_093, w_136_133, w_136_307, w_136_319, w_136_504, w_136_588, w_136_694, w_136_920;
  wire w_137_009, w_137_019, w_137_044, w_137_068, w_137_119, w_137_150, w_137_165, w_137_199, w_137_202, w_137_249, w_137_265, w_137_297, w_137_383, w_137_394, w_137_424, w_137_478, w_137_554, w_137_579, w_137_594, w_137_613, w_137_643;
  wire w_138_021, w_138_023, w_138_061, w_138_065, w_138_084, w_138_127, w_138_145, w_138_147, w_138_183, w_138_187, w_138_191, w_138_192, w_138_261, w_138_269, w_138_416, w_138_465, w_138_569, w_138_674, w_138_690, w_138_693, w_138_726, w_138_738;
  wire w_139_001, w_139_002, w_139_003, w_139_005, w_139_006, w_139_007, w_139_009, w_139_012, w_139_013;
  wire w_140_051, w_140_101, w_140_150, w_140_219, w_140_273, w_140_280, w_140_284, w_140_289, w_140_308, w_140_319, w_140_333, w_140_630;
  wire w_141_052, w_141_061, w_141_078, w_141_088, w_141_342, w_141_358, w_141_409, w_141_465, w_141_610, w_141_673, w_141_706, w_141_707, w_141_726, w_141_823;
  wire w_142_011, w_142_062, w_142_087, w_142_130, w_142_158, w_142_208, w_142_340, w_142_493, w_142_567, w_142_598;
  wire w_143_002, w_143_055, w_143_115, w_143_129, w_143_159, w_143_241, w_143_253, w_143_256, w_143_279, w_143_311, w_143_328, w_143_356, w_143_402, w_143_418, w_143_510, w_143_549, w_143_576, w_143_577, w_143_578;
  wire w_144_022, w_144_097, w_144_128, w_144_131, w_144_158, w_144_234, w_144_282, w_144_289, w_144_299, w_144_323, w_144_347, w_144_394, w_144_412, w_144_417;
  wire w_145_008, w_145_017, w_145_023, w_145_029, w_145_030, w_145_046, w_145_047, w_145_050, w_145_052, w_145_054, w_145_059, w_145_062, w_145_091, w_145_097;
  wire w_146_012, w_146_065, w_146_073, w_146_106, w_146_122, w_146_124, w_146_129, w_146_170, w_146_196, w_146_222, w_146_224, w_146_231, w_146_264, w_146_274, w_146_296, w_146_314, w_146_328;
  wire w_147_047, w_147_085, w_147_125, w_147_140, w_147_152, w_147_189, w_147_213, w_147_263, w_147_269, w_147_338, w_147_491, w_147_520;
  wire w_148_028, w_148_102, w_148_111, w_148_280, w_148_311, w_148_327, w_148_364, w_148_371, w_148_379, w_148_417, w_148_429, w_148_441, w_148_444, w_148_460, w_148_495;
  wire w_149_065, w_149_069, w_149_145, w_149_161, w_149_232, w_149_239, w_149_266, w_149_315, w_149_353, w_149_355, w_149_392, w_149_449, w_149_546, w_149_559, w_149_707;
  wire w_150_043, w_150_122, w_150_140, w_150_154, w_150_160, w_150_194;
  wire w_151_000, w_151_003, w_151_034, w_151_109, w_151_196, w_151_210, w_151_223, w_151_226, w_151_246, w_151_249, w_151_255, w_151_282, w_151_283, w_151_288, w_151_298, w_151_307;
  wire w_152_042, w_152_059, w_152_087, w_152_116, w_152_130, w_152_278, w_152_395, w_152_422, w_152_460, w_152_476, w_152_479, w_152_505, w_152_611, w_152_621, w_152_632, w_152_696, w_152_770, w_152_771, w_152_772, w_152_773, w_152_774, w_152_775, w_152_779, w_152_780, w_152_781, w_152_782, w_152_783, w_152_784, w_152_786;
  wire w_153_056, w_153_072, w_153_114, w_153_152, w_153_177, w_153_210, w_153_385, w_153_415, w_153_457, w_153_471;
  wire w_154_004, w_154_083, w_154_113, w_154_137, w_154_148, w_154_154, w_154_243, w_154_297, w_154_555, w_154_563, w_154_586, w_154_799;
  wire w_155_011, w_155_013, w_155_027, w_155_054, w_155_061, w_155_079, w_155_108, w_155_109, w_155_124;
  wire w_156_092, w_156_302, w_156_315, w_156_422, w_156_456, w_156_622, w_156_661, w_156_708, w_156_709, w_156_710, w_156_711, w_156_712, w_156_713;
  wire w_157_016, w_157_038, w_157_105, w_157_180, w_157_528, w_157_539, w_157_557, w_157_739, w_157_754, w_157_814;
  wire w_158_009, w_158_069, w_158_076, w_158_079, w_158_082, w_158_145, w_158_198, w_158_213, w_158_225, w_158_356, w_158_392, w_158_546, w_158_633, w_158_643, w_158_841, w_158_847;
  wire w_159_004, w_159_062, w_159_064, w_159_074, w_159_102, w_159_149, w_159_169, w_159_192, w_159_221, w_159_227, w_159_245, w_159_253, w_159_260, w_159_264, w_159_285;
  wire w_160_072, w_160_073, w_160_081, w_160_088, w_160_155, w_160_181, w_160_320, w_160_359, w_160_431, w_160_599, w_160_638;
  wire w_161_081, w_161_104, w_161_124, w_161_221;
  wire w_162_051, w_162_133, w_162_139, w_162_146, w_162_154, w_162_173, w_162_181, w_162_210, w_162_244, w_162_249, w_162_298, w_162_321, w_162_326, w_162_359, w_162_396, w_162_427, w_162_466;
  wire w_163_002, w_163_047, w_163_068, w_163_095, w_163_120, w_163_176, w_163_181, w_163_215, w_163_235, w_163_237, w_163_341, w_163_536, w_163_642;
  wire w_164_035, w_164_037, w_164_042, w_164_069, w_164_109, w_164_129, w_164_131, w_164_155, w_164_183, w_164_186, w_164_193, w_164_314, w_164_326, w_164_375;
  wire w_165_098, w_165_120, w_165_140, w_165_187, w_165_203, w_165_277, w_165_362, w_165_550;
  wire w_166_015, w_166_020, w_166_041, w_166_047, w_166_120, w_166_219, w_166_269, w_166_294, w_166_327, w_166_331, w_166_360, w_166_531;
  wire w_167_031, w_167_042, w_167_069, w_167_234, w_167_265, w_167_275, w_167_280, w_167_290, w_167_406, w_167_416, w_167_458, w_167_495, w_167_557, w_167_656;
  wire w_168_104, w_168_128, w_168_133, w_168_361, w_168_387, w_168_412, w_168_541, w_168_767;
  wire w_169_017, w_169_021, w_169_022, w_169_034, w_169_036, w_169_042, w_169_050, w_169_068;
  wire w_170_032, w_170_045, w_170_166, w_170_171, w_170_199, w_170_220, w_170_275, w_170_289, w_170_407;
  wire w_171_042, w_171_188, w_171_189, w_171_215, w_171_242, w_171_264, w_171_280, w_171_296, w_171_326, w_171_333, w_171_359, w_171_369, w_171_391, w_171_472;
  wire w_172_030, w_172_060, w_172_109, w_172_299, w_172_315, w_172_357, w_172_365, w_172_388, w_172_405;
  wire w_173_043, w_173_069, w_173_110, w_173_120, w_173_158, w_173_432;
  wire w_174_149, w_174_189, w_174_269, w_174_453, w_174_516, w_174_538, w_174_762, w_174_857;
  wire w_175_182, w_175_456, w_175_551, w_175_828;
  wire w_176_067, w_176_154, w_176_180, w_176_201, w_176_270, w_176_361, w_176_380, w_176_479;
  wire w_177_030, w_177_072, w_177_095, w_177_278, w_177_347, w_177_395, w_177_524, w_177_549, w_177_639, w_177_701, w_177_790, w_177_863, w_177_912;
  wire w_178_014, w_178_016, w_178_351, w_178_504, w_178_590, w_178_600, w_178_883, w_178_943;
  wire w_179_022, w_179_218, w_179_549, w_179_713, w_179_724, w_179_888;
  wire w_180_005, w_180_050, w_180_075, w_180_160, w_180_172, w_180_210, w_180_269, w_180_305, w_180_333;
  wire w_181_103, w_181_162, w_181_211, w_181_234, w_181_388, w_181_495, w_181_516, w_181_790, w_181_802;
  wire w_182_038, w_182_039, w_182_073, w_182_091, w_182_115, w_182_120, w_182_122, w_182_159, w_182_188, w_182_193, w_182_210, w_182_223, w_182_227, w_182_228, w_182_274;
  wire w_183_035, w_183_041, w_183_053, w_183_067, w_183_070, w_183_110, w_183_224;
  wire w_184_008, w_184_039, w_184_049, w_184_085, w_184_157, w_184_173, w_184_191, w_184_243;
  wire w_185_031, w_185_061, w_185_078, w_185_100, w_185_103, w_185_118, w_185_149, w_185_202, w_185_277;
  wire w_186_001, w_186_007, w_186_042, w_186_070, w_186_198, w_186_304, w_186_442, w_186_479, w_186_544, w_186_609, w_186_618, w_186_642;
  wire w_187_011, w_187_022, w_187_024, w_187_096, w_187_099, w_187_131, w_187_148, w_187_153, w_187_161, w_187_175, w_187_183, w_187_203;
  wire w_188_073, w_188_087, w_188_123, w_188_161, w_188_427, w_188_430, w_188_491, w_188_535, w_188_536, w_188_537, w_188_538, w_188_539, w_188_543, w_188_544, w_188_545, w_188_546, w_188_547, w_188_548, w_188_550;
  wire w_189_071, w_189_115, w_189_117, w_189_298, w_189_346, w_189_525, w_189_974;
  wire w_190_000, w_190_068, w_190_168, w_190_222, w_190_237, w_190_261, w_190_289, w_190_348, w_190_394;
  wire w_191_036, w_191_037, w_191_083, w_191_118, w_191_135, w_191_142, w_191_174, w_191_211, w_191_278, w_191_294, w_191_316, w_191_325, w_191_385, w_191_392;
  wire w_192_000, w_192_001, w_192_002;
  wire w_193_003, w_193_042, w_193_197, w_193_252, w_193_290, w_193_291, w_193_314, w_193_340, w_193_416, w_193_418, w_193_454, w_193_669;
  wire w_194_011, w_194_077, w_194_089, w_194_211, w_194_219, w_194_268, w_194_283, w_194_433, w_194_453, w_194_471, w_194_495, w_194_593, w_194_699, w_194_909;
  wire w_195_029, w_195_070, w_195_082, w_195_181, w_195_256, w_195_335, w_195_348, w_195_487, w_195_517;
  wire w_196_045, w_196_274, w_196_306, w_196_453, w_196_712, w_196_728, w_196_808;
  wire w_197_140, w_197_143, w_197_189, w_197_237, w_197_352, w_197_422, w_197_541, w_197_674, w_197_746, w_197_778, w_197_838, w_197_896;
  wire w_198_040, w_198_074, w_198_220, w_198_315, w_198_322, w_198_330, w_198_578, w_198_741;
  wire w_199_044, w_199_056, w_199_060, w_199_131, w_199_419, w_199_751, w_199_795, w_199_829;
  wire w_200_029, w_200_166, w_200_262, w_200_683;
  wire w_201_076, w_201_095, w_201_276, w_201_514, w_201_655, w_201_698, w_201_719;
  wire w_202_003, w_202_009, w_202_011, w_202_012, w_202_015, w_202_018, w_202_019, w_202_020;
  wire w_203_061, w_203_082, w_203_098, w_203_110, w_203_156, w_203_258, w_203_304, w_203_312, w_203_407, w_203_512;
  wire w_204_218, w_204_257, w_204_342, w_204_363;
  wire w_205_113, w_205_126, w_205_427, w_205_566;
  wire w_206_057, w_206_126, w_206_334;
  wire w_207_005, w_207_023, w_207_104, w_207_147, w_207_226, w_207_236, w_207_244, w_207_353;
  wire w_208_026, w_208_028, w_208_032, w_208_267;
  wire w_209_171, w_209_179, w_209_180, w_209_203;
  wire w_210_314, w_210_523, w_210_574, w_210_681;
  wire w_211_029, w_211_040, w_211_050, w_211_052, w_211_133, w_211_150, w_211_241, w_211_276, w_211_498, w_211_528;
  wire w_212_013, w_212_084, w_212_102, w_212_109;
  wire w_213_041, w_213_433, w_213_538;
  wire w_214_005, w_214_027, w_214_039, w_214_052, w_214_070, w_214_075, w_214_092, w_214_100, w_214_107;
  wire w_215_092, w_215_170, w_215_267, w_215_322, w_215_422, w_215_428, w_215_565;
  wire w_216_050, w_216_102, w_216_126, w_216_129;
  wire w_217_209, w_217_279, w_217_372, w_217_797, w_217_819;
  wire w_218_004, w_218_016, w_218_141, w_218_204, w_218_428, w_218_582;
  wire w_219_030, w_219_038, w_219_064, w_219_069, w_219_146, w_219_217, w_219_277;
  wire w_220_034, w_220_055, w_220_257, w_220_604, w_220_608, w_220_821;
  wire w_221_070, w_221_136, w_221_396, w_221_550;
  wire w_222_045, w_222_259, w_222_477, w_222_662;
  wire w_223_023, w_223_141, w_223_157, w_223_278, w_223_379, w_223_493, w_223_582, w_223_631, w_223_840, w_223_925;
  wire w_224_009, w_224_038, w_224_041, w_224_042, w_224_052, w_224_058, w_224_075;
  wire w_225_002, w_225_022, w_225_026;
  wire w_226_000, w_226_001, w_226_005, w_226_008, w_226_010, w_226_013;
  wire w_227_012, w_227_067, w_227_199, w_227_260, w_227_408, w_227_416, w_227_522, w_227_547;
  wire w_228_267, w_228_288, w_228_329, w_228_637, w_228_745;
  wire w_229_076, w_229_125, w_229_274, w_229_295;
  wire w_230_032, w_230_036, w_230_048, w_230_082, w_230_238, w_230_246, w_230_248, w_230_251, w_230_252, w_230_262, w_230_295;
  wire w_231_002, w_231_026, w_231_036, w_231_049, w_231_057, w_231_083;
  wire w_232_008, w_232_029, w_232_032, w_232_146, w_232_202, w_232_235, w_232_363;
  wire w_233_078, w_233_128, w_233_319, w_233_342, w_233_384, w_233_391;
  wire w_234_050, w_234_515, w_234_554;
  wire w_235_019, w_235_058, w_235_140;
  wire w_236_047, w_236_050, w_236_151, w_236_154, w_236_162, w_236_300, w_236_315, w_236_410, w_236_606;
  wire w_237_228, w_237_276, w_237_376, w_237_379, w_237_423;
  wire w_238_033, w_238_053, w_238_080, w_238_159, w_238_218, w_238_231, w_238_251, w_238_285, w_238_312, w_238_350, w_238_360, w_238_389;
  wire w_239_054, w_239_174, w_239_183, w_239_648, w_239_678, w_239_728;
  wire w_240_011, w_240_178, w_240_754, w_240_814, w_240_815, w_240_816, w_240_817, w_240_818, w_240_819, w_240_820, w_240_821;
  wire w_241_027, w_241_065, w_241_142, w_241_276, w_241_336, w_241_344;
  wire w_242_106, w_242_173, w_242_223;
  wire w_243_003, w_243_013, w_243_075, w_243_109, w_243_141, w_243_147, w_243_152, w_243_205, w_243_223;
  wire w_244_160, w_244_220;
  wire w_245_076, w_245_090, w_245_236, w_245_277, w_245_297;
  wire w_246_002, w_246_107, w_246_253, w_246_274, w_246_276, w_246_287;
  wire w_247_091, w_247_092, w_247_496, w_247_498, w_247_610, w_247_611;
  wire w_248_014, w_248_299, w_248_327, w_248_459, w_248_648;
  wire w_249_036, w_249_065, w_249_193, w_249_223, w_249_255;
  wire w_250_003, w_250_055, w_250_059, w_250_068, w_250_226, w_250_287, w_250_420, w_250_445;
  wire w_251_026, w_251_031, w_251_208, w_251_229, w_251_259, w_251_262;
  wire w_252_190, w_252_225, w_252_358, w_252_383;
  wire w_253_000, w_253_003, w_253_005, w_253_009, w_253_031, w_253_032, w_253_048;
  wire w_254_057, w_254_184, w_254_269, w_254_306;
  wire w_255_000, w_255_003, w_255_007, w_255_033, w_255_036;
  wire w_256_020, w_256_047, w_256_124;
  wire w_257_044, w_257_146, w_257_271, w_257_402, w_257_428, w_257_512, w_257_562;
  wire w_258_122, w_258_236, w_258_754;
  wire w_259_099, w_259_167, w_259_234, w_259_308, w_259_372, w_259_461, w_259_505;
  wire w_260_123, w_260_154, w_260_373, w_260_510, w_260_578, w_260_616, w_260_751, w_260_812;
  wire w_261_418, w_261_469;
  wire w_262_035, w_262_059, w_262_086, w_262_110, w_262_146;
  wire w_263_069, w_263_077, w_263_093, w_263_174, w_263_189, w_263_199;
  wire w_264_132, w_264_371, w_264_439, w_264_606, w_264_782, w_264_796, w_264_900;
  wire w_265_059, w_265_060, w_265_065, w_265_068, w_265_075, w_265_202, w_265_414, w_265_528;
  wire w_266_295, w_266_429, w_266_451;
  wire w_267_076, w_267_088, w_267_111, w_267_141, w_267_225, w_267_550, w_267_602;
  wire w_268_116, w_268_172, w_268_353, w_268_446;
  wire w_269_017, w_269_031, w_269_035;
  wire w_270_103, w_270_166, w_270_174, w_270_473, w_270_681;
  wire w_271_002, w_271_038, w_271_039, w_271_074, w_271_107, w_271_157;
  wire w_272_135;
  wire w_273_061, w_273_127, w_273_366;
  wire w_274_000, w_274_002;
  wire w_275_000, w_275_002, w_275_003;
  wire w_276_645, w_276_686;
  wire w_277_033, w_277_088, w_277_106, w_277_109;
  wire w_278_065, w_278_216, w_278_224, w_278_359, w_278_442;
  wire w_279_032, w_279_088, w_279_344;
  wire w_280_002, w_280_016, w_280_018, w_280_019, w_280_023;
  wire w_281_029, w_281_115, w_281_197, w_281_344, w_281_706;
  wire w_282_074, w_282_103;
  wire w_283_079, w_283_250, w_283_283, w_283_335, w_283_355, w_283_373, w_283_498;
  wire w_284_079, w_284_092, w_284_102, w_284_229, w_284_312, w_284_405, w_284_430, w_284_462;
  wire w_285_102, w_285_158;
  wire w_286_249;
  wire w_287_109, w_287_110, w_287_395, w_287_695;
  wire w_288_135, w_288_203, w_288_353, w_288_665;
  wire w_289_304, w_289_480, w_289_855;
  wire w_290_052, w_290_115, w_290_183, w_290_260;
  wire w_291_035, w_291_052, w_291_707;
  wire w_292_109, w_292_160, w_292_235, w_292_413, w_292_705, w_292_706, w_292_707, w_292_708, w_292_709, w_292_710, w_292_711, w_292_712, w_292_713, w_292_714;
  wire w_293_051, w_293_087, w_293_573, w_293_625, w_293_697;
  wire w_294_010, w_294_038, w_294_279, w_294_644, w_294_710;
  wire w_295_009, w_295_080, w_295_116, w_295_170;
  wire w_296_000, w_296_017, w_296_067;
  wire w_297_114, w_297_117, w_297_138, w_297_150, w_297_196;
  wire w_298_205;
  wire w_299_079, w_299_134;
  wire w_300_036, w_300_208, w_300_507, w_300_631, w_300_854;
  wire w_301_070, w_301_356, w_301_478;
  wire w_302_000, w_302_016, w_302_020, w_302_023, w_302_029;
  wire w_304_041, w_304_046, w_304_064, w_304_079;
  wire w_305_009, w_305_046, w_305_083, w_305_091, w_305_093, w_305_097, w_305_151;
  wire w_306_015, w_306_018, w_306_028, w_306_072, w_306_088, w_306_091, w_306_137;
  wire w_307_312;
  wire w_308_061, w_308_084;
  wire w_309_002, w_309_115, w_309_151, w_309_164, w_309_193;
  wire w_310_259;
  wire w_311_140, w_311_169;
  wire w_312_051, w_312_791, w_312_894;
  wire w_313_027, w_313_166, w_313_170, w_313_228, w_313_246, w_313_446, w_313_477;
  wire w_314_086, w_314_388, w_314_765;
  wire w_315_105, w_315_129, w_315_455, w_315_491;
  wire w_316_056, w_316_137, w_316_320, w_316_635, w_316_731, w_316_852, w_316_853, w_316_854, w_316_855, w_316_856, w_316_857, w_316_858, w_316_859, w_316_860, w_316_861, w_316_862;
  wire w_317_043, w_317_059, w_317_533, w_317_562, w_317_740;
  wire w_318_024, w_318_026, w_318_031, w_318_038, w_318_051, w_318_063, w_318_064, w_318_065, w_318_066, w_318_067, w_318_068, w_318_069, w_318_070, w_318_071, w_318_072;
  wire w_319_072, w_319_254;
  wire w_320_029, w_320_101, w_320_365, w_320_609;
  wire w_321_011, w_321_277, w_321_543, w_321_763;
  wire w_322_585;
  wire w_323_219, w_323_372, w_323_678, w_323_902;
  wire w_324_020, w_324_030, w_324_151, w_324_589;
  wire w_325_027, w_325_156, w_325_265;
  wire w_326_011, w_326_193;
  wire w_327_007, w_327_025, w_327_728, w_327_873;
  wire w_328_273;
  wire w_329_037, w_329_379, w_329_502;
  wire w_330_072, w_330_107, w_330_151;
  wire w_331_007, w_331_050, w_331_087, w_331_095;
  wire w_332_075, w_332_147, w_332_161, w_332_184, w_332_407;
  wire w_333_108, w_333_374, w_333_540;
  wire w_334_000, w_334_002;
  wire w_335_094, w_335_105;
  wire w_336_047, w_336_056;
  wire w_338_448, w_338_783;
  wire w_339_117;
  wire w_340_120, w_340_224, w_340_315, w_340_328;
  wire w_341_018, w_341_025, w_341_044, w_341_045, w_341_046;
  wire w_342_109, w_342_140, w_342_172, w_342_504;
  wire w_343_076, w_343_160, w_343_172;
  wire w_344_000, w_344_001;
  wire w_345_197;
  wire w_346_012, w_346_022, w_346_024, w_346_038;
  wire w_347_123, w_347_130;
  wire w_348_000;
  wire w_349_067, w_349_088;
  wire w_350_011, w_350_226;
  wire w_351_002, w_351_004, w_351_041, w_351_044, w_351_045;
  wire w_352_075, w_352_100;
  wire w_353_055, w_353_057, w_353_080, w_353_088, w_353_102;
  wire w_354_345, w_354_649;
  wire w_355_160;
  wire w_356_012, w_356_475, w_356_701, w_356_756;
  wire w_357_147;
  wire w_358_031, w_358_421, w_358_438, w_358_607, w_358_750;
  wire w_359_460;
  wire w_360_035;
  wire w_361_000, w_361_026, w_361_029, w_361_032, w_361_059;
  wire w_362_019, w_362_069, w_362_083;
  wire w_363_006;
  wire w_364_383, w_364_803;
  wire w_365_043, w_365_069, w_365_145;
  wire w_366_160, w_366_444;
  wire w_367_053, w_367_133, w_367_180, w_367_243;
  wire w_368_005, w_368_006;
  wire w_369_005, w_369_081, w_369_305;
  wire w_370_154;
  wire w_371_053;
  wire w_372_378, w_372_442, w_372_455;
  wire w_373_024, w_373_069;
  wire w_374_011, w_374_012;
  wire w_375_045;
  wire w_376_277, w_376_391;
  wire w_377_168, w_377_284, w_377_395, w_377_418;
  wire w_378_247;
  wire w_379_001, w_379_050, w_379_060;
  wire w_380_030, w_380_104, w_380_107, w_380_238;
  wire w_381_222, w_381_632;
  wire w_382_232, w_382_405, w_382_610;
  wire w_383_005, w_383_095, w_383_156, w_383_337, w_383_420;
  wire w_385_375;
  wire w_386_036, w_386_195, w_386_630;
  wire w_387_049;
  wire w_388_023, w_388_079, w_388_098, w_388_100, w_388_223, w_388_244;
  wire w_389_061, w_389_068, w_389_092, w_389_335;
  wire w_390_033;
  wire w_391_028;
  wire w_392_000;
  wire w_393_163, w_393_323;
  wire w_394_103, w_394_118, w_394_129, w_394_195;
  wire w_395_026, w_395_081, w_395_103, w_395_161;
  wire w_396_533;
  wire w_397_098, w_397_194, w_397_197, w_397_322;
  wire w_398_362;
  wire w_399_008, w_399_050, w_399_061, w_399_064, w_399_091;
  wire w_400_025, w_400_203, w_400_790, w_400_791, w_400_792, w_400_793, w_400_794, w_400_795, w_400_796, w_400_797, w_400_798;
  wire w_401_500, w_401_636, w_401_729, w_401_785;
  wire w_402_188, w_402_217;
  wire w_403_085, w_403_140, w_403_276, w_403_277, w_403_278;
  wire w_404_022, w_404_049;
  wire w_405_131, w_405_146, w_405_393, w_405_439, w_405_808;
  wire w_406_013, w_406_047, w_406_263, w_406_437, w_406_577;
  wire w_407_039, w_407_066;
  wire w_408_011, w_408_090;
  wire w_410_001, w_410_093;
  wire w_411_948;
  wire w_412_106, w_412_147, w_412_746;
  wire w_413_287, w_413_446;
  wire w_414_008, w_414_153, w_414_162;
  wire w_415_059, w_415_247, w_415_370;
  wire w_416_134, w_416_301, w_416_719, w_416_776, w_416_777, w_416_778, w_416_779, w_416_780, w_416_781;
  wire w_417_005, w_417_149, w_417_156;
  wire w_418_005, w_418_034;
  wire w_420_527;
  wire w_421_003, w_421_146, w_421_159;
  wire w_422_026, w_422_041;
  wire w_423_027, w_423_151, w_423_235;
  wire w_424_038, w_424_083, w_424_336, w_424_509;
  wire w_427_082, w_427_096, w_427_358;
  wire w_428_557, w_428_765;
  wire w_429_111, w_429_135, w_429_153, w_429_244;
  wire w_430_279;
  wire w_431_019, w_431_024, w_431_025;
  wire w_432_022, w_432_026;
  wire w_433_066, w_433_391;
  wire w_435_077, w_435_087, w_435_090;
  wire w_436_087, w_436_096, w_436_111;
  wire w_437_005, w_437_050, w_437_069;
  wire w_438_352;
  wire w_439_237;
  wire w_440_157, w_440_458, w_440_479, w_440_495;
  wire w_441_004, w_441_011, w_441_013;
  wire w_442_003, w_442_014, w_442_020, w_442_053, w_442_089;
  wire w_444_000, w_444_005, w_444_007;
  wire w_445_010, w_445_017, w_445_024, w_445_037;
  wire w_446_650;
  wire w_447_210, w_447_349, w_447_499;
  wire w_449_078, w_449_110;
  wire w_450_081, w_450_116, w_450_117, w_450_118, w_450_119, w_450_120, w_450_121, w_450_122, w_450_123;
  wire w_451_379;
  wire w_452_044, w_452_487;
  wire w_453_179;
  wire w_454_165, w_454_685;
  wire w_455_040, w_455_105, w_455_112;
  wire w_457_023, w_457_071, w_457_092;
  wire w_459_131;
  wire w_460_255, w_460_536;
  wire w_461_112, w_461_186;
  wire w_462_369;
  wire w_464_156;
  wire w_465_326, w_465_523;
  wire w_466_177, w_466_287;
  wire w_467_016, w_467_042;
  wire w_468_004, w_468_052, w_468_080;
  wire w_469_058, w_469_209, w_469_565;
  wire w_470_021;
  wire w_471_332, w_471_893;
  wire w_474_405, w_474_430, w_474_431, w_474_432, w_474_433, w_474_434, w_474_438, w_474_439, w_474_440, w_474_441, w_474_442, w_474_443, w_474_444, w_474_445, w_474_446, w_474_447, w_474_449;
  wire w_476_110, w_476_174, w_476_782;
  wire w_477_060, w_477_460, w_477_648, w_477_713;
  wire w_478_050;
  wire w_479_086, w_479_183, w_479_188;
  wire w_480_046, w_480_285;
  wire w_482_031;
  wire w_483_180, w_483_216, w_483_217, w_483_218, w_483_219, w_483_220, w_483_221, w_483_222, w_483_223, w_483_224, w_483_225, w_483_226, w_483_227;
  wire w_484_159, w_484_422, w_484_522, w_484_601;
  wire w_486_233;
  wire w_487_023, w_487_195, w_487_231;
  wire w_488_004, w_488_061, w_488_066, w_488_117;
  wire w_489_029;
  wire w_490_392;
  wire w_491_184, w_491_222, w_491_453;
  wire w_493_023;
  wire w_494_418, w_494_428;
  wire w_495_061;
  wire w_497_072, w_497_367;
  wire w_498_003, w_498_527;
  wire w_499_113, w_499_268, w_499_278;
  wire w_500_173;
  wire w_501_029, w_501_049;
  wire w_502_002, w_502_014;
  wire w_503_031, w_503_730, w_503_731, w_503_732, w_503_733, w_503_734, w_503_735, w_503_736, w_503_737, w_503_738, w_503_739, w_503_743, w_503_744, w_503_745, w_503_746, w_503_747, w_503_748, w_503_749, w_503_750, w_503_751, w_503_752, w_503_754;
  wire w_504_203;
  wire w_505_085, w_505_686;
  wire w_508_000;
  wire w_509_022, w_509_040;
  wire w_510_377, w_510_748;
  wire w_511_108, w_511_753;
  wire w_512_001, w_512_120, w_512_345;
  wire w_513_218;
  wire w_514_204;
  wire w_515_129, w_515_169, w_515_535;
  wire w_517_397;
  wire w_518_369, w_518_760;
  wire w_519_060, w_519_098;
  wire w_520_251, w_520_860;
  wire w_521_000;
  wire w_524_068, w_524_639;
  wire w_525_019, w_525_027;
  wire w_526_150;
  wire w_527_041, w_527_056, w_527_095, w_527_113;
  wire w_528_000, w_528_087;
  wire w_529_240, w_529_542, w_529_947;
  wire w_530_171, w_530_524;
  wire w_531_104, w_531_273, w_531_352;
  wire w_534_277;
  wire w_536_295;
  wire w_537_074;
  wire w_538_778;
  wire w_539_036, w_539_064;
  wire w_541_008, w_541_013, w_541_068;
  wire w_543_064;
  wire w_545_264, w_545_270;
  wire w_546_205;
  wire w_547_131, w_547_377, w_547_427;
  wire w_550_001, w_550_051;
  wire w_551_922;
  wire w_552_506, w_552_556;
  wire w_553_655;
  wire w_555_112;
  wire w_556_244;
  wire w_558_351;
  wire w_559_126, w_559_352;
  wire w_560_550, w_560_731;
  wire w_561_112;
  wire w_562_064;
  wire w_563_002, w_563_007, w_563_029;
  wire w_564_518, w_564_612;
  wire w_565_169, w_565_447, w_565_579, w_565_627, w_565_653;
  wire w_566_252, w_566_464;
  wire w_567_204, w_567_775;
  wire w_568_144;
  wire w_569_371;
  wire w_570_277;
  wire w_571_125;
  wire w_572_339, w_572_469;
  wire w_573_015;
  wire w_576_060, w_576_076;
  wire w_577_770;
  wire w_578_013, w_578_116, w_578_266;
  wire w_580_001, w_580_034;
  wire w_581_048, w_581_068, w_581_206;
  wire w_582_163;
  wire w_584_143, w_584_242;
  wire w_585_305;
  wire w_586_005;
  wire w_588_655, w_588_660, w_588_885;
  wire w_589_435, w_589_696;
  wire w_590_483;
  wire w_592_237;
  wire w_593_338, w_593_555;
  wire w_594_047, w_594_071, w_594_088;
  wire w_595_052, w_595_289;
  wire w_597_010, w_597_154, w_597_305, w_597_329, w_597_330, w_597_331, w_597_332, w_597_333, w_597_334, w_597_335, w_597_336, w_597_337, w_597_341, w_597_342, w_597_343, w_597_344, w_597_345, w_597_346, w_597_347, w_597_348, w_597_349, w_597_351;
  wire w_600_055;
  wire w_601_099;
  wire w_604_292, w_604_585, w_604_740;
  wire w_606_125, w_606_297, w_606_398;
  wire w_610_161, w_610_178;
  wire w_611_013;
  wire w_612_023;
  wire w_613_169, w_613_372;
  wire w_614_603;
  wire w_615_006;
  wire w_617_055;
  wire w_618_328;
  wire w_619_158;
  wire w_620_386, w_620_448;
  wire w_622_073;
  wire w_623_290;
  wire w_624_007, w_624_026;
  wire w_625_023;
  wire w_626_001;
  wire w_628_163;
  wire w_630_006, w_630_101;
  wire w_633_074, w_633_156;
  wire w_635_153;
  wire w_637_226, w_637_537;
  wire w_638_381;
  wire w_639_173;
  wire w_643_784, w_643_889;
  wire w_644_029, w_644_288, w_644_363, w_644_394;
  wire w_646_006, w_646_027;
  wire w_651_087;
  wire w_652_169, w_652_187;
  wire w_654_033;
  wire w_656_184;
  wire w_657_576;
  wire w_658_148;
  wire w_665_155;
  wire w_667_474;
  wire w_671_004, w_671_349;
  wire w_673_893;
  wire w_675_073;
  wire w_677_133;
  wire w_679_446;
  wire w_681_125;
  wire w_684_004, w_684_012, w_684_680;
  wire w_685_052, w_685_145;
  wire w_686_000, w_686_047;
  wire w_687_067, w_687_271;
  wire w_689_222, w_689_272, w_689_291;
  wire w_690_226, w_690_459;
  wire w_691_066;
  wire w_692_415;
  wire w_693_100;
  wire w_694_016;
  wire w_698_419;
  wire w_700_169;
  wire w_701_285, w_701_509;
  wire w_702_177;
  wire w_703_212, w_703_395, w_703_396, w_703_397, w_703_398, w_703_399, w_703_400, w_703_401, w_703_402, w_703_403, w_703_404, w_703_405, w_703_406;
  wire w_705_598;
  wire w_706_150, w_706_155;
  wire w_707_071, w_707_146;
  wire w_713_009, w_713_133, w_713_134, w_713_135, w_713_139, w_713_140, w_713_141, w_713_142, w_713_143, w_713_144, w_713_145, w_713_146, w_713_147, w_713_148, w_713_149, w_713_151;
  wire w_716_133;
  wire w_718_257;
  wire w_719_615, w_719_616, w_719_617, w_719_618, w_719_619, w_719_620, w_719_621, w_719_622, w_719_623;
  wire w_720_811, w_720_812, w_720_813, w_720_814, w_720_815, w_720_816;
  wire w_721_179, w_721_271;
  wire w_722_521;
  wire w_723_185;
  wire w_729_129;
  wire w_730_090;
  wire w_731_104;
  wire w_732_078;
  wire w_737_368, w_737_555, w_737_556, w_737_557, w_737_558, w_737_559, w_737_560, w_737_561;
  wire w_739_365;
  wire w_740_340;
  wire w_742_037, w_742_744;
  wire w_743_142, w_743_143, w_743_144, w_743_145, w_743_146;
  wire w_745_143;
  wire w_746_004;
  wire w_749_165;
  wire w_751_361;
  wire w_753_047;
  wire w_754_035, w_754_554;
  wire w_755_022;
  wire w_756_019;
  wire w_757_254;
  wire w_759_380;
  wire w_761_008;
  wire w_762_761;
  wire w_764_052, w_764_518;
  wire w_768_177;
  wire w_771_065;
  wire w_775_531, w_775_618;
  wire w_777_041;
  wire w_778_142, w_778_263;
  wire w_780_073;
  wire w_783_313;
  wire w_784_017;
  wire w_787_430;
  wire w_788_201, w_788_202, w_788_203, w_788_204, w_788_205, w_788_209, w_788_210, w_788_211, w_788_212, w_788_213, w_788_214, w_788_215, w_788_216, w_788_217, w_788_219;
  wire w_789_570;
  wire w_790_729;
  wire w_791_166;
  wire w_795_038, w_795_155;
  wire w_796_256;
  wire w_797_385;
  wire w_802_628, w_802_629, w_802_630, w_802_631, w_802_632, w_802_633, w_802_634;
  wire w_804_005;
  wire w_805_240;
  wire w_807_002;
  wire w_809_082;
  wire w_813_317;
  wire w_820_016;
  wire w_821_033;
  wire w_822_988, w_822_989, w_822_990;
  wire w_826_020, w_826_130;
  wire w_828_076, w_828_088;
  wire w_829_086, w_829_467;
  wire w_832_482;
  wire w_838_328;
  wire w_842_229;
  wire w_843_544;
  wire w_844_288;
  wire w_845_074;
  wire w_846_004;
  wire w_847_002, w_847_003, w_847_004, w_847_005, w_847_006;
  wire w_848_326, w_848_335;
  wire w_850_023;
  wire w_853_747;
  wire w_856_011;
  wire w_860_088, w_860_491;
  wire w_863_324;
  wire w_866_111;
  wire w_869_114;
  wire w_871_145, w_871_351;
  wire w_873_255;
  wire w_875_165, w_875_251;
  wire w_876_001;
  wire w_878_548, w_878_681, w_878_748, w_878_749, w_878_750, w_878_751, w_878_752, w_878_753, w_878_754, w_878_755, w_878_759, w_878_760, w_878_761, w_878_762, w_878_763, w_878_764, w_878_766;
  wire w_881_105;
  wire w_882_423;
  wire w_883_420;
  wire w_887_066;
  wire w_888_266;
  wire w_889_143, w_889_239, w_889_352;
  wire w_891_119, w_891_163;
  wire w_893_103, w_893_145;
  wire w_894_262, w_894_263, w_894_264, w_894_265, w_894_266, w_894_267, w_894_268, w_894_269, w_894_270, w_894_271, w_894_272, w_894_273, w_894_277, w_894_278, w_894_279, w_894_280, w_894_281, w_894_282, w_894_283, w_894_284, w_894_285, w_894_287;
  wire w_896_755, w_896_756, w_896_757, w_896_758;
  wire w_899_531, w_899_532, w_899_533, w_899_534, w_899_535, w_899_536, w_899_537, w_899_538, w_899_539, w_899_540;
  wire w_901_380;
  wire w_904_126;
  wire w_905_810, w_905_811, w_905_812, w_905_816, w_905_817, w_905_818, w_905_819, w_905_820, w_905_821, w_905_823;
  wire w_907_282;
  wire w_908_298;
  wire w_914_427;
  wire w_916_185, w_916_358;
  wire w_919_108, w_919_354;
  wire w_921_163;
  wire w_924_279, w_924_298;
  wire w_927_320;
  wire w_928_157;
  wire w_930_000;
  wire w_931_517;
  wire w_933_375;
  wire w_935_942, w_935_969, w_935_970, w_935_971, w_935_972, w_935_973, w_935_977, w_935_978, w_935_979, w_935_981;
  wire w_938_341;
  wire w_942_549;
  wire w_943_456;
  wire w_945_256;
  wire w_949_032;
  wire w_952_565, w_952_772;
  wire w_954_012;
  wire w_955_092, w_955_348, w_955_349, w_955_350, w_955_351, w_955_352, w_955_353, w_955_354, w_955_355, w_955_356, w_955_357;
  wire w_966_010, w_966_534;
  wire w_967_137;
  wire w_968_916, w_968_917, w_968_918, w_968_919, w_968_920, w_968_921, w_968_922, w_968_923, w_968_924, w_968_925, w_968_926, w_968_927, w_968_931, w_968_932, w_968_933, w_968_934, w_968_936;
  wire w_971_280, w_971_281, w_971_282, w_971_283, w_971_284, w_971_285, w_971_286, w_971_287, w_971_288;
  wire w_973_121;
  wire w_974_075;
  wire w_975_059;
  wire w_977_099;
  wire w_978_339;
  wire w_980_815;
  wire w_982_324;
  wire w_986_106, w_986_714;
  wire w_991_282;
  wire w_996_052;
  wire w_1000_000, w_1000_001, w_1000_002, w_1000_003, w_1000_004, w_1000_005, w_1000_006, w_1000_007, w_1000_008, w_1000_009, w_1000_010, w_1000_011, w_1000_012, w_1000_013, w_1000_014, w_1000_015, w_1000_016, w_1000_017, w_1000_018, w_1000_019, w_1000_020, w_1000_021, w_1000_022, w_1000_023, w_1000_024, w_1000_025, w_1000_026, w_1000_027, w_1000_028, w_1000_029, w_1000_030, w_1000_031, w_1000_032, w_1000_033, w_1000_034, w_1000_035, w_1000_036, w_1000_037, w_1000_038, w_1000_039, w_1000_040, w_1000_041, w_1000_042, w_1000_043, w_1000_044, w_1000_045, w_1000_046, w_1000_047, w_1000_048, w_1000_049, w_1000_050, w_1000_051, w_1000_052, w_1000_053, w_1000_054, w_1000_055, w_1000_056, w_1000_057, w_1000_058, w_1000_059, w_1000_060, w_1000_061, w_1000_062, w_1000_063, w_1000_064, w_1000_065, w_1000_066, w_1000_067, w_1000_068, w_1000_069, w_1000_070, w_1000_071, w_1000_072, w_1000_073, w_1000_074, w_1000_075, w_1000_076, w_1000_077, w_1000_078, w_1000_079, w_1000_080, w_1000_081, w_1000_082, w_1000_083, w_1000_084, w_1000_085, w_1000_086, w_1000_087, w_1000_088, w_1000_089, w_1000_090, w_1000_091, w_1000_092, w_1000_093, w_1000_094, w_1000_095, w_1000_096, w_1000_097, w_1000_098, w_1000_099, w_1000_100, w_1000_101, w_1000_102, w_1000_103, w_1000_104, w_1000_105, w_1000_106, w_1000_107, w_1000_108, w_1000_109, w_1000_110, w_1000_111, w_1000_112, w_1000_113, w_1000_114, w_1000_115, w_1000_116, w_1000_117, w_1000_118, w_1000_119, w_1000_120, w_1000_121, w_1000_122, w_1000_123, w_1000_124, w_1000_125, w_1000_126, w_1000_127, w_1000_128, w_1000_129, w_1000_130, w_1000_131, w_1000_132, w_1000_133, w_1000_134, w_1000_135, w_1000_136, w_1000_137, w_1000_138, w_1000_139, w_1000_140, w_1000_141, w_1000_142, w_1000_143, w_1000_144, w_1000_145, w_1000_146, w_1000_147, w_1000_148, w_1000_149, w_1000_150, w_1000_151, w_1000_152, w_1000_153, w_1000_154, w_1000_155, w_1000_156, w_1000_157, w_1000_158, w_1000_159, w_1000_160, w_1000_161, w_1000_162, w_1000_163, w_1000_164, w_1000_165, w_1000_166, w_1000_167, w_1000_168, w_1000_169, w_1000_170, w_1000_171, w_1000_172, w_1000_173, w_1000_174, w_1000_175, w_1000_176, w_1000_177, w_1000_178, w_1000_179, w_1000_180, w_1000_181, w_1000_182, w_1000_183, w_1000_184, w_1000_185;
  not1 I001_000(w_001_000, w_000_000);
  nand2 I001_001(w_001_001, w_000_001, w_000_002);
  not1 I001_002(w_001_002, w_000_003);
  or2  I001_003(w_001_003, w_000_004, w_000_005);
  nand2 I001_004(w_001_004, w_000_006, w_000_007);
  nand2 I001_005(w_001_005, w_000_008, w_000_009);
  not1 I001_006(w_001_006, w_000_010);
  and2 I001_007(w_001_007, w_000_011, w_000_012);
  nand2 I001_008(w_001_008, w_000_013, w_000_014);
  not1 I001_009(w_001_009, w_000_015);
  nand2 I001_010(w_001_010, w_000_016, w_000_017);
  or2  I001_011(w_001_011, w_000_018, w_000_019);
  not1 I001_012(w_001_012, w_000_020);
  nand2 I001_013(w_001_013, w_000_021, w_000_022);
  nand2 I001_014(w_001_014, w_000_023, w_000_024);
  or2  I001_015(w_001_015, w_000_025, w_000_026);
  and2 I001_016(w_001_016, w_000_027, w_000_028);
  and2 I001_017(w_001_017, w_000_029, w_000_030);
  or2  I001_018(w_001_018, w_000_031, w_000_032);
  and2 I001_019(w_001_019, w_000_033, w_000_034);
  not1 I001_020(w_001_020, w_000_035);
  and2 I001_021(w_001_021, w_000_036, w_000_037);
  or2  I001_022(w_001_022, w_000_038, w_000_039);
  and2 I001_023(w_001_023, w_000_040, w_000_041);
  or2  I001_024(w_001_024, w_000_042, w_000_043);
  or2  I001_026(w_001_026, w_000_046, w_000_047);
  not1 I001_027(w_001_027, w_000_048);
  nand2 I001_028(w_001_028, w_000_049, w_000_050);
  and2 I001_029(w_001_029, w_000_051, w_000_052);
  and2 I001_030(w_001_030, w_000_053, w_000_054);
  nand2 I001_031(w_001_031, w_000_055, w_000_056);
  and2 I001_032(w_001_032, w_000_057, w_000_058);
  and2 I001_033(w_001_033, w_000_059, w_000_012);
  not1 I001_034(w_001_034, w_000_060);
  not1 I001_035(w_001_035, w_000_061);
  nand2 I001_036(w_001_036, w_000_062, w_000_063);
  not1 I001_037(w_001_037, w_000_064);
  or2  I001_038(w_001_038, w_000_065, w_000_066);
  or2  I001_039(w_001_039, w_000_067, w_000_068);
  and2 I001_040(w_001_040, w_000_069, w_000_070);
  not1 I001_041(w_001_041, w_000_071);
  or2  I001_042(w_001_042, w_000_072, w_000_073);
  nand2 I001_043(w_001_043, w_000_074, w_000_075);
  nand2 I001_044(w_001_044, w_000_076, w_000_077);
  or2  I001_046(w_001_046, w_000_080, w_000_081);
  and2 I001_047(w_001_047, w_000_082, w_000_083);
  not1 I001_048(w_001_048, w_000_084);
  nand2 I001_050(w_001_050, w_000_086, w_000_087);
  nand2 I001_051(w_001_051, w_000_088, w_000_089);
  nand2 I001_052(w_001_052, w_000_019, w_000_090);
  and2 I001_053(w_001_053, w_000_091, w_000_092);
  and2 I001_054(w_001_054, w_000_093, w_000_094);
  nand2 I001_055(w_001_055, w_000_095, w_000_096);
  not1 I001_056(w_001_056, w_000_097);
  or2  I001_057(w_001_057, w_000_098, w_000_099);
  and2 I001_058(w_001_058, w_000_100, w_000_101);
  or2  I001_059(w_001_059, w_000_102, w_000_103);
  and2 I001_060(w_001_060, w_000_034, w_000_104);
  and2 I001_061(w_001_061, w_000_105, w_000_106);
  and2 I001_062(w_001_062, w_000_107, w_000_108);
  nand2 I001_063(w_001_063, w_000_109, w_000_110);
  and2 I001_064(w_001_064, w_000_111, w_000_112);
  or2  I001_065(w_001_065, w_000_113, w_000_114);
  nand2 I001_066(w_001_066, w_000_115, w_000_116);
  or2  I001_068(w_001_068, w_000_118, w_000_119);
  or2  I001_069(w_001_069, w_000_120, w_000_121);
  nand2 I001_070(w_001_070, w_000_011, w_000_122);
  or2  I001_071(w_001_071, w_000_123, w_000_124);
  nand2 I001_072(w_001_072, w_000_125, w_000_126);
  not1 I001_073(w_001_073, w_000_127);
  and2 I001_074(w_001_074, w_000_128, w_000_129);
  and2 I001_075(w_001_075, w_000_130, w_000_131);
  or2  I001_076(w_001_076, w_000_132, w_000_133);
  and2 I001_077(w_001_077, w_000_134, w_000_135);
  nand2 I001_078(w_001_078, w_000_136, w_000_137);
  and2 I001_079(w_001_079, w_000_138, w_000_139);
  not1 I001_080(w_001_080, w_000_140);
  nand2 I001_081(w_001_081, w_000_141, w_000_142);
  or2  I001_082(w_001_082, w_000_082, w_000_143);
  and2 I001_083(w_001_083, w_000_144, w_000_145);
  nand2 I001_084(w_001_084, w_000_146, w_000_147);
  nand2 I001_085(w_001_085, w_000_148, w_000_149);
  nand2 I001_086(w_001_086, w_000_150, w_000_151);
  and2 I001_087(w_001_087, w_000_152, w_000_153);
  nand2 I001_088(w_001_088, w_000_154, w_000_155);
  or2  I001_089(w_001_089, w_000_156, w_000_157);
  not1 I001_090(w_001_090, w_000_158);
  and2 I001_091(w_001_091, w_000_159, w_000_160);
  not1 I001_092(w_001_092, w_000_161);
  or2  I001_093(w_001_093, w_000_162, w_000_163);
  not1 I001_094(w_001_094, w_000_164);
  and2 I001_095(w_001_095, w_000_165, w_000_062);
  and2 I001_096(w_001_096, w_000_166, w_000_036);
  and2 I001_097(w_001_097, w_000_167, w_000_168);
  not1 I001_098(w_001_098, w_000_169);
  nand2 I001_099(w_001_099, w_000_170, w_000_131);
  or2  I001_100(w_001_100, w_000_171, w_000_172);
  not1 I001_101(w_001_101, w_000_173);
  nand2 I001_102(w_001_102, w_000_174, w_000_175);
  nand2 I001_103(w_001_103, w_000_176, w_000_177);
  or2  I001_104(w_001_104, w_000_178, w_000_179);
  and2 I001_107(w_001_107, w_000_181, w_000_090);
  and2 I001_108(w_001_108, w_000_182, w_000_183);
  and2 I001_109(w_001_109, w_000_107, w_000_184);
  and2 I001_110(w_001_110, w_000_179, w_000_185);
  nand2 I001_111(w_001_111, w_000_186, w_000_187);
  and2 I001_112(w_001_112, w_000_188, w_000_009);
  nand2 I001_114(w_001_114, w_000_191, w_000_192);
  or2  I001_115(w_001_115, w_000_193, w_000_194);
  nand2 I001_118(w_001_118, w_000_199, w_000_200);
  or2  I001_119(w_001_119, w_000_201, w_000_127);
  not1 I001_120(w_001_120, w_000_202);
  not1 I001_121(w_001_121, w_000_203);
  and2 I001_122(w_001_122, w_000_204, w_000_205);
  and2 I001_123(w_001_123, w_000_081, w_000_206);
  and2 I001_124(w_001_124, w_000_207, w_000_208);
  and2 I001_125(w_001_125, w_000_209, w_000_210);
  or2  I001_126(w_001_126, w_000_211, w_000_212);
  and2 I001_127(w_001_127, w_000_042, w_000_213);
  or2  I001_128(w_001_128, w_000_214, w_000_190);
  and2 I001_129(w_001_129, w_000_215, w_000_209);
  or2  I001_130(w_001_130, w_000_216, w_000_217);
  and2 I001_131(w_001_131, w_000_155, w_000_218);
  and2 I001_132(w_001_132, w_000_219, w_000_220);
  or2  I001_133(w_001_133, w_000_221, w_000_222);
  nand2 I001_134(w_001_134, w_000_223, w_000_142);
  or2  I001_136(w_001_136, w_000_226, w_000_227);
  not1 I001_138(w_001_138, w_000_230);
  nand2 I001_139(w_001_139, w_000_231, w_000_202);
  not1 I001_140(w_001_140, w_000_232);
  and2 I001_141(w_001_141, w_000_021, w_000_233);
  and2 I001_142(w_001_142, w_000_234, w_000_189);
  and2 I001_143(w_001_143, w_000_235, w_000_236);
  not1 I001_144(w_001_144, w_000_036);
  nand2 I001_146(w_001_146, w_000_239, w_000_133);
  and2 I001_147(w_001_147, w_000_240, w_000_241);
  nand2 I001_148(w_001_148, w_000_242, w_000_243);
  or2  I001_149(w_001_149, w_000_244, w_000_046);
  and2 I001_150(w_001_150, w_000_245, w_000_246);
  not1 I001_151(w_001_151, w_000_247);
  or2  I001_152(w_001_152, w_000_248, w_000_249);
  or2  I001_154(w_001_154, w_000_152, w_000_252);
  nand2 I001_155(w_001_155, w_000_188, w_000_157);
  or2  I001_156(w_001_156, w_000_253, w_000_254);
  not1 I001_157(w_001_157, w_000_255);
  and2 I001_158(w_001_158, w_000_256, w_000_028);
  and2 I001_160(w_001_160, w_000_258, w_000_259);
  nand2 I001_163(w_001_163, w_000_262, w_000_263);
  nand2 I001_164(w_001_164, w_000_264, w_000_159);
  nand2 I001_165(w_001_165, w_000_265, w_000_134);
  nand2 I001_167(w_001_167, w_000_267, w_000_268);
  or2  I001_168(w_001_168, w_000_269, w_000_270);
  or2  I001_170(w_001_170, w_000_273, w_000_238);
  nand2 I001_171(w_001_171, w_000_274, w_000_275);
  nand2 I001_173(w_001_173, w_000_278, w_000_144);
  or2  I001_174(w_001_174, w_000_279, w_000_280);
  and2 I001_175(w_001_175, w_000_281, w_000_282);
  not1 I001_176(w_001_176, w_000_232);
  or2  I001_177(w_001_177, w_000_042, w_000_283);
  or2  I001_178(w_001_178, w_000_023, w_000_284);
  or2  I001_179(w_001_179, w_000_285, w_000_190);
  or2  I001_180(w_001_180, w_000_286, w_000_287);
  or2  I001_181(w_001_181, w_000_234, w_000_288);
  not1 I001_182(w_001_182, w_000_289);
  or2  I001_184(w_001_184, w_000_291, w_000_292);
  not1 I001_186(w_001_186, w_000_293);
  not1 I001_187(w_001_187, w_000_294);
  and2 I001_188(w_001_188, w_000_295, w_000_296);
  not1 I001_189(w_001_189, w_000_290);
  nand2 I001_190(w_001_190, w_000_297, w_000_051);
  and2 I001_191(w_001_191, w_000_298, w_000_299);
  or2  I001_192(w_001_192, w_000_300, w_000_301);
  not1 I001_193(w_001_193, w_000_214);
  nand2 I001_194(w_001_194, w_000_302, w_000_090);
  and2 I001_195(w_001_195, w_000_303, w_000_304);
  or2  I001_196(w_001_196, w_000_189, w_000_274);
  nand2 I001_197(w_001_197, w_000_305, w_000_306);
  or2  I001_198(w_001_198, w_000_307, w_000_308);
  not1 I001_199(w_001_199, w_000_309);
  and2 I001_201(w_001_201, w_000_310, w_000_311);
  and2 I001_202(w_001_202, w_000_312, w_000_237);
  or2  I001_203(w_001_203, w_000_059, w_000_217);
  nand2 I001_205(w_001_205, w_000_314, w_000_315);
  or2  I001_206(w_001_206, w_000_316, w_000_289);
  nand2 I001_207(w_001_207, w_000_317, w_000_318);
  not1 I001_210(w_001_210, w_000_321);
  or2  I001_211(w_001_211, w_000_322, w_000_074);
  or2  I001_213(w_001_213, w_000_324, w_000_270);
  nand2 I001_214(w_001_214, w_000_325, w_000_326);
  or2  I001_215(w_001_215, w_000_327, w_000_328);
  not1 I001_216(w_001_216, w_000_173);
  nand2 I001_217(w_001_217, w_000_329, w_000_330);
  not1 I001_218(w_001_218, w_000_331);
  and2 I001_219(w_001_219, w_000_332, w_000_057);
  not1 I001_221(w_001_221, w_000_334);
  nand2 I001_222(w_001_222, w_000_335, w_000_231);
  not1 I001_224(w_001_224, w_000_030);
  not1 I001_225(w_001_225, w_000_325);
  or2  I001_226(w_001_226, w_000_338, w_000_339);
  nand2 I001_228(w_001_228, w_000_340, w_000_341);
  not1 I001_229(w_001_229, w_000_342);
  not1 I001_230(w_001_230, w_000_021);
  not1 I001_231(w_001_231, w_000_343);
  or2  I001_233(w_001_233, w_000_346, w_000_347);
  and2 I001_234(w_001_234, w_000_348, w_000_207);
  nand2 I001_235(w_001_235, w_000_349, w_000_350);
  nand2 I001_236(w_001_236, w_000_351, w_000_127);
  not1 I001_237(w_001_237, w_000_236);
  and2 I001_238(w_001_238, w_000_352, w_000_105);
  nand2 I001_239(w_001_239, w_000_049, w_000_244);
  nand2 I001_241(w_001_241, w_000_355, w_000_356);
  and2 I001_243(w_001_243, w_000_358, w_000_359);
  or2  I001_244(w_001_244, w_000_360, w_000_361);
  not1 I001_245(w_001_245, w_000_362);
  not1 I001_246(w_001_246, w_000_093);
  not1 I001_247(w_001_247, w_000_126);
  nand2 I001_249(w_001_249, w_000_074, w_000_364);
  or2  I001_250(w_001_250, w_000_179, w_000_365);
  not1 I001_251(w_001_251, w_000_366);
  and2 I001_253(w_001_253, w_000_294, w_000_017);
  or2  I001_255(w_001_255, w_000_369, w_000_153);
  nand2 I001_256(w_001_256, w_000_370, w_000_328);
  or2  I001_257(w_001_257, w_000_291, w_000_371);
  and2 I001_259(w_001_259, w_000_372, w_000_055);
  not1 I001_260(w_001_260, w_000_373);
  not1 I001_261(w_001_261, w_000_374);
  or2  I001_263(w_001_263, w_000_377, w_000_073);
  and2 I001_264(w_001_264, w_000_378, w_000_379);
  not1 I001_265(w_001_265, w_000_380);
  nand2 I001_266(w_001_266, w_000_381, w_000_006);
  nand2 I001_267(w_001_267, w_000_382, w_000_383);
  and2 I001_268(w_001_268, w_000_384, w_000_226);
  nand2 I001_269(w_001_269, w_000_385, w_000_386);
  or2  I001_270(w_001_270, w_000_387, w_000_388);
  and2 I001_271(w_001_271, w_000_389, w_000_390);
  and2 I001_274(w_001_274, w_000_379, w_000_321);
  not1 I001_275(w_001_275, w_000_392);
  and2 I001_276(w_001_276, w_000_393, w_000_234);
  and2 I001_277(w_001_277, w_000_283, w_000_072);
  not1 I001_278(w_001_278, w_000_394);
  nand2 I001_279(w_001_279, w_000_347, w_000_395);
  not1 I001_280(w_001_280, w_000_396);
  not1 I001_281(w_001_281, w_000_059);
  not1 I001_282(w_001_282, w_000_047);
  and2 I001_283(w_001_283, w_000_082, w_000_397);
  and2 I001_284(w_001_284, w_000_204, w_000_398);
  nand2 I001_285(w_001_285, w_000_399, w_000_400);
  and2 I001_286(w_001_286, w_000_278, w_000_159);
  not1 I001_287(w_001_287, w_000_262);
  nand2 I001_288(w_001_288, w_000_041, w_000_401);
  not1 I001_290(w_001_290, w_000_154);
  nand2 I001_291(w_001_291, w_000_402, w_000_403);
  and2 I001_293(w_001_293, w_000_269, w_000_218);
  or2  I001_295(w_001_295, w_000_407, w_000_408);
  and2 I001_296(w_001_296, w_000_409, w_000_410);
  and2 I001_297(w_001_297, w_000_084, w_000_308);
  nand2 I001_299(w_001_299, w_000_376, w_000_412);
  nand2 I001_300(w_001_300, w_000_052, w_000_171);
  or2  I001_301(w_001_301, w_000_413, w_000_414);
  and2 I001_303(w_001_303, w_000_109, w_000_415);
  and2 I001_304(w_001_304, w_000_378, w_000_109);
  or2  I001_305(w_001_305, w_000_081, w_000_114);
  not1 I001_306(w_001_306, w_000_416);
  not1 I001_307(w_001_307, w_000_067);
  nand2 I001_308(w_001_308, w_000_223, w_000_417);
  or2  I001_310(w_001_310, w_000_419, w_000_420);
  nand2 I001_311(w_001_311, w_000_421, w_000_254);
  not1 I001_312(w_001_312, w_000_131);
  or2  I001_313(w_001_313, w_000_422, w_000_423);
  or2  I001_314(w_001_314, w_000_081, w_000_424);
  or2  I001_316(w_001_316, w_000_427, w_000_415);
  and2 I001_317(w_001_317, w_000_428, w_000_404);
  not1 I001_318(w_001_318, w_000_429);
  nand2 I001_319(w_001_319, w_000_297, w_000_032);
  not1 I001_320(w_001_320, w_000_181);
  not1 I001_321(w_001_321, w_000_415);
  or2  I001_322(w_001_322, w_000_430, w_000_431);
  nand2 I001_323(w_001_323, w_000_432, w_000_297);
  nand2 I001_324(w_001_324, w_000_433, w_000_154);
  or2  I001_325(w_001_325, w_000_309, w_000_434);
  and2 I001_326(w_001_326, w_000_382, w_000_021);
  not1 I001_327(w_001_327, w_000_435);
  and2 I001_328(w_001_328, w_000_436, w_000_211);
  or2  I001_329(w_001_329, w_000_086, w_000_285);
  not1 I001_330(w_001_330, w_000_437);
  and2 I001_332(w_001_332, w_000_439, w_000_440);
  or2  I001_333(w_001_333, w_000_441, w_000_442);
  or2  I001_334(w_001_334, w_000_443, w_000_136);
  and2 I001_335(w_001_335, w_000_444, w_000_445);
  not1 I001_339(w_001_339, w_000_437);
  or2  I001_340(w_001_340, w_000_008, w_000_450);
  nand2 I001_341(w_001_341, w_000_350, w_000_451);
  or2  I001_342(w_001_342, w_000_452, w_000_126);
  or2  I001_343(w_001_343, w_000_071, w_000_453);
  nand2 I001_345(w_001_345, w_000_398, w_000_456);
  not1 I001_346(w_001_346, w_000_393);
  or2  I001_347(w_001_347, w_000_457, w_000_458);
  nand2 I001_348(w_001_348, w_000_459, w_000_460);
  nand2 I001_349(w_001_349, w_000_461, w_000_099);
  or2  I001_350(w_001_350, w_000_462, w_000_463);
  or2  I001_351(w_001_351, w_000_464, w_000_465);
  and2 I001_352(w_001_352, w_000_298, w_000_184);
  nand2 I001_353(w_001_353, w_000_466, w_000_467);
  not1 I001_354(w_001_354, w_000_428);
  not1 I001_355(w_001_355, w_000_468);
  and2 I001_356(w_001_356, w_000_469, w_000_278);
  or2  I001_357(w_001_357, w_000_470, w_000_471);
  not1 I001_358(w_001_358, w_000_445);
  nand2 I001_360(w_001_360, w_000_412, w_000_127);
  not1 I001_361(w_001_361, w_000_421);
  or2  I001_362(w_001_362, w_000_334, w_000_439);
  not1 I001_363(w_001_363, w_000_421);
  not1 I001_365(w_001_365, w_000_475);
  not1 I001_366(w_001_366, w_000_476);
  or2  I001_367(w_001_367, w_000_477, w_000_478);
  not1 I001_368(w_001_368, w_000_479);
  not1 I001_369(w_001_369, w_000_399);
  or2  I001_370(w_001_370, w_000_154, w_000_173);
  nand2 I001_371(w_001_371, w_000_480, w_000_481);
  or2  I001_374(w_001_374, w_000_483, w_000_484);
  nand2 I001_375(w_001_375, w_000_280, w_000_485);
  and2 I001_376(w_001_376, w_000_486, w_000_341);
  not1 I001_377(w_001_377, w_000_352);
  or2  I001_378(w_001_378, w_000_487, w_000_069);
  nand2 I001_380(w_001_380, w_000_112, w_000_300);
  not1 I001_381(w_001_381, w_000_488);
  nand2 I001_382(w_001_382, w_000_364, w_000_489);
  and2 I001_385(w_001_385, w_000_491, w_000_492);
  and2 I001_387(w_001_387, w_000_494, w_000_495);
  not1 I001_388(w_001_388, w_000_465);
  not1 I001_390(w_001_390, w_000_183);
  nand2 I001_391(w_001_391, w_000_496, w_000_497);
  not1 I001_393(w_001_393, w_000_289);
  or2  I001_394(w_001_394, w_000_499, w_000_500);
  and2 I001_395(w_001_395, w_000_501, w_000_502);
  nand2 I001_396(w_001_396, w_000_503, w_000_313);
  or2  I001_397(w_001_397, w_000_198, w_000_504);
  nand2 I001_398(w_001_398, w_000_155, w_000_505);
  and2 I001_399(w_001_399, w_000_156, w_000_506);
  or2  I001_400(w_001_400, w_000_507, w_000_286);
  nand2 I001_401(w_001_401, w_000_358, w_000_508);
  and2 I001_402(w_001_402, w_000_245, w_000_181);
  or2  I001_403(w_001_403, w_000_509, w_000_323);
  not1 I001_405(w_001_405, w_000_075);
  and2 I001_406(w_001_406, w_000_042, w_000_510);
  nand2 I001_407(w_001_407, w_000_511, w_000_289);
  and2 I001_408(w_001_408, w_000_469, w_000_238);
  nand2 I001_409(w_001_409, w_000_512, w_000_383);
  nand2 I001_410(w_001_410, w_000_133, w_000_343);
  and2 I001_411(w_001_411, w_000_513, w_000_514);
  nand2 I001_412(w_001_412, w_000_515, w_000_011);
  or2  I001_414(w_001_414, w_000_517, w_000_518);
  nand2 I001_415(w_001_415, w_000_002, w_000_174);
  nand2 I001_416(w_001_416, w_000_519, w_000_216);
  nand2 I001_417(w_001_417, w_000_377, w_000_487);
  and2 I001_418(w_001_418, w_000_520, w_000_521);
  or2  I001_420(w_001_420, w_000_522, w_000_496);
  or2  I001_422(w_001_422, w_000_523, w_000_474);
  and2 I001_423(w_001_423, w_000_393, w_000_485);
  or2  I001_425(w_001_425, w_000_524, w_000_525);
  and2 I001_426(w_001_426, w_000_526, w_000_424);
  nand2 I001_427(w_001_427, w_000_280, w_000_527);
  not1 I001_428(w_001_428, w_000_010);
  and2 I001_429(w_001_429, w_000_528, w_000_529);
  or2  I001_430(w_001_430, w_000_140, w_000_530);
  or2  I001_432(w_001_432, w_000_431, w_000_533);
  and2 I001_433(w_001_433, w_000_534, w_000_535);
  not1 I001_435(w_001_435, w_000_421);
  nand2 I001_436(w_001_436, w_000_537, w_000_538);
  and2 I001_437(w_001_437, w_000_539, w_000_095);
  nand2 I001_438(w_001_438, w_000_024, w_000_088);
  not1 I001_439(w_001_439, w_000_386);
  or2  I001_440(w_001_440, w_000_232, w_000_540);
  not1 I001_441(w_001_441, w_000_373);
  not1 I001_442(w_001_442, w_000_433);
  nand2 I001_443(w_001_443, w_000_541, w_000_279);
  nand2 I001_445(w_001_445, w_000_351, w_000_339);
  and2 I001_446(w_001_446, w_000_543, w_000_330);
  not1 I001_447(w_001_447, w_000_515);
  or2  I001_448(w_001_448, w_000_544, w_000_186);
  or2  I001_449(w_001_449, w_000_011, w_000_545);
  nand2 I001_451(w_001_451, w_000_547, w_000_548);
  nand2 I001_452(w_001_452, w_000_549, w_000_354);
  and2 I001_453(w_001_453, w_000_124, w_000_139);
  nand2 I001_454(w_001_454, w_000_063, w_000_418);
  or2  I001_455(w_001_455, w_000_550, w_000_269);
  or2  I001_456(w_001_456, w_000_404, w_000_551);
  nand2 I001_457(w_001_457, w_000_552, w_000_553);
  nand2 I001_458(w_001_458, w_000_435, w_000_087);
  or2  I001_459(w_001_459, w_000_554, w_000_450);
  nand2 I001_460(w_001_460, w_000_555, w_000_556);
  not1 I001_462(w_001_462, w_000_205);
  or2  I001_464(w_001_464, w_000_559, w_000_403);
  and2 I001_465(w_001_465, w_000_560, w_000_561);
  not1 I001_466(w_001_466, w_000_562);
  nand2 I001_467(w_001_467, w_000_563, w_000_361);
  and2 I001_468(w_001_468, w_000_378, w_000_447);
  and2 I001_469(w_001_469, w_000_045, w_000_564);
  nand2 I001_470(w_001_470, w_000_565, w_000_551);
  or2  I001_471(w_001_471, w_000_386, w_000_353);
  not1 I001_472(w_001_472, w_000_566);
  not1 I001_473(w_001_473, w_000_036);
  not1 I001_474(w_001_474, w_000_107);
  and2 I001_475(w_001_475, w_000_417, w_000_567);
  or2  I001_476(w_001_476, w_000_568, w_000_480);
  not1 I001_477(w_001_477, w_000_569);
  not1 I001_478(w_001_478, w_000_123);
  or2  I001_479(w_001_479, w_000_570, w_000_484);
  or2  I001_480(w_001_480, w_000_312, w_000_571);
  or2  I001_481(w_001_481, w_000_572, w_000_165);
  and2 I001_482(w_001_482, w_000_573, w_000_069);
  or2  I001_483(w_001_483, w_000_574, w_000_422);
  nand2 I001_484(w_001_484, w_000_295, w_000_569);
  nand2 I001_485(w_001_485, w_000_575, w_000_576);
  and2 I001_486(w_001_486, w_000_571, w_000_340);
  or2  I001_487(w_001_487, w_000_577, w_000_172);
  nand2 I001_488(w_001_488, w_000_089, w_000_527);
  not1 I001_489(w_001_489, w_000_578);
  and2 I001_490(w_001_490, w_000_050, w_000_196);
  and2 I001_491(w_001_491, w_000_333, w_000_213);
  not1 I001_492(w_001_492, w_000_499);
  not1 I001_493(w_001_493, w_000_579);
  and2 I001_494(w_001_494, w_000_115, w_000_141);
  not1 I001_495(w_001_495, w_000_580);
  or2  I001_496(w_001_496, w_000_263, w_000_198);
  not1 I001_497(w_001_497, w_000_581);
  not1 I001_498(w_001_498, w_000_513);
  and2 I001_500(w_001_500, w_000_571, w_000_346);
  nand2 I001_501(w_001_501, w_000_138, w_000_225);
  nand2 I001_502(w_001_502, w_000_540, w_000_421);
  and2 I001_503(w_001_503, w_000_226, w_000_582);
  not1 I001_504(w_001_504, w_000_583);
  and2 I001_505(w_001_505, w_000_584, w_000_585);
  and2 I001_506(w_001_506, w_000_446, w_000_339);
  nand2 I001_507(w_001_507, w_000_586, w_000_587);
  or2  I001_508(w_001_508, w_000_588, w_000_542);
  and2 I001_509(w_001_509, w_000_339, w_000_174);
  and2 I001_510(w_001_510, w_000_589, w_000_330);
  or2  I001_512(w_001_512, w_000_519, w_000_590);
  not1 I001_513(w_001_513, w_000_292);
  and2 I001_514(w_001_514, w_000_591, w_000_279);
  not1 I001_515(w_001_515, w_000_592);
  nand2 I001_516(w_001_516, w_000_295, w_000_593);
  not1 I001_518(w_001_518, w_000_596);
  and2 I001_519(w_001_519, w_000_584, w_000_597);
  or2  I001_521(w_001_521, w_000_496, w_000_440);
  nand2 I001_522(w_001_522, w_000_599, w_000_600);
  and2 I001_523(w_001_523, w_000_601, w_000_602);
  and2 I001_524(w_001_524, w_000_523, w_000_251);
  or2  I001_525(w_001_525, w_000_603, w_000_530);
  not1 I001_527(w_001_527, w_000_302);
  or2  I001_528(w_001_528, w_000_079, w_000_591);
  nand2 I001_529(w_001_529, w_000_407, w_000_484);
  nand2 I001_531(w_001_531, w_000_053, w_000_528);
  nand2 I001_532(w_001_532, w_000_494, w_000_606);
  nand2 I001_533(w_001_533, w_000_581, w_000_123);
  and2 I001_534(w_001_534, w_000_187, w_000_607);
  and2 I001_537(w_001_537, w_000_098, w_000_486);
  not1 I001_538(w_001_538, w_000_609);
  nand2 I001_539(w_001_539, w_000_098, w_000_610);
  not1 I001_540(w_001_540, w_000_505);
  not1 I001_542(w_001_542, w_000_425);
  and2 I001_543(w_001_543, w_000_611, w_000_612);
  not1 I001_544(w_001_544, w_000_613);
  and2 I001_546(w_001_546, w_000_086, w_000_614);
  nand2 I001_547(w_001_547, w_000_615, w_000_616);
  or2  I001_548(w_001_548, w_000_197, w_000_617);
  nand2 I001_549(w_001_549, w_000_035, w_000_618);
  not1 I001_551(w_001_551, w_000_619);
  nand2 I001_553(w_001_553, w_000_325, w_000_620);
  or2  I001_555(w_001_555, w_000_115, w_000_560);
  or2  I001_557(w_001_557, w_000_100, w_000_097);
  and2 I001_558(w_001_558, w_000_329, w_000_349);
  or2  I001_559(w_001_559, w_000_623, w_000_624);
  nand2 I001_561(w_001_561, w_000_626, w_000_627);
  not1 I001_562(w_001_562, w_000_626);
  or2  I001_564(w_001_564, w_000_629, w_000_409);
  not1 I001_565(w_001_565, w_000_515);
  nand2 I001_566(w_001_566, w_000_630, w_000_428);
  and2 I001_567(w_001_567, w_000_631, w_000_613);
  not1 I001_568(w_001_568, w_000_300);
  not1 I001_569(w_001_569, w_000_632);
  or2  I001_570(w_001_570, w_000_633, w_000_100);
  and2 I001_571(w_001_571, w_000_397, w_000_416);
  nand2 I001_572(w_001_572, w_000_634, w_000_544);
  and2 I001_573(w_001_573, w_000_320, w_000_635);
  not1 I001_574(w_001_574, w_000_565);
  not1 I001_575(w_001_575, w_000_499);
  not1 I001_576(w_001_576, w_000_546);
  and2 I001_577(w_001_577, w_000_636, w_000_062);
  nand2 I001_578(w_001_578, w_000_637, w_000_638);
  and2 I001_579(w_001_579, w_000_534, w_000_639);
  not1 I001_580(w_001_580, w_000_640);
  or2  I001_581(w_001_581, w_000_596, w_000_641);
  and2 I001_582(w_001_582, w_000_642, w_000_324);
  nand2 I001_584(w_001_584, w_000_643, w_000_361);
  nand2 I001_585(w_001_585, w_000_037, w_000_187);
  or2  I001_586(w_001_586, w_000_602, w_000_644);
  and2 I001_587(w_001_587, w_000_088, w_000_645);
  and2 I001_589(w_001_589, w_000_628, w_000_135);
  and2 I001_590(w_001_590, w_000_162, w_000_647);
  not1 I001_591(w_001_591, w_000_648);
  nand2 I001_592(w_001_592, w_000_466, w_000_649);
  and2 I001_593(w_001_593, w_000_515, w_000_487);
  not1 I001_595(w_001_595, w_000_650);
  and2 I001_597(w_001_597, w_000_494, w_000_293);
  or2  I001_598(w_001_598, w_000_651, w_000_382);
  and2 I001_599(w_001_599, w_000_475, w_000_323);
  not1 I001_600(w_001_600, w_000_652);
  nand2 I001_601(w_001_601, w_000_653, w_000_654);
  or2  I001_602(w_001_602, w_000_168, w_000_655);
  or2  I001_603(w_001_603, w_000_656, w_000_499);
  or2  I001_604(w_001_604, w_000_535, w_000_014);
  and2 I001_605(w_001_605, w_000_657, w_000_346);
  nand2 I001_606(w_001_606, w_000_072, w_000_391);
  and2 I001_607(w_001_607, w_000_411, w_000_623);
  nand2 I001_608(w_001_608, w_000_057, w_000_658);
  or2  I001_609(w_001_609, w_000_439, w_000_281);
  nand2 I001_611(w_001_611, w_000_418, w_000_596);
  not1 I001_612(w_001_612, w_000_659);
  and2 I001_613(w_001_613, w_000_567, w_000_660);
  and2 I001_614(w_001_614, w_000_067, w_000_661);
  nand2 I001_615(w_001_615, w_000_433, w_000_490);
  or2  I001_616(w_001_616, w_000_132, w_000_662);
  or2  I001_617(w_001_617, w_000_523, w_000_663);
  and2 I001_618(w_001_618, w_000_147, w_000_629);
  or2  I001_619(w_001_619, w_000_335, w_000_422);
  and2 I001_620(w_001_620, w_000_664, w_000_043);
  or2  I001_622(w_001_622, w_000_666, w_000_653);
  and2 I001_623(w_001_623, w_000_052, w_000_220);
  or2  I001_624(w_001_624, w_000_204, w_000_287);
  nand2 I001_625(w_001_625, w_000_540, w_000_667);
  or2  I001_627(w_001_627, w_000_127, w_000_669);
  nand2 I001_629(w_001_629, w_000_670, w_000_520);
  nand2 I001_631(w_001_631, w_000_616, w_000_267);
  nand2 I001_632(w_001_632, w_000_382, w_000_292);
  nand2 I001_633(w_001_633, w_000_035, w_000_553);
  nand2 I001_634(w_001_634, w_000_608, w_000_671);
  and2 I001_635(w_001_635, w_000_672, w_000_198);
  and2 I001_636(w_001_636, w_000_673, w_000_376);
  or2  I001_637(w_001_637, w_000_173, w_000_503);
  nand2 I001_638(w_001_638, w_000_254, w_000_673);
  or2  I001_639(w_001_639, w_000_481, w_000_674);
  or2  I001_640(w_001_640, w_000_396, w_000_044);
  not1 I001_641(w_001_641, w_000_280);
  and2 I001_642(w_001_642, w_000_209, w_000_675);
  not1 I001_644(w_001_644, w_000_677);
  or2  I001_645(w_001_645, w_000_678, w_000_679);
  or2  I001_647(w_001_647, w_000_680, w_000_681);
  and2 I001_650(w_001_650, w_000_071, w_000_682);
  and2 I001_652(w_001_652, w_000_683, w_000_684);
  and2 I001_653(w_001_653, w_000_504, w_000_685);
  nand2 I001_654(w_001_654, w_000_358, w_000_525);
  not1 I001_655(w_001_655, w_000_117);
  not1 I001_656(w_001_656, w_000_636);
  not1 I001_657(w_001_657, w_000_560);
  not1 I001_658(w_001_658, w_000_614);
  or2  I001_659(w_001_659, w_000_686, w_000_687);
  or2  I001_661(w_001_661, w_000_688, w_000_400);
  and2 I001_662(w_001_662, w_000_689, w_000_004);
  or2  I001_663(w_001_663, w_000_458, w_000_356);
  nand2 I001_665(w_001_665, w_000_569, w_000_128);
  or2  I001_666(w_001_666, w_000_446, w_000_374);
  not1 I001_667(w_001_667, w_000_605);
  or2  I001_669(w_001_669, w_000_691, w_000_692);
  not1 I001_670(w_001_670, w_000_693);
  and2 I001_671(w_001_671, w_000_238, w_000_694);
  or2  I001_672(w_001_672, w_000_000, w_000_562);
  or2  I001_673(w_001_673, w_000_695, w_000_348);
  or2  I001_674(w_001_674, w_000_017, w_000_696);
  or2  I001_675(w_001_675, w_000_497, w_000_569);
  nand2 I001_677(w_001_677, w_000_018, w_000_470);
  or2  I001_678(w_001_678, w_000_392, w_000_280);
  not1 I001_679(w_001_679, w_000_697);
  or2  I001_680(w_001_680, w_000_698, w_000_699);
  and2 I001_681(w_001_681, w_000_550, w_000_021);
  not1 I001_683(w_001_683, w_000_140);
  not1 I001_684(w_001_684, w_000_647);
  or2  I001_685(w_001_685, w_000_702, w_000_461);
  not1 I001_686(w_001_686, w_000_142);
  not1 I001_687(w_001_687, w_000_191);
  nand2 I001_688(w_001_688, w_000_520, w_000_320);
  not1 I001_689(w_001_689, w_000_538);
  not1 I001_690(w_001_690, w_000_492);
  not1 I001_691(w_001_691, w_000_422);
  not1 I001_692(w_001_692, w_000_685);
  and2 I001_694(w_001_694, w_000_644, w_000_704);
  or2  I001_695(w_001_695, w_000_705, w_000_522);
  nand2 I001_696(w_001_696, w_000_706, w_000_157);
  nand2 I001_697(w_001_697, w_000_602, w_000_492);
  and2 I001_698(w_001_698, w_000_296, w_000_707);
  or2  I001_700(w_001_700, w_000_051, w_000_512);
  and2 I001_701(w_001_701, w_000_589, w_000_654);
  and2 I001_702(w_001_702, w_000_709, w_000_428);
  not1 I001_703(w_001_703, w_000_557);
  and2 I001_704(w_001_704, w_000_576, w_000_337);
  not1 I001_706(w_001_706, w_000_005);
  not1 I001_707(w_001_707, w_000_710);
  or2  I001_709(w_001_709, w_000_236, w_000_015);
  or2  I001_710(w_001_710, w_000_711, w_000_353);
  nand2 I001_711(w_001_711, w_000_712, w_000_713);
  not1 I001_712(w_001_712, w_000_236);
  not1 I001_713(w_001_713, w_000_292);
  not1 I001_714(w_001_714, w_000_158);
  or2  I001_716(w_001_716, w_000_111, w_000_569);
  not1 I001_717(w_001_717, w_000_260);
  not1 I001_718(w_001_718, w_000_714);
  nand2 I001_719(w_001_719, w_000_147, w_000_715);
  or2  I001_720(w_001_720, w_000_716, w_000_439);
  not1 I001_721(w_001_721, w_000_017);
  not1 I001_722(w_001_722, w_000_375);
  or2  I001_723(w_001_723, w_000_511, w_000_674);
  or2  I001_725(w_001_725, w_000_566, w_000_717);
  or2  I001_726(w_001_726, w_000_161, w_000_134);
  or2  I001_727(w_001_727, w_000_536, w_000_127);
  not1 I001_728(w_001_728, w_000_718);
  or2  I001_729(w_001_729, w_000_316, w_000_260);
  nand2 I001_730(w_001_730, w_000_570, w_000_567);
  not1 I001_731(w_001_731, w_000_486);
  and2 I001_732(w_001_732, w_000_719, w_000_277);
  nand2 I001_734(w_001_734, w_000_693, w_000_037);
  not1 I001_737(w_001_737, w_000_540);
  or2  I001_738(w_001_738, w_000_095, w_000_674);
  or2  I001_742(w_001_742, w_000_242, w_000_690);
  nand2 I001_743(w_001_743, w_000_161, w_000_676);
  not1 I001_744(w_001_744, w_000_169);
  nand2 I001_745(w_001_745, w_000_563, w_000_135);
  nand2 I001_746(w_001_746, w_000_351, w_000_180);
  and2 I001_748(w_001_748, w_000_722, w_000_723);
  not1 I001_750(w_001_750, w_000_069);
  and2 I001_751(w_001_751, w_000_416, w_000_052);
  not1 I001_752(w_001_752, w_000_625);
  not1 I001_753(w_001_753, w_000_433);
  nand2 I001_755(w_001_755, w_000_724, w_000_725);
  nand2 I001_756(w_001_756, w_000_235, w_000_726);
  not1 I001_757(w_001_757, w_000_727);
  and2 I001_759(w_001_759, w_000_549, w_000_728);
  and2 I001_760(w_001_760, w_000_589, w_000_013);
  and2 I001_761(w_001_761, w_000_563, w_000_729);
  not1 I001_762(w_001_762, w_000_730);
  not1 I001_763(w_001_763, w_000_731);
  and2 I001_764(w_001_764, w_000_732, w_000_384);
  nand2 I001_765(w_001_765, w_000_209, w_000_238);
  and2 I001_766(w_001_766, w_000_684, w_000_539);
  not1 I001_767(w_001_767, w_000_733);
  nand2 I001_768(w_001_768, w_000_450, w_000_734);
  not1 I001_769(w_001_769, w_000_250);
  not1 I001_770(w_001_770, w_000_428);
  not1 I001_771(w_001_771, w_000_264);
  nand2 I001_772(w_001_772, w_000_735, w_000_736);
  and2 I001_773(w_001_773, w_000_634, w_000_737);
  nand2 I001_774(w_001_774, w_000_738, w_000_105);
  or2  I001_775(w_001_775, w_000_736, w_000_142);
  or2  I001_777(w_001_777, w_000_595, w_000_710);
  or2  I001_778(w_001_778, w_000_632, w_000_249);
  nand2 I001_779(w_001_779, w_000_467, w_000_376);
  not1 I001_780(w_001_780, w_000_601);
  nand2 I001_782(w_001_782, w_000_082, w_000_038);
  nand2 I001_783(w_001_783, w_000_014, w_000_739);
  or2  I001_784(w_001_784, w_000_740, w_000_430);
  not1 I001_785(w_001_785, w_000_669);
  nand2 I001_786(w_001_786, w_000_659, w_000_741);
  nand2 I001_787(w_001_787, w_000_742, w_000_313);
  nand2 I001_788(w_001_788, w_000_718, w_000_260);
  or2  I001_789(w_001_789, w_000_335, w_000_743);
  nand2 I001_790(w_001_790, w_000_443, w_000_712);
  nand2 I001_791(w_001_791, w_000_353, w_000_313);
  not1 I001_792(w_001_792, w_000_513);
  and2 I001_793(w_001_793, w_000_096, w_000_551);
  and2 I001_794(w_001_794, w_000_110, w_000_699);
  nand2 I001_796(w_001_796, w_000_090, w_000_744);
  not1 I001_797(w_001_797, w_000_369);
  and2 I001_798(w_001_798, w_000_008, w_000_682);
  and2 I001_799(w_001_799, w_000_726, w_000_295);
  or2  I001_800(w_001_800, w_000_414, w_000_187);
  and2 I001_801(w_001_801, w_000_745, w_000_251);
  and2 I001_802(w_001_802, w_000_210, w_000_564);
  not1 I001_803(w_001_803, w_000_723);
  or2  I001_804(w_001_804, w_000_746, w_000_626);
  or2  I001_805(w_001_805, w_000_747, w_000_325);
  not1 I001_807(w_001_807, w_000_589);
  not1 I001_809(w_001_809, w_000_749);
  nand2 I001_810(w_001_810, w_000_750, w_000_751);
  not1 I001_811(w_001_811, w_000_155);
  or2  I001_812(w_001_812, w_000_648, w_000_695);
  not1 I001_813(w_001_813, w_000_505);
  not1 I001_814(w_001_814, w_000_366);
  not1 I001_816(w_001_816, w_000_408);
  not1 I001_817(w_001_817, w_000_753);
  or2  I001_818(w_001_818, w_000_235, w_000_093);
  nand2 I001_819(w_001_819, w_000_601, w_000_251);
  and2 I001_820(w_001_820, w_000_410, w_000_651);
  nand2 I001_822(w_001_822, w_000_448, w_000_275);
  or2  I001_824(w_001_824, w_000_651, w_000_755);
  not1 I001_825(w_001_825, w_000_756);
  and2 I001_826(w_001_826, w_000_757, w_000_164);
  and2 I001_827(w_001_827, w_000_043, w_000_572);
  nand2 I001_828(w_001_828, w_000_758, w_000_733);
  not1 I001_829(w_001_829, w_000_256);
  and2 I001_832(w_001_832, w_000_760, w_000_297);
  and2 I001_834(w_001_834, w_000_250, w_000_125);
  or2  I001_835(w_001_835, w_000_253, w_000_319);
  nand2 I001_838(w_001_838, w_000_644, w_000_203);
  not1 I001_839(w_001_839, w_000_729);
  or2  I001_842(w_001_842, w_000_765, w_000_766);
  and2 I001_843(w_001_843, w_000_286, w_000_698);
  or2  I001_844(w_001_844, w_000_513, w_000_344);
  not1 I001_845(w_001_845, w_000_421);
  nand2 I001_846(w_001_846, w_000_207, w_000_658);
  and2 I001_847(w_001_847, w_000_767, w_000_729);
  nand2 I001_848(w_001_848, w_000_758, w_000_053);
  nand2 I001_850(w_001_850, w_000_210, w_000_302);
  not1 I001_852(w_001_852, w_000_769);
  not1 I001_853(w_001_853, w_000_485);
  not1 I001_854(w_001_854, w_000_770);
  or2  I001_856(w_001_856, w_000_501, w_000_772);
  not1 I001_857(w_001_857, w_000_448);
  and2 I001_858(w_001_858, w_000_069, w_000_000);
  nand2 I001_859(w_001_859, w_000_150, w_000_108);
  or2  I001_860(w_001_860, w_000_556, w_000_287);
  and2 I001_861(w_001_861, w_000_328, w_000_462);
  not1 I001_864(w_001_864, w_000_774);
  not1 I001_865(w_001_865, w_000_775);
  nand2 I001_866(w_001_866, w_000_657, w_000_129);
  nand2 I001_867(w_001_867, w_000_294, w_000_630);
  and2 I001_868(w_001_868, w_000_057, w_000_078);
  and2 I001_870(w_001_870, w_000_628, w_000_186);
  or2  I001_871(w_001_871, w_000_184, w_000_776);
  not1 I001_872(w_001_872, w_000_777);
  not1 I001_874(w_001_874, w_000_444);
  or2  I001_876(w_001_876, w_000_589, w_000_283);
  nand2 I001_878(w_001_878, w_000_780, w_000_042);
  or2  I001_880(w_001_880, w_000_428, w_000_550);
  or2  I001_881(w_001_881, w_000_056, w_000_737);
  not1 I001_882(w_001_882, w_000_241);
  not1 I001_883(w_001_883, w_000_782);
  not1 I001_884(w_001_884, w_000_554);
  or2  I001_885(w_001_885, w_000_658, w_000_264);
  not1 I001_886(w_001_886, w_000_281);
  and2 I001_888(w_001_888, w_000_499, w_000_763);
  not1 I001_889(w_001_889, w_000_263);
  not1 I001_890(w_001_890, w_000_399);
  or2  I001_892(w_001_892, w_000_111, w_000_129);
  and2 I001_893(w_001_893, w_000_012, w_000_186);
  or2  I001_894(w_001_894, w_000_055, w_000_779);
  nand2 I001_895(w_001_895, w_000_784, w_000_589);
  or2  I001_896(w_001_896, w_000_089, w_000_247);
  nand2 I002_000(w_002_000, w_000_524, w_001_102);
  and2 I002_001(w_002_001, w_001_114, w_001_326);
  and2 I002_002(w_002_002, w_000_632, w_001_096);
  or2  I002_003(w_002_003, w_000_225, w_001_231);
  nand2 I002_004(w_002_004, w_000_286, w_000_785);
  or2  I002_005(w_002_005, w_001_483, w_000_082);
  not1 I002_007(w_002_007, w_000_680);
  and2 I002_008(w_002_008, w_001_006, w_000_035);
  not1 I002_009(w_002_009, w_001_131);
  and2 I002_010(w_002_010, w_000_709, w_001_825);
  and2 I002_011(w_002_011, w_000_463, w_001_002);
  and2 I002_012(w_002_012, w_000_485, w_001_092);
  not1 I002_013(w_002_013, w_000_656);
  and2 I002_014(w_002_014, w_001_073, w_000_786);
  not1 I002_015(w_002_015, w_001_848);
  not1 I002_016(w_002_016, w_000_787);
  not1 I002_017(w_002_017, w_000_788);
  and2 I002_019(w_002_019, w_000_206, w_000_356);
  or2  I002_020(w_002_020, w_001_847, w_000_789);
  and2 I002_021(w_002_021, w_000_702, w_001_432);
  and2 I002_022(w_002_022, w_001_886, w_001_299);
  and2 I002_023(w_002_023, w_001_489, w_000_539);
  and2 I002_024(w_002_024, w_000_790, w_000_043);
  and2 I002_026(w_002_026, w_000_676, w_001_253);
  nand2 I002_027(w_002_027, w_001_215, w_001_028);
  or2  I002_028(w_002_028, w_001_709, w_001_680);
  nand2 I002_029(w_002_029, w_000_331, w_000_522);
  and2 I002_030(w_002_030, w_000_413, w_000_029);
  and2 I002_031(w_002_031, w_000_424, w_000_448);
  and2 I002_032(w_002_032, w_000_618, w_000_791);
  and2 I002_033(w_002_033, w_001_267, w_001_619);
  or2  I002_034(w_002_034, w_001_848, w_000_770);
  and2 I002_035(w_002_035, w_000_355, w_001_350);
  or2  I002_036(w_002_036, w_001_148, w_000_792);
  or2  I002_038(w_002_038, w_000_303, w_001_470);
  nand2 I002_039(w_002_039, w_001_469, w_000_003);
  and2 I002_040(w_002_040, w_001_064, w_000_526);
  not1 I002_041(w_002_041, w_000_376);
  or2  I002_042(w_002_042, w_001_078, w_000_059);
  not1 I002_043(w_002_043, w_001_399);
  and2 I002_044(w_002_044, w_001_070, w_000_532);
  and2 I002_045(w_002_045, w_000_187, w_000_230);
  not1 I002_046(w_002_046, w_001_051);
  and2 I002_047(w_002_047, w_000_492, w_000_306);
  and2 I002_048(w_002_048, w_000_493, w_001_001);
  not1 I002_049(w_002_049, w_000_793);
  not1 I002_051(w_002_051, w_001_458);
  and2 I002_052(w_002_052, w_001_146, w_000_720);
  not1 I002_053(w_002_053, w_000_014);
  not1 I002_054(w_002_054, w_000_739);
  and2 I002_055(w_002_055, w_000_735, w_001_334);
  or2  I002_056(w_002_056, w_000_635, w_001_546);
  and2 I002_057(w_002_057, w_001_055, w_001_037);
  and2 I002_059(w_002_059, w_000_446, w_001_040);
  or2  I002_060(w_002_060, w_001_303, w_001_221);
  not1 I002_061(w_002_061, w_001_775);
  or2  I002_062(w_002_062, w_000_462, w_000_794);
  or2  I002_063(w_002_063, w_001_417, w_001_728);
  and2 I002_064(w_002_064, w_001_766, w_000_795);
  not1 I002_065(w_002_065, w_001_259);
  not1 I002_066(w_002_066, w_001_057);
  nand2 I002_067(w_002_067, w_000_030, w_001_702);
  or2  I002_068(w_002_068, w_000_096, w_001_492);
  not1 I002_069(w_002_069, w_001_306);
  and2 I002_070(w_002_070, w_000_403, w_000_163);
  or2  I002_071(w_002_071, w_000_339, w_000_352);
  or2  I002_072(w_002_072, w_001_818, w_000_504);
  or2  I002_073(w_002_073, w_000_796, w_000_302);
  and2 I002_074(w_002_074, w_001_004, w_001_256);
  or2  I002_075(w_002_075, w_000_748, w_001_050);
  not1 I002_076(w_002_076, w_001_796);
  or2  I002_077(w_002_077, w_001_311, w_000_680);
  not1 I002_078(w_002_078, w_000_032);
  and2 I002_079(w_002_079, w_001_203, w_000_661);
  and2 I002_080(w_002_080, w_000_797, w_000_553);
  nand2 I002_081(w_002_081, w_000_557, w_000_048);
  not1 I002_082(w_002_082, w_001_148);
  not1 I002_085(w_002_085, w_000_139);
  not1 I002_086(w_002_086, w_000_342);
  or2  I002_087(w_002_087, w_001_005, w_001_704);
  not1 I002_088(w_002_088, w_000_575);
  not1 I002_089(w_002_089, w_000_160);
  not1 I002_090(w_002_090, w_000_623);
  not1 I002_091(w_002_091, w_000_488);
  and2 I002_092(w_002_092, w_001_149, w_000_693);
  or2  I002_093(w_002_093, w_000_448, w_001_360);
  nand2 I002_094(w_002_094, w_000_124, w_001_062);
  not1 I002_096(w_002_096, w_001_167);
  not1 I002_097(w_002_097, w_000_798);
  or2  I002_099(w_002_099, w_001_451, w_001_173);
  not1 I002_100(w_002_100, w_000_585);
  and2 I002_101(w_002_101, w_001_339, w_000_799);
  and2 I002_102(w_002_102, w_001_368, w_000_432);
  and2 I002_104(w_002_104, w_001_571, w_000_794);
  or2  I002_105(w_002_105, w_001_255, w_000_400);
  nand2 I002_106(w_002_106, w_001_573, w_001_157);
  nand2 I002_107(w_002_107, w_001_095, w_000_457);
  not1 I002_108(w_002_108, w_000_801);
  nand2 I002_110(w_002_110, w_000_803, w_000_477);
  or2  I002_111(w_002_111, w_000_271, w_000_287);
  nand2 I002_112(w_002_112, w_000_687, w_000_279);
  and2 I002_114(w_002_114, w_000_066, w_001_229);
  nand2 I002_115(w_002_115, w_000_660, w_001_484);
  or2  I002_116(w_002_116, w_001_329, w_000_203);
  not1 I002_117(w_002_117, w_001_215);
  not1 I002_118(w_002_118, w_000_503);
  or2  I002_119(w_002_119, w_000_542, w_001_500);
  nand2 I002_120(w_002_120, w_000_804, w_001_571);
  or2  I002_121(w_002_121, w_000_638, w_000_187);
  or2  I002_122(w_002_122, w_000_199, w_000_770);
  and2 I002_123(w_002_123, w_001_451, w_000_805);
  not1 I002_124(w_002_124, w_000_098);
  and2 I002_125(w_002_125, w_000_806, w_001_802);
  nand2 I002_126(w_002_126, w_000_654, w_001_614);
  nand2 I002_127(w_002_127, w_000_538, w_000_807);
  and2 I002_128(w_002_128, w_000_483, w_001_422);
  not1 I002_129(w_002_129, w_001_544);
  nand2 I002_130(w_002_130, w_001_099, w_001_247);
  not1 I002_131(w_002_131, w_001_697);
  not1 I002_132(w_002_132, w_001_002);
  nand2 I002_133(w_002_133, w_000_808, w_001_892);
  or2  I002_134(w_002_134, w_001_835, w_001_014);
  nand2 I002_135(w_002_135, w_000_439, w_001_323);
  and2 I002_136(w_002_136, w_001_358, w_000_302);
  or2  I002_137(w_002_137, w_001_650, w_000_690);
  and2 I002_138(w_002_138, w_000_388, w_000_057);
  not1 I002_139(w_002_139, w_001_295);
  and2 I002_140(w_002_140, w_000_540, w_001_141);
  nand2 I002_141(w_002_141, w_001_053, w_001_829);
  and2 I002_142(w_002_142, w_000_152, w_001_316);
  not1 I002_143(w_002_143, w_001_073);
  nand2 I002_144(w_002_144, w_000_809, w_000_040);
  and2 I002_145(w_002_145, w_000_780, w_000_810);
  nand2 I002_146(w_002_146, w_001_479, w_001_019);
  nand2 I002_147(w_002_147, w_001_512, w_000_254);
  or2  I002_148(w_002_148, w_001_083, w_000_528);
  nand2 I002_149(w_002_149, w_001_196, w_000_554);
  not1 I002_150(w_002_150, w_001_256);
  not1 I002_151(w_002_151, w_001_296);
  not1 I002_152(w_002_152, w_001_429);
  and2 I002_153(w_002_153, w_001_600, w_001_718);
  nand2 I002_154(w_002_154, w_000_737, w_000_390);
  not1 I002_156(w_002_156, w_001_257);
  or2  I002_157(w_002_157, w_001_707, w_001_399);
  and2 I002_158(w_002_158, w_001_889, w_000_527);
  nand2 I002_159(w_002_159, w_001_059, w_001_412);
  and2 I002_160(w_002_160, w_000_130, w_000_304);
  nand2 I002_161(w_002_161, w_000_046, w_001_839);
  not1 I002_162(w_002_162, w_000_508);
  and2 I002_163(w_002_163, w_001_765, w_001_130);
  and2 I002_164(w_002_164, w_000_529, w_001_403);
  not1 I002_165(w_002_165, w_001_283);
  or2  I002_166(w_002_166, w_000_591, w_000_069);
  and2 I002_167(w_002_167, w_000_551, w_000_026);
  nand2 I002_168(w_002_168, w_000_072, w_000_811);
  nand2 I002_169(w_002_169, w_000_484, w_001_094);
  or2  I002_170(w_002_170, w_001_473, w_000_812);
  not1 I002_171(w_002_171, w_001_737);
  and2 I002_172(w_002_172, w_000_020, w_001_874);
  nand2 I002_173(w_002_173, w_001_046, w_001_167);
  nand2 I002_174(w_002_174, w_001_193, w_000_780);
  or2  I002_175(w_002_175, w_000_107, w_000_298);
  nand2 I002_176(w_002_176, w_000_289, w_001_817);
  and2 I002_178(w_002_178, w_000_813, w_000_572);
  nand2 I002_179(w_002_179, w_001_446, w_001_538);
  or2  I002_181(w_002_181, w_000_250, w_001_814);
  nand2 I002_182(w_002_182, w_001_024, w_000_765);
  or2  I002_183(w_002_183, w_000_406, w_000_441);
  and2 I002_184(w_002_184, w_001_591, w_000_679);
  nand2 I002_185(w_002_185, w_000_251, w_000_814);
  or2  I002_186(w_002_186, w_001_859, w_001_352);
  and2 I002_187(w_002_187, w_000_386, w_000_815);
  and2 I002_188(w_002_188, w_001_814, w_001_001);
  nand2 I002_189(w_002_189, w_000_816, w_001_396);
  not1 I002_190(w_002_190, w_001_073);
  or2  I002_192(w_002_192, w_001_707, w_001_746);
  or2  I002_193(w_002_193, w_001_605, w_000_653);
  or2  I002_194(w_002_194, w_001_039, w_001_276);
  nand2 I002_195(w_002_195, w_001_091, w_000_130);
  not1 I002_196(w_002_196, w_001_108);
  and2 I002_198(w_002_198, w_001_681, w_001_192);
  or2  I002_199(w_002_199, w_001_042, w_000_370);
  and2 I002_200(w_002_200, w_000_023, w_000_817);
  not1 I002_201(w_002_201, w_001_604);
  or2  I002_202(w_002_202, w_000_695, w_001_069);
  or2  I002_203(w_002_203, w_000_177, w_001_680);
  nand2 I002_204(w_002_204, w_001_257, w_000_766);
  not1 I002_205(w_002_205, w_001_061);
  nand2 I002_206(w_002_206, w_000_249, w_001_224);
  not1 I002_207(w_002_207, w_000_247);
  and2 I002_208(w_002_208, w_001_661, w_001_451);
  not1 I002_209(w_002_209, w_000_498);
  and2 I002_210(w_002_210, w_001_568, w_000_818);
  or2  I002_211(w_002_211, w_000_021, w_000_819);
  or2  I002_212(w_002_212, w_000_196, w_001_777);
  and2 I002_214(w_002_214, w_001_429, w_000_772);
  nand2 I002_215(w_002_215, w_000_576, w_001_886);
  not1 I002_216(w_002_216, w_001_323);
  not1 I002_217(w_002_217, w_000_289);
  and2 I002_218(w_002_218, w_000_662, w_000_424);
  and2 I002_219(w_002_219, w_001_620, w_001_640);
  nand2 I002_220(w_002_220, w_000_018, w_000_222);
  nand2 I002_221(w_002_221, w_001_004, w_001_053);
  nand2 I002_222(w_002_222, w_001_878, w_000_387);
  and2 I002_223(w_002_223, w_000_062, w_001_032);
  nand2 I002_224(w_002_224, w_001_005, w_000_743);
  not1 I002_225(w_002_225, w_000_820);
  not1 I002_226(w_002_226, w_001_053);
  not1 I002_227(w_002_227, w_001_072);
  not1 I002_228(w_002_228, w_000_512);
  and2 I002_229(w_002_229, w_000_821, w_000_255);
  or2  I002_231(w_002_231, w_001_415, w_001_854);
  not1 I002_232(w_002_232, w_000_220);
  not1 I002_233(w_002_233, w_000_270);
  and2 I002_234(w_002_234, w_001_107, w_001_439);
  or2  I002_235(w_002_235, w_000_189, w_001_304);
  or2  I002_236(w_002_236, w_001_151, w_001_011);
  and2 I002_237(w_002_237, w_001_423, w_001_572);
  or2  I002_238(w_002_238, w_000_339, w_000_822);
  and2 I002_240(w_002_240, w_001_789, w_000_710);
  not1 I002_242(w_002_242, w_001_103);
  and2 I002_243(w_002_243, w_000_607, w_001_696);
  nand2 I002_244(w_002_244, w_001_471, w_000_591);
  and2 I002_245(w_002_245, w_000_823, w_001_143);
  and2 I002_246(w_002_246, w_001_662, w_000_334);
  nand2 I002_247(w_002_247, w_001_396, w_000_296);
  or2  I002_248(w_002_248, w_000_096, w_000_824);
  nand2 I002_249(w_002_249, w_000_617, w_000_367);
  or2  I002_250(w_002_250, w_000_386, w_001_074);
  or2  I002_251(w_002_251, w_001_271, w_000_500);
  and2 I002_253(w_002_253, w_001_400, w_001_038);
  or2  I002_254(w_002_254, w_000_334, w_000_386);
  not1 I002_255(w_002_255, w_000_216);
  not1 I002_256(w_002_256, w_000_185);
  and2 I002_257(w_002_257, w_000_825, w_000_826);
  and2 I002_258(w_002_258, w_001_033, w_001_864);
  not1 I002_259(w_002_259, w_000_630);
  not1 I002_260(w_002_260, w_000_762);
  nand2 I002_261(w_002_261, w_000_697, w_001_221);
  or2  I002_262(w_002_262, w_000_620, w_000_442);
  not1 I002_263(w_002_263, w_000_424);
  or2  I002_264(w_002_264, w_001_269, w_001_380);
  nand2 I002_265(w_002_265, w_001_720, w_000_309);
  not1 I002_266(w_002_266, w_000_499);
  and2 I002_267(w_002_267, w_000_038, w_000_827);
  or2  I002_268(w_002_268, w_000_828, w_001_398);
  nand2 I002_269(w_002_269, w_001_370, w_001_457);
  and2 I002_270(w_002_270, w_001_234, w_001_021);
  nand2 I002_271(w_002_271, w_000_753, w_000_829);
  not1 I002_272(w_002_272, w_001_305);
  and2 I002_273(w_002_273, w_001_157, w_000_326);
  nand2 I002_274(w_002_274, w_000_258, w_000_012);
  and2 I002_275(w_002_275, w_001_762, w_000_538);
  and2 I002_276(w_002_276, w_001_348, w_001_307);
  not1 I002_277(w_002_277, w_000_328);
  or2  I002_278(w_002_278, w_001_433, w_001_023);
  nand2 I002_279(w_002_279, w_000_328, w_001_146);
  or2  I002_280(w_002_280, w_001_472, w_000_830);
  not1 I002_281(w_002_281, w_001_196);
  nand2 I002_283(w_002_283, w_000_667, w_000_761);
  or2  I002_284(w_002_284, w_000_441, w_000_397);
  or2  I002_286(w_002_286, w_000_832, w_000_745);
  and2 I002_288(w_002_288, w_000_125, w_001_008);
  nand2 I002_289(w_002_289, w_000_679, w_000_577);
  not1 I002_290(w_002_290, w_000_690);
  nand2 I002_291(w_002_291, w_001_132, w_001_310);
  nand2 I002_292(w_002_292, w_001_083, w_001_507);
  and2 I002_293(w_002_293, w_001_409, w_000_833);
  nand2 I002_294(w_002_294, w_001_021, w_001_377);
  nand2 I002_295(w_002_295, w_001_738, w_000_197);
  or2  I002_296(w_002_296, w_001_774, w_000_834);
  or2  I002_297(w_002_297, w_001_868, w_001_753);
  nand2 I002_298(w_002_298, w_000_835, w_000_801);
  nand2 I002_299(w_002_299, w_000_397, w_000_836);
  not1 I002_300(w_002_300, w_001_126);
  and2 I002_301(w_002_301, w_000_837, w_001_277);
  or2  I002_302(w_002_302, w_001_475, w_001_101);
  or2  I002_303(w_002_303, w_001_306, w_000_542);
  not1 I002_304(w_002_304, w_001_647);
  or2  I002_305(w_002_305, w_001_503, w_001_477);
  not1 I002_306(w_002_306, w_001_226);
  not1 I002_307(w_002_307, w_000_838);
  or2  I002_308(w_002_308, w_000_839, w_000_779);
  nand2 I002_309(w_002_309, w_001_725, w_000_840);
  and2 I002_310(w_002_310, w_001_566, w_001_321);
  and2 I002_311(w_002_311, w_001_495, w_000_757);
  or2  I002_312(w_002_312, w_001_260, w_000_841);
  nand2 I002_313(w_002_313, w_000_082, w_001_788);
  not1 I002_314(w_002_314, w_001_712);
  not1 I002_315(w_002_315, w_001_491);
  or2  I002_316(w_002_316, w_000_216, w_000_497);
  and2 I002_317(w_002_317, w_001_063, w_001_154);
  nand2 I002_318(w_002_318, w_001_001, w_001_090);
  nand2 I002_320(w_002_320, w_001_533, w_001_070);
  nand2 I002_321(w_002_321, w_001_468, w_000_842);
  nand2 I002_322(w_002_322, w_001_760, w_000_843);
  or2  I002_323(w_002_323, w_000_370, w_001_291);
  or2  I002_324(w_002_324, w_001_797, w_001_190);
  nand2 I002_325(w_002_325, w_000_280, w_001_771);
  not1 I002_326(w_002_326, w_000_759);
  and2 I002_327(w_002_327, w_001_181, w_001_050);
  or2  I002_328(w_002_328, w_001_319, w_000_270);
  and2 I002_329(w_002_329, w_001_143, w_001_347);
  not1 I002_330(w_002_330, w_000_639);
  nand2 I002_331(w_002_331, w_001_788, w_000_793);
  and2 I002_333(w_002_333, w_001_063, w_000_567);
  and2 I002_334(w_002_334, w_001_072, w_000_244);
  or2  I002_335(w_002_335, w_000_514, w_001_327);
  or2  I002_336(w_002_336, w_000_675, w_001_876);
  not1 I002_337(w_002_337, w_001_480);
  not1 I002_338(w_002_338, w_001_625);
  not1 I002_339(w_002_339, w_000_403);
  nand2 I002_340(w_002_340, w_001_515, w_000_672);
  nand2 I002_341(w_002_341, w_001_020, w_000_844);
  nand2 I002_342(w_002_342, w_000_586, w_001_624);
  nand2 I002_343(w_002_343, w_001_633, w_001_308);
  or2  I002_344(w_002_344, w_001_077, w_000_845);
  and2 I002_345(w_002_345, w_001_475, w_000_846);
  not1 I002_346(w_002_346, w_001_481);
  or2  I002_347(w_002_347, w_000_153, w_000_541);
  not1 I002_348(w_002_348, w_000_838);
  or2  I002_349(w_002_349, w_000_424, w_001_192);
  nand2 I002_350(w_002_350, w_000_177, w_000_832);
  not1 I002_351(w_002_351, w_000_806);
  not1 I002_352(w_002_352, w_001_586);
  not1 I002_353(w_002_353, w_000_409);
  not1 I002_354(w_002_354, w_000_847);
  nand2 I002_355(w_002_355, w_001_484, w_000_189);
  not1 I002_356(w_002_356, w_001_647);
  and2 I002_357(w_002_357, w_000_215, w_001_455);
  nand2 I002_358(w_002_358, w_000_848, w_001_301);
  nand2 I002_359(w_002_359, w_001_895, w_001_810);
  not1 I002_360(w_002_360, w_000_212);
  or2  I002_361(w_002_361, w_001_486, w_001_235);
  or2  I002_362(w_002_362, w_001_072, w_001_192);
  not1 I002_363(w_002_363, w_000_840);
  not1 I002_364(w_002_364, w_001_055);
  nand2 I002_365(w_002_365, w_000_815, w_000_184);
  or2  I002_367(w_002_367, w_001_077, w_001_101);
  and2 I002_369(w_002_369, w_000_201, w_000_849);
  nand2 I002_370(w_002_370, w_000_080, w_000_559);
  and2 I002_371(w_002_371, w_001_764, w_001_177);
  and2 I002_372(w_002_372, w_001_270, w_001_782);
  not1 I002_373(w_002_373, w_000_672);
  or2  I002_374(w_002_374, w_001_773, w_000_379);
  or2  I002_375(w_002_375, w_001_509, w_001_557);
  not1 I002_376(w_002_376, w_001_446);
  not1 I002_377(w_002_377, w_000_850);
  and2 I002_378(w_002_378, w_001_366, w_001_357);
  or2  I002_379(w_002_379, w_001_657, w_000_625);
  or2  I002_380(w_002_380, w_001_884, w_001_531);
  not1 I002_383(w_002_383, w_000_206);
  and2 I002_384(w_002_384, w_000_085, w_000_354);
  nand2 I002_385(w_002_385, w_001_711, w_001_800);
  or2  I002_386(w_002_386, w_001_426, w_000_704);
  not1 I002_387(w_002_387, w_001_235);
  nand2 I002_388(w_002_388, w_000_540, w_000_649);
  or2  I002_389(w_002_389, w_001_700, w_000_732);
  not1 I002_390(w_002_390, w_001_290);
  not1 I002_391(w_002_391, w_001_375);
  not1 I002_392(w_002_392, w_001_179);
  and2 I002_393(w_002_393, w_001_300, w_000_446);
  or2  I002_394(w_002_394, w_000_824, w_000_300);
  and2 I002_396(w_002_396, w_001_591, w_001_279);
  nand2 I002_397(w_002_397, w_001_094, w_000_602);
  and2 I002_398(w_002_398, w_000_329, w_001_279);
  not1 I002_400(w_002_400, w_000_614);
  not1 I002_401(w_002_401, w_000_852);
  not1 I002_402(w_002_402, w_001_698);
  and2 I002_403(w_002_403, w_001_057, w_001_081);
  or2  I002_404(w_002_404, w_000_037, w_001_684);
  and2 I002_405(w_002_405, w_001_773, w_000_128);
  and2 I002_406(w_002_406, w_001_092, w_001_546);
  nand2 I002_408(w_002_408, w_001_799, w_001_429);
  or2  I002_409(w_002_409, w_001_816, w_001_820);
  not1 I002_410(w_002_410, w_000_058);
  nand2 I002_411(w_002_411, w_001_095, w_001_332);
  and2 I002_412(w_002_412, w_001_813, w_000_853);
  not1 I002_413(w_002_413, w_001_473);
  nand2 I002_414(w_002_414, w_001_525, w_001_442);
  and2 I002_415(w_002_415, w_000_593, w_001_319);
  not1 I002_416(w_002_416, w_000_487);
  or2  I002_417(w_002_417, w_000_633, w_001_777);
  or2  I002_418(w_002_418, w_001_872, w_000_799);
  and2 I002_419(w_002_419, w_000_612, w_000_365);
  not1 I002_420(w_002_420, w_001_190);
  not1 I002_421(w_002_421, w_000_715);
  or2  I002_422(w_002_422, w_000_272, w_001_779);
  or2  I002_423(w_002_423, w_001_221, w_000_582);
  not1 I002_424(w_002_424, w_000_568);
  and2 I002_425(w_002_425, w_001_089, w_001_871);
  nand2 I002_427(w_002_427, w_000_749, w_000_134);
  nand2 I002_428(w_002_428, w_001_202, w_000_854);
  not1 I002_429(w_002_429, w_000_649);
  nand2 I002_430(w_002_430, w_001_222, w_001_157);
  or2  I002_431(w_002_431, w_000_725, w_001_213);
  not1 I002_432(w_002_432, w_000_437);
  and2 I002_433(w_002_433, w_000_752, w_001_717);
  and2 I002_434(w_002_434, w_000_467, w_000_855);
  not1 I002_435(w_002_435, w_001_168);
  not1 I002_437(w_002_437, w_000_856);
  or2  I002_438(w_002_438, w_001_371, w_001_633);
  and2 I002_439(w_002_439, w_001_799, w_000_282);
  nand2 I002_440(w_002_440, w_001_034, w_001_388);
  not1 I002_441(w_002_441, w_001_207);
  or2  I002_442(w_002_442, w_001_494, w_000_258);
  or2  I002_443(w_002_443, w_001_604, w_000_489);
  not1 I002_444(w_002_444, w_000_820);
  and2 I002_445(w_002_445, w_001_191, w_001_246);
  and2 I002_446(w_002_446, w_000_046, w_000_558);
  or2  I002_447(w_002_447, w_001_048, w_000_056);
  nand2 I002_448(w_002_448, w_001_263, w_000_009);
  or2  I002_449(w_002_449, w_001_619, w_000_456);
  nand2 I002_450(w_002_450, w_000_298, w_000_016);
  not1 I002_451(w_002_451, w_000_857);
  or2  I002_452(w_002_452, w_001_228, w_001_818);
  not1 I002_453(w_002_453, w_000_728);
  and2 I002_454(w_002_454, w_001_673, w_000_145);
  or2  I002_455(w_002_455, w_000_409, w_001_505);
  not1 I002_456(w_002_456, w_000_124);
  or2  I002_457(w_002_457, w_001_347, w_001_731);
  or2  I002_458(w_002_458, w_000_849, w_001_478);
  not1 I002_459(w_002_459, w_001_058);
  and2 I002_460(w_002_460, w_001_685, w_000_503);
  or2  I002_461(w_002_461, w_001_529, w_001_593);
  not1 I002_462(w_002_462, w_001_354);
  nand2 I002_463(w_002_463, w_000_224, w_000_518);
  or2  I002_464(w_002_464, w_001_218, w_001_192);
  nand2 I002_465(w_002_465, w_001_041, w_001_551);
  nand2 I002_466(w_002_466, w_000_609, w_001_023);
  not1 I002_467(w_002_467, w_001_878);
  or2  I002_469(w_002_469, w_000_296, w_001_789);
  and2 I002_470(w_002_470, w_001_307, w_000_394);
  or2  I002_471(w_002_471, w_001_586, w_001_019);
  nand2 I002_472(w_002_472, w_000_467, w_000_858);
  and2 I002_473(w_002_473, w_000_315, w_001_078);
  or2  I002_474(w_002_474, w_000_859, w_001_339);
  not1 I002_475(w_002_475, w_000_734);
  not1 I002_476(w_002_476, w_001_523);
  and2 I002_478(w_002_478, w_000_032, w_001_812);
  nand2 I002_479(w_002_479, w_001_631, w_000_149);
  nand2 I002_480(w_002_480, w_000_816, w_000_295);
  not1 I002_482(w_002_482, w_001_746);
  or2  I002_483(w_002_483, w_000_621, w_000_645);
  and2 I002_484(w_002_484, w_001_091, w_000_185);
  and2 I002_485(w_002_485, w_001_349, w_001_590);
  and2 I002_486(w_002_486, w_001_091, w_001_053);
  nand2 I002_487(w_002_487, w_000_701, w_000_847);
  or2  I002_488(w_002_488, w_001_211, w_001_464);
  not1 I002_489(w_002_489, w_000_760);
  nand2 I002_490(w_002_490, w_000_757, w_001_533);
  or2  I002_491(w_002_491, w_001_718, w_001_388);
  nand2 I002_492(w_002_492, w_000_860, w_001_546);
  or2  I002_493(w_002_493, w_001_054, w_000_669);
  and2 I002_494(w_002_494, w_001_868, w_001_884);
  nand2 I002_495(w_002_495, w_001_700, w_001_052);
  and2 I002_496(w_002_496, w_001_194, w_000_112);
  nand2 I002_497(w_002_497, w_001_120, w_000_096);
  or2  I003_000(w_003_000, w_000_839, w_002_308);
  and2 I003_001(w_003_001, w_002_110, w_000_429);
  not1 I003_002(w_003_002, w_001_297);
  and2 I003_003(w_003_003, w_001_728, w_000_474);
  not1 I003_004(w_003_004, w_002_286);
  nand2 I003_005(w_003_005, w_000_856, w_002_106);
  nand2 I003_006(w_003_006, w_002_402, w_000_236);
  nand2 I003_007(w_003_007, w_001_427, w_002_494);
  nand2 I003_008(w_003_008, w_001_604, w_000_073);
  nand2 I003_009(w_003_009, w_002_224, w_000_861);
  nand2 I003_010(w_003_010, w_001_766, w_000_278);
  or2  I003_011(w_003_011, w_000_155, w_001_671);
  nand2 I003_012(w_003_012, w_001_399, w_000_316);
  nand2 I003_013(w_003_013, w_000_004, w_001_721);
  nand2 I003_014(w_003_014, w_001_365, w_001_730);
  nand2 I003_015(w_003_015, w_000_862, w_000_389);
  or2  I003_016(w_003_016, w_002_337, w_000_589);
  and2 I003_017(w_003_017, w_002_005, w_001_622);
  or2  I003_018(w_003_018, w_000_215, w_000_451);
  nand2 I003_019(w_003_019, w_000_583, w_001_829);
  and2 I003_020(w_003_020, w_001_282, w_000_194);
  and2 I003_021(w_003_021, w_001_721, w_000_382);
  not1 I003_022(w_003_022, w_000_051);
  and2 I003_023(w_003_023, w_001_640, w_000_062);
  not1 I003_024(w_003_024, w_002_036);
  nand2 I003_025(w_003_025, w_002_105, w_002_280);
  not1 I003_026(w_003_026, w_002_215);
  not1 I003_027(w_003_027, w_001_872);
  or2  I003_028(w_003_028, w_001_246, w_001_097);
  nand2 I003_029(w_003_029, w_001_255, w_002_345);
  or2  I003_030(w_003_030, w_002_497, w_002_189);
  nand2 I003_031(w_003_031, w_002_337, w_001_856);
  not1 I003_032(w_003_032, w_000_459);
  or2  I003_033(w_003_033, w_000_863, w_001_683);
  and2 I003_034(w_003_034, w_000_864, w_001_515);
  or2  I003_035(w_003_035, w_000_509, w_002_385);
  and2 I003_036(w_003_036, w_001_078, w_002_112);
  not1 I003_037(w_003_037, w_002_301);
  or2  I003_038(w_003_038, w_002_136, w_002_201);
  and2 I003_039(w_003_039, w_002_162, w_002_057);
  not1 I003_040(w_003_040, w_001_590);
  nand2 I003_041(w_003_041, w_001_497, w_001_697);
  not1 I003_042(w_003_042, w_002_061);
  not1 I003_043(w_003_043, w_001_675);
  nand2 I003_044(w_003_044, w_000_145, w_000_010);
  or2  I003_045(w_003_045, w_000_200, w_002_228);
  and2 I003_046(w_003_046, w_001_574, w_002_227);
  nand2 I003_047(w_003_047, w_001_537, w_000_332);
  and2 I003_048(w_003_048, w_002_331, w_002_065);
  nand2 I003_049(w_003_049, w_001_122, w_002_272);
  or2  I003_050(w_003_050, w_001_707, w_000_022);
  or2  I003_051(w_003_051, w_000_115, w_000_681);
  or2  I003_052(w_003_052, w_000_247, w_002_205);
  not1 I003_053(w_003_053, w_001_050);
  and2 I003_054(w_003_054, w_000_632, w_000_056);
  or2  I003_055(w_003_055, w_001_074, w_000_142);
  or2  I003_056(w_003_056, w_002_265, w_001_827);
  and2 I003_057(w_003_057, w_001_202, w_001_205);
  or2  I003_058(w_003_058, w_000_865, w_000_328);
  or2  I003_059(w_003_059, w_000_866, w_000_786);
  or2  I003_060(w_003_060, w_000_867, w_002_264);
  or2  I003_061(w_003_061, w_001_142, w_001_275);
  or2  I003_062(w_003_062, w_001_022, w_002_101);
  or2  I003_063(w_003_063, w_001_094, w_001_267);
  and2 I003_064(w_003_064, w_000_226, w_002_085);
  nand2 I003_065(w_003_065, w_000_213, w_000_287);
  nand2 I003_066(w_003_066, w_002_169, w_002_146);
  and2 I003_067(w_003_067, w_002_279, w_001_127);
  and2 I003_068(w_003_068, w_000_281, w_001_317);
  nand2 I003_069(w_003_069, w_000_543, w_001_031);
  nand2 I003_070(w_003_070, w_000_104, w_000_412);
  nand2 I003_071(w_003_071, w_000_035, w_000_441);
  nand2 I003_072(w_003_072, w_000_770, w_001_284);
  or2  I003_073(w_003_073, w_000_702, w_001_053);
  or2  I003_074(w_003_074, w_000_116, w_001_229);
  not1 I003_075(w_003_075, w_002_359);
  or2  I003_076(w_003_076, w_000_868, w_002_254);
  and2 I003_077(w_003_077, w_000_018, w_001_178);
  or2  I003_078(w_003_078, w_002_121, w_002_240);
  not1 I003_079(w_003_079, w_001_876);
  nand2 I003_080(w_003_080, w_002_433, w_002_102);
  and2 I003_081(w_003_081, w_000_571, w_000_088);
  or2  I003_082(w_003_082, w_002_447, w_001_401);
  not1 I003_083(w_003_083, w_002_157);
  not1 I003_084(w_003_084, w_000_673);
  not1 I003_085(w_003_085, w_001_079);
  not1 I003_086(w_003_086, w_000_159);
  not1 I003_087(w_003_087, w_000_582);
  not1 I003_088(w_003_088, w_001_087);
  or2  I003_089(w_003_089, w_000_086, w_000_584);
  or2  I003_090(w_003_090, w_000_673, w_002_411);
  not1 I003_091(w_003_091, w_001_812);
  and2 I003_092(w_003_092, w_000_468, w_002_203);
  or2  I003_093(w_003_093, w_001_644, w_000_151);
  nand2 I003_094(w_003_094, w_002_293, w_000_018);
  nand2 I003_095(w_003_095, w_002_002, w_000_257);
  or2  I003_096(w_003_096, w_000_842, w_002_256);
  nand2 I003_097(w_003_097, w_002_169, w_002_132);
  and2 I003_098(w_003_098, w_002_420, w_000_385);
  nand2 I003_099(w_003_099, w_000_690, w_002_070);
  or2  I003_100(w_003_100, w_000_506, w_002_245);
  and2 I003_101(w_003_101, w_000_276, w_001_706);
  or2  I003_102(w_003_102, w_002_179, w_001_474);
  not1 I003_103(w_003_103, w_000_347);
  or2  I003_104(w_003_104, w_000_869, w_001_130);
  nand2 I003_105(w_003_105, w_001_515, w_001_287);
  or2  I003_106(w_003_106, w_001_709, w_001_417);
  nand2 I003_107(w_003_107, w_000_512, w_001_681);
  and2 I003_108(w_003_108, w_000_740, w_000_346);
  or2  I003_109(w_003_109, w_002_323, w_000_700);
  and2 I003_110(w_003_110, w_002_484, w_001_498);
  not1 I003_111(w_003_111, w_002_288);
  or2  I003_112(w_003_112, w_001_030, w_002_206);
  and2 I003_113(w_003_113, w_001_078, w_001_024);
  nand2 I003_114(w_003_114, w_000_057, w_002_471);
  or2  I003_115(w_003_115, w_002_169, w_001_111);
  and2 I003_116(w_003_116, w_001_811, w_000_870);
  nand2 I003_117(w_003_117, w_001_482, w_000_604);
  not1 I003_118(w_003_118, w_000_871);
  or2  I003_119(w_003_119, w_000_478, w_000_272);
  or2  I003_120(w_003_120, w_002_296, w_002_238);
  not1 I003_121(w_003_121, w_002_061);
  nand2 I003_122(w_003_122, w_002_227, w_000_038);
  nand2 I003_123(w_003_123, w_002_202, w_001_028);
  or2  I003_124(w_003_124, w_002_012, w_002_394);
  and2 I003_125(w_003_125, w_002_164, w_000_746);
  nand2 I003_126(w_003_126, w_001_018, w_001_366);
  nand2 I003_127(w_003_127, w_001_060, w_000_662);
  and2 I003_128(w_003_128, w_002_443, w_001_595);
  and2 I003_129(w_003_129, w_000_640, w_001_046);
  and2 I003_130(w_003_130, w_002_231, w_001_198);
  nand2 I003_131(w_003_131, w_002_460, w_001_253);
  not1 I003_132(w_003_132, w_001_027);
  and2 I003_133(w_003_133, w_000_746, w_000_824);
  nand2 I003_134(w_003_134, w_001_487, w_002_291);
  and2 I003_135(w_003_135, w_002_238, w_000_872);
  and2 I003_136(w_003_136, w_001_181, w_001_678);
  and2 I003_137(w_003_137, w_000_873, w_000_147);
  and2 I003_138(w_003_138, w_002_254, w_000_161);
  nand2 I003_139(w_003_139, w_000_244, w_000_362);
  or2  I003_140(w_003_140, w_002_129, w_002_358);
  and2 I003_141(w_003_141, w_000_227, w_001_449);
  or2  I003_142(w_003_142, w_001_743, w_002_482);
  or2  I003_143(w_003_143, w_001_260, w_001_650);
  nand2 I003_144(w_003_144, w_001_529, w_000_233);
  nand2 I003_145(w_003_145, w_001_704, w_001_224);
  not1 I003_146(w_003_146, w_000_156);
  or2  I003_147(w_003_147, w_002_364, w_002_009);
  nand2 I003_148(w_003_148, w_000_458, w_000_874);
  or2  I003_149(w_003_149, w_001_234, w_001_522);
  not1 I003_150(w_003_150, w_000_524);
  or2  I003_151(w_003_151, w_002_054, w_002_106);
  or2  I003_152(w_003_152, w_000_660, w_002_188);
  nand2 I003_153(w_003_153, w_000_195, w_000_469);
  nand2 I003_154(w_003_154, w_000_830, w_001_663);
  and2 I003_155(w_003_155, w_001_020, w_002_078);
  nand2 I003_156(w_003_156, w_001_600, w_000_202);
  or2  I003_157(w_003_157, w_001_573, w_001_422);
  not1 I003_158(w_003_158, w_001_236);
  not1 I003_159(w_003_159, w_000_875);
  or2  I003_160(w_003_160, w_000_470, w_000_743);
  or2  I003_161(w_003_161, w_001_028, w_002_403);
  not1 I003_162(w_003_162, w_002_320);
  and2 I003_163(w_003_163, w_002_325, w_000_876);
  and2 I003_164(w_003_164, w_002_416, w_001_112);
  nand2 I003_165(w_003_165, w_002_290, w_000_785);
  or2  I003_166(w_003_166, w_001_060, w_000_877);
  not1 I003_167(w_003_167, w_000_068);
  nand2 I003_168(w_003_168, w_001_096, w_002_494);
  nand2 I003_169(w_003_169, w_002_166, w_001_858);
  and2 I003_170(w_003_170, w_001_149, w_002_401);
  or2  I003_171(w_003_171, w_002_364, w_000_878);
  not1 I003_172(w_003_172, w_001_768);
  nand2 I003_173(w_003_173, w_001_828, w_001_816);
  not1 I003_174(w_003_174, w_001_236);
  not1 I003_175(w_003_175, w_001_581);
  not1 I003_176(w_003_176, w_000_493);
  not1 I003_177(w_003_177, w_000_516);
  and2 I003_178(w_003_178, w_000_877, w_001_128);
  and2 I003_179(w_003_179, w_002_065, w_000_840);
  not1 I003_180(w_003_180, w_000_631);
  nand2 I003_181(w_003_181, w_000_474, w_000_224);
  not1 I003_182(w_003_182, w_000_879);
  not1 I003_183(w_003_183, w_001_634);
  and2 I003_184(w_003_184, w_002_451, w_001_872);
  and2 I003_185(w_003_185, w_000_484, w_000_402);
  not1 I003_186(w_003_186, w_002_033);
  not1 I003_187(w_003_187, w_000_023);
  not1 I003_188(w_003_188, w_000_522);
  or2  I003_189(w_003_189, w_000_157, w_001_011);
  or2  I003_190(w_003_190, w_000_466, w_000_449);
  not1 I003_191(w_003_191, w_000_613);
  and2 I003_192(w_003_192, w_001_270, w_001_260);
  nand2 I003_193(w_003_193, w_001_360, w_002_127);
  and2 I003_194(w_003_194, w_001_053, w_001_104);
  nand2 I003_195(w_003_195, w_001_627, w_000_593);
  and2 I003_196(w_003_196, w_002_355, w_002_363);
  nand2 I003_197(w_003_197, w_001_164, w_001_592);
  or2  I003_198(w_003_198, w_002_220, w_001_044);
  and2 I003_199(w_003_199, w_002_323, w_001_448);
  and2 I003_200(w_003_200, w_002_031, w_001_271);
  not1 I003_201(w_003_201, w_001_803);
  or2  I003_202(w_003_202, w_002_396, w_001_885);
  or2  I003_203(w_003_203, w_001_600, w_000_588);
  and2 I003_204(w_003_204, w_001_181, w_002_044);
  or2  I003_205(w_003_205, w_001_483, w_001_895);
  or2  I003_206(w_003_206, w_002_343, w_002_261);
  or2  I003_207(w_003_207, w_002_386, w_000_131);
  nand2 I003_208(w_003_208, w_000_224, w_002_333);
  not1 I003_209(w_003_209, w_002_007);
  not1 I003_210(w_003_210, w_000_596);
  nand2 I003_211(w_003_211, w_002_129, w_001_202);
  not1 I003_212(w_003_212, w_000_037);
  nand2 I003_213(w_003_213, w_001_694, w_000_307);
  and2 I003_214(w_003_214, w_002_034, w_000_445);
  nand2 I003_215(w_003_215, w_001_484, w_001_319);
  and2 I003_216(w_003_216, w_000_429, w_002_170);
  nand2 I003_217(w_003_217, w_000_264, w_001_030);
  or2  I003_218(w_003_218, w_000_129, w_002_314);
  nand2 I003_219(w_003_219, w_000_776, w_001_098);
  nand2 I003_220(w_003_220, w_000_659, w_001_476);
  and2 I003_221(w_003_221, w_002_425, w_001_743);
  not1 I003_222(w_003_222, w_001_403);
  nand2 I003_223(w_003_223, w_000_071, w_002_439);
  nand2 I003_224(w_003_224, w_001_718, w_002_430);
  and2 I003_225(w_003_225, w_002_242, w_001_016);
  and2 I004_000(w_004_000, w_003_077, w_002_022);
  nand2 I004_001(w_004_001, w_002_478, w_003_197);
  nand2 I004_002(w_004_002, w_002_439, w_000_537);
  not1 I004_003(w_004_003, w_003_157);
  or2  I004_004(w_004_004, w_002_296, w_002_312);
  or2  I004_005(w_004_005, w_002_014, w_000_590);
  nand2 I004_006(w_004_006, w_002_458, w_000_825);
  or2  I004_007(w_004_007, w_002_350, w_001_884);
  not1 I004_008(w_004_008, w_000_082);
  or2  I004_009(w_004_009, w_002_375, w_001_447);
  and2 I004_010(w_004_010, w_000_056, w_001_478);
  or2  I004_011(w_004_011, w_003_113, w_002_141);
  nand2 I004_012(w_004_012, w_002_233, w_003_218);
  or2  I004_013(w_004_013, w_003_044, w_002_459);
  not1 I004_014(w_004_014, w_003_193);
  and2 I004_015(w_004_015, w_003_049, w_002_429);
  or2  I004_016(w_004_016, w_003_199, w_001_019);
  or2  I004_017(w_004_017, w_002_394, w_002_257);
  or2  I004_018(w_004_018, w_000_750, w_001_759);
  or2  I004_019(w_004_019, w_000_203, w_002_225);
  or2  I004_020(w_004_020, w_000_032, w_003_124);
  or2  I004_021(w_004_021, w_000_643, w_001_394);
  or2  I004_022(w_004_022, w_002_425, w_002_101);
  or2  I004_023(w_004_023, w_003_113, w_000_880);
  not1 I004_024(w_004_024, w_001_058);
  and2 I004_025(w_004_025, w_002_169, w_001_138);
  or2  I004_026(w_004_026, w_003_213, w_002_069);
  or2  I004_027(w_004_027, w_002_043, w_003_064);
  nand2 I004_028(w_004_028, w_000_684, w_000_734);
  or2  I004_029(w_004_029, w_002_187, w_003_057);
  not1 I004_030(w_004_030, w_003_113);
  and2 I004_031(w_004_031, w_000_398, w_000_223);
  nand2 I004_032(w_004_032, w_001_361, w_000_348);
  nand2 I004_033(w_004_033, w_003_011, w_000_689);
  nand2 I004_034(w_004_034, w_003_075, w_002_375);
  nand2 I004_035(w_004_035, w_002_461, w_000_881);
  not1 I004_036(w_004_036, w_003_085);
  and2 I004_037(w_004_037, w_002_183, w_000_882);
  nand2 I004_038(w_004_038, w_000_150, w_002_295);
  nand2 I005_000(w_005_000, w_001_790, w_000_409);
  nand2 I005_001(w_005_001, w_004_017, w_002_210);
  not1 I005_002(w_005_002, w_000_225);
  and2 I005_003(w_005_003, w_001_701, w_002_002);
  or2  I005_004(w_005_004, w_003_098, w_002_486);
  nand2 I005_005(w_005_005, w_004_020, w_002_378);
  and2 I005_006(w_005_006, w_001_092, w_000_883);
  not1 I005_007(w_005_007, w_000_303);
  or2  I005_008(w_005_008, w_001_023, w_002_100);
  or2  I005_009(w_005_009, w_002_175, w_003_127);
  and2 I005_010(w_005_010, w_002_305, w_004_035);
  not1 I005_011(w_005_011, w_002_179);
  or2  I005_012(w_005_012, w_003_043, w_000_260);
  nand2 I005_013(w_005_013, w_003_126, w_004_033);
  not1 I005_014(w_005_014, w_001_843);
  and2 I005_015(w_005_015, w_002_369, w_000_325);
  and2 I005_016(w_005_016, w_004_033, w_004_030);
  and2 I005_017(w_005_017, w_001_615, w_000_514);
  or2  I005_018(w_005_018, w_004_037, w_004_019);
  nand2 I005_019(w_005_019, w_004_006, w_000_340);
  not1 I005_020(w_005_020, w_004_022);
  nand2 I005_023(w_005_023, w_002_243, w_004_004);
  nand2 I005_024(w_005_024, w_000_853, w_000_327);
  and2 I005_026(w_005_026, w_002_362, w_000_241);
  or2  I005_028(w_005_028, w_003_018, w_003_091);
  or2  I005_029(w_005_029, w_003_160, w_002_304);
  nand2 I005_030(w_005_030, w_003_040, w_003_125);
  not1 I005_031(w_005_031, w_001_452);
  and2 I005_032(w_005_032, w_000_323, w_003_155);
  or2  I005_033(w_005_033, w_000_201, w_001_847);
  or2  I005_034(w_005_034, w_004_007, w_001_284);
  and2 I005_035(w_005_035, w_001_053, w_004_032);
  or2  I005_036(w_005_036, w_003_115, w_000_026);
  or2  I005_037(w_005_037, w_001_504, w_004_030);
  and2 I005_038(w_005_038, w_002_309, w_002_257);
  nand2 I005_039(w_005_039, w_004_021, w_003_153);
  and2 I005_040(w_005_040, w_004_021, w_004_027);
  not1 I005_042(w_005_042, w_003_205);
  nand2 I005_043(w_005_043, w_003_036, w_001_091);
  not1 I005_045(w_005_045, w_003_171);
  not1 I005_047(w_005_047, w_004_003);
  and2 I005_048(w_005_048, w_001_090, w_001_464);
  or2  I005_049(w_005_049, w_000_885, w_001_020);
  or2  I005_050(w_005_050, w_001_408, w_004_020);
  and2 I005_051(w_005_051, w_000_531, w_001_457);
  and2 I005_053(w_005_053, w_001_760, w_000_825);
  or2  I005_054(w_005_054, w_000_098, w_004_020);
  not1 I005_055(w_005_055, w_004_031);
  and2 I005_056(w_005_056, w_000_831, w_000_203);
  nand2 I005_057(w_005_057, w_000_496, w_004_008);
  and2 I005_058(w_005_058, w_001_442, w_001_613);
  and2 I005_059(w_005_059, w_003_166, w_003_165);
  and2 I005_060(w_005_060, w_000_217, w_000_198);
  nand2 I005_061(w_005_061, w_001_647, w_004_027);
  not1 I005_062(w_005_062, w_001_692);
  not1 I005_063(w_005_063, w_004_038);
  or2  I005_064(w_005_064, w_001_744, w_003_009);
  and2 I005_065(w_005_065, w_004_014, w_001_074);
  not1 I005_066(w_005_066, w_001_466);
  nand2 I005_067(w_005_067, w_004_033, w_001_558);
  and2 I005_069(w_005_069, w_002_096, w_003_008);
  and2 I005_070(w_005_070, w_002_310, w_004_016);
  and2 I005_071(w_005_071, w_002_183, w_004_001);
  not1 I005_072(w_005_072, w_002_279);
  and2 I005_073(w_005_073, w_000_595, w_002_256);
  or2  I005_074(w_005_074, w_001_313, w_004_024);
  nand2 I005_075(w_005_075, w_001_018, w_001_885);
  and2 I005_076(w_005_076, w_004_032, w_000_504);
  not1 I005_078(w_005_078, w_001_319);
  and2 I005_080(w_005_080, w_002_431, w_000_635);
  not1 I005_081(w_005_081, w_004_011);
  or2  I005_082(w_005_082, w_002_389, w_004_003);
  nand2 I005_083(w_005_083, w_001_504, w_001_350);
  or2  I005_084(w_005_084, w_003_199, w_000_337);
  not1 I005_085(w_005_085, w_003_204);
  nand2 I005_086(w_005_086, w_003_105, w_004_035);
  and2 I005_088(w_005_088, w_001_027, w_001_098);
  or2  I005_089(w_005_089, w_000_886, w_002_386);
  or2  I005_090(w_005_090, w_000_887, w_000_245);
  and2 I005_091(w_005_091, w_003_219, w_003_002);
  nand2 I005_092(w_005_092, w_002_161, w_003_004);
  and2 I005_093(w_005_093, w_002_040, w_003_126);
  nand2 I005_094(w_005_094, w_000_032, w_002_293);
  not1 I005_095(w_005_095, w_000_325);
  and2 I005_096(w_005_096, w_000_064, w_002_160);
  not1 I005_097(w_005_097, w_004_016);
  not1 I005_098(w_005_098, w_000_655);
  not1 I005_099(w_005_099, w_002_040);
  and2 I005_100(w_005_100, w_001_396, w_002_045);
  not1 I005_101(w_005_101, w_000_015);
  not1 I005_102(w_005_102, w_003_098);
  nand2 I005_103(w_005_103, w_001_743, w_003_035);
  or2  I005_104(w_005_104, w_001_878, w_000_810);
  nand2 I005_105(w_005_105, w_001_412, w_002_154);
  nand2 I005_106(w_005_106, w_002_102, w_004_030);
  and2 I005_107(w_005_107, w_003_090, w_004_024);
  and2 I005_108(w_005_108, w_000_585, w_002_452);
  nand2 I005_109(w_005_109, w_003_092, w_004_012);
  not1 I005_110(w_005_110, w_000_205);
  nand2 I005_112(w_005_112, w_001_085, w_003_128);
  not1 I005_113(w_005_113, w_003_144);
  not1 I005_114(w_005_114, w_003_008);
  and2 I005_116(w_005_116, w_003_093, w_003_023);
  not1 I005_117(w_005_117, w_001_437);
  not1 I005_118(w_005_118, w_001_277);
  nand2 I005_119(w_005_119, w_001_157, w_000_005);
  or2  I005_120(w_005_120, w_003_138, w_004_025);
  nand2 I005_121(w_005_121, w_001_219, w_004_010);
  not1 I005_123(w_005_123, w_003_077);
  and2 I005_124(w_005_124, w_000_657, w_000_762);
  or2  I005_126(w_005_126, w_002_389, w_004_019);
  nand2 I005_128(w_005_128, w_003_034, w_002_424);
  and2 I005_129(w_005_129, w_002_259, w_001_226);
  and2 I005_131(w_005_131, w_002_168, w_003_143);
  not1 I005_132(w_005_132, w_000_673);
  nand2 I005_133(w_005_133, w_002_415, w_003_152);
  and2 I005_134(w_005_134, w_004_014, w_001_631);
  and2 I005_135(w_005_135, w_001_569, w_003_039);
  or2  I005_136(w_005_136, w_003_072, w_004_025);
  and2 I005_137(w_005_137, w_003_084, w_000_000);
  not1 I005_138(w_005_138, w_004_028);
  and2 I005_139(w_005_139, w_004_014, w_004_020);
  nand2 I005_141(w_005_141, w_004_029, w_004_008);
  not1 I005_142(w_005_142, w_000_163);
  not1 I005_143(w_005_143, w_003_058);
  or2  I005_144(w_005_144, w_003_207, w_003_068);
  and2 I005_145(w_005_145, w_002_012, w_002_467);
  or2  I005_147(w_005_147, w_000_876, w_002_196);
  nand2 I005_148(w_005_148, w_003_093, w_000_889);
  nand2 I005_149(w_005_149, w_003_130, w_001_041);
  not1 I005_150(w_005_150, w_000_445);
  or2  I005_151(w_005_151, w_000_317, w_002_403);
  or2  I005_152(w_005_152, w_004_018, w_001_490);
  or2  I005_153(w_005_153, w_003_028, w_001_801);
  and2 I005_154(w_005_154, w_000_495, w_000_633);
  and2 I005_155(w_005_155, w_002_102, w_002_405);
  not1 I005_156(w_005_156, w_000_447);
  and2 I005_157(w_005_157, w_001_244, w_002_076);
  or2  I005_158(w_005_158, w_004_012, w_000_144);
  nand2 I005_159(w_005_159, w_003_082, w_001_669);
  not1 I005_160(w_005_160, w_004_002);
  not1 I005_161(w_005_161, w_000_890);
  and2 I005_163(w_005_163, w_001_122, w_000_880);
  nand2 I005_164(w_005_164, w_002_181, w_002_190);
  not1 I005_165(w_005_165, w_001_249);
  or2  I005_166(w_005_166, w_002_492, w_001_003);
  and2 I005_167(w_005_167, w_002_456, w_001_040);
  nand2 I005_168(w_005_168, w_001_015, w_000_457);
  not1 I005_169(w_005_169, w_001_267);
  not1 I005_170(w_005_170, w_004_000);
  nand2 I005_171(w_005_171, w_004_029, w_003_068);
  and2 I005_172(w_005_172, w_001_038, w_001_858);
  and2 I005_173(w_005_173, w_000_702, w_001_198);
  not1 I005_174(w_005_174, w_000_654);
  and2 I005_175(w_005_175, w_002_062, w_002_274);
  or2  I005_176(w_005_176, w_001_362, w_000_891);
  and2 I005_177(w_005_177, w_001_088, w_001_793);
  or2  I005_178(w_005_178, w_004_024, w_001_492);
  and2 I005_179(w_005_179, w_002_204, w_002_106);
  and2 I005_180(w_005_180, w_000_803, w_004_028);
  or2  I005_181(w_005_181, w_002_404, w_001_454);
  nand2 I005_184(w_005_184, w_000_438, w_003_134);
  nand2 I005_185(w_005_185, w_001_081, w_003_092);
  or2  I005_186(w_005_186, w_000_374, w_002_106);
  not1 I005_188(w_005_188, w_002_092);
  or2  I005_189(w_005_189, w_000_125, w_001_759);
  nand2 I005_190(w_005_190, w_000_404, w_002_312);
  not1 I005_191(w_005_191, w_000_296);
  and2 I005_193(w_005_193, w_003_150, w_000_596);
  or2  I005_194(w_005_194, w_004_004, w_003_129);
  or2  I005_195(w_005_195, w_003_071, w_004_000);
  and2 I005_196(w_005_196, w_003_189, w_002_335);
  or2  I005_197(w_005_197, w_004_021, w_002_097);
  not1 I005_199(w_005_199, w_004_032);
  not1 I005_200(w_005_200, w_002_130);
  nand2 I005_201(w_005_201, w_003_180, w_004_036);
  or2  I005_202(w_005_202, w_002_078, w_004_020);
  and2 I005_203(w_005_203, w_002_107, w_001_342);
  and2 I005_204(w_005_204, w_003_012, w_000_200);
  nand2 I005_205(w_005_205, w_002_482, w_001_271);
  not1 I005_206(w_005_206, w_003_204);
  and2 I005_207(w_005_207, w_002_138, w_001_590);
  and2 I005_208(w_005_208, w_000_094, w_003_141);
  nand2 I005_210(w_005_210, w_003_195, w_000_197);
  and2 I005_211(w_005_211, w_003_210, w_002_130);
  nand2 I005_212(w_005_212, w_004_034, w_001_792);
  or2  I005_213(w_005_213, w_004_020, w_000_286);
  or2  I005_214(w_005_214, w_001_228, w_002_300);
  or2  I005_216(w_005_216, w_001_564, w_003_220);
  not1 I005_217(w_005_217, w_000_602);
  not1 I005_218(w_005_218, w_002_085);
  or2  I005_219(w_005_219, w_003_096, w_001_662);
  or2  I005_220(w_005_220, w_003_011, w_004_038);
  and2 I005_221(w_005_221, w_002_345, w_001_555);
  not1 I005_223(w_005_223, w_004_021);
  nand2 I005_224(w_005_224, w_003_017, w_002_394);
  nand2 I005_225(w_005_225, w_001_080, w_001_259);
  or2  I005_226(w_005_226, w_002_273, w_000_832);
  and2 I005_227(w_005_227, w_004_013, w_000_504);
  not1 I005_228(w_005_228, w_002_059);
  not1 I005_229(w_005_229, w_001_039);
  nand2 I005_230(w_005_230, w_001_870, w_002_330);
  and2 I005_232(w_005_232, w_004_028, w_004_036);
  nand2 I005_233(w_005_233, w_004_036, w_000_351);
  nand2 I005_234(w_005_234, w_001_652, w_002_040);
  not1 I005_235(w_005_235, w_001_452);
  not1 I005_237(w_005_237, w_000_746);
  nand2 I005_238(w_005_238, w_003_070, w_000_065);
  and2 I005_239(w_005_239, w_001_522, w_004_024);
  or2  I005_240(w_005_240, w_003_093, w_001_251);
  not1 I005_242(w_005_242, w_000_732);
  nand2 I005_243(w_005_243, w_000_472, w_003_148);
  not1 I005_244(w_005_244, w_000_246);
  or2  I005_245(w_005_245, w_000_542, w_003_132);
  nand2 I005_246(w_005_246, w_004_022, w_001_013);
  not1 I005_247(w_005_247, w_001_260);
  not1 I005_248(w_005_248, w_004_007);
  not1 I005_249(w_005_249, w_003_096);
  not1 I005_250(w_005_250, w_003_208);
  nand2 I005_251(w_005_251, w_003_016, w_001_728);
  and2 I005_252(w_005_252, w_001_888, w_000_507);
  not1 I005_253(w_005_253, w_000_133);
  and2 I005_254(w_005_254, w_002_472, w_001_500);
  nand2 I005_256(w_005_256, w_001_460, w_003_020);
  not1 I005_257(w_005_257, w_003_128);
  or2  I005_258(w_005_258, w_001_822, w_004_015);
  not1 I005_259(w_005_259, w_000_606);
  and2 I005_260(w_005_260, w_004_007, w_000_447);
  or2  I005_261(w_005_261, w_004_038, w_000_321);
  nand2 I005_262(w_005_262, w_001_509, w_004_025);
  nand2 I005_264(w_005_264, w_002_355, w_004_024);
  or2  I005_265(w_005_265, w_003_093, w_002_342);
  nand2 I005_266(w_005_266, w_000_155, w_002_227);
  not1 I005_268(w_005_268, w_003_190);
  or2  I005_269(w_005_269, w_002_232, w_004_035);
  nand2 I005_270(w_005_270, w_002_107, w_000_314);
  not1 I005_271(w_005_271, w_002_022);
  not1 I005_272(w_005_272, w_004_005);
  and2 I005_273(w_005_273, w_002_273, w_003_087);
  nand2 I005_274(w_005_274, w_000_635, w_003_038);
  and2 I005_275(w_005_275, w_000_264, w_002_438);
  not1 I005_276(w_005_276, w_001_666);
  or2  I005_277(w_005_277, w_000_737, w_003_155);
  and2 I005_278(w_005_278, w_000_325, w_004_011);
  or2  I005_280(w_005_280, w_001_778, w_002_334);
  not1 I005_281(w_005_281, w_001_222);
  not1 I005_282(w_005_282, w_003_160);
  not1 I005_283(w_005_283, w_004_001);
  and2 I005_284(w_005_284, w_002_182, w_000_639);
  and2 I005_285(w_005_285, w_004_033, w_002_072);
  nand2 I005_286(w_005_286, w_001_598, w_002_369);
  not1 I005_287(w_005_287, w_004_021);
  not1 I005_288(w_005_288, w_003_101);
  not1 I005_289(w_005_289, w_004_006);
  nand2 I005_291(w_005_291, w_001_163, w_000_633);
  and2 I005_292(w_005_292, w_000_426, w_003_072);
  nand2 I005_293(w_005_293, w_003_158, w_004_018);
  not1 I005_294(w_005_294, w_001_279);
  and2 I005_295(w_005_295, w_001_445, w_001_476);
  and2 I005_296(w_005_296, w_000_614, w_004_011);
  or2  I005_297(w_005_297, w_000_429, w_001_527);
  or2  I005_298(w_005_298, w_003_060, w_003_140);
  not1 I005_299(w_005_299, w_001_147);
  not1 I005_300(w_005_300, w_001_883);
  or2  I005_302(w_005_302, w_000_849, w_001_343);
  or2  I005_303(w_005_303, w_000_787, w_002_451);
  nand2 I005_304(w_005_304, w_000_504, w_004_016);
  and2 I005_305(w_005_305, w_003_126, w_001_270);
  not1 I005_306(w_005_306, w_004_015);
  and2 I005_307(w_005_307, w_003_021, w_000_386);
  or2  I005_308(w_005_308, w_001_011, w_001_854);
  or2  I005_309(w_005_309, w_004_002, w_002_279);
  and2 I005_310(w_005_310, w_001_083, w_002_418);
  nand2 I005_311(w_005_311, w_003_128, w_002_278);
  and2 I005_313(w_005_313, w_003_118, w_001_865);
  and2 I005_314(w_005_314, w_004_002, w_001_202);
  nand2 I005_315(w_005_315, w_001_099, w_001_785);
  and2 I005_316(w_005_316, w_002_271, w_001_700);
  and2 I005_317(w_005_317, w_002_070, w_000_174);
  nand2 I005_319(w_005_319, w_001_666, w_001_569);
  nand2 I005_320(w_005_320, w_004_009, w_004_007);
  or2  I005_322(w_005_322, w_001_221, w_002_376);
  or2  I005_323(w_005_323, w_002_379, w_003_014);
  nand2 I005_324(w_005_324, w_002_001, w_003_110);
  and2 I005_325(w_005_325, w_001_097, w_001_112);
  nand2 I005_327(w_005_327, w_000_177, w_000_893);
  not1 I005_328(w_005_328, w_001_082);
  nand2 I005_329(w_005_329, w_004_021, w_004_003);
  not1 I005_330(w_005_330, w_002_126);
  or2  I005_331(w_005_331, w_002_475, w_002_212);
  and2 I005_333(w_005_333, w_002_226, w_003_007);
  or2  I005_334(w_005_334, w_003_185, w_003_201);
  nand2 I005_335(w_005_335, w_001_314, w_002_370);
  nand2 I005_336(w_005_336, w_001_804, w_004_028);
  not1 I005_337(w_005_337, w_003_067);
  or2  I005_338(w_005_338, w_003_100, w_002_448);
  nand2 I005_339(w_005_339, w_000_381, w_004_003);
  not1 I005_342(w_005_342, w_001_893);
  nand2 I005_344(w_005_344, w_001_491, w_001_349);
  not1 I005_346(w_005_346, w_003_112);
  or2  I005_347(w_005_347, w_002_233, w_001_697);
  or2  I005_349(w_005_349, w_000_164, w_002_198);
  not1 I005_350(w_005_350, w_002_247);
  and2 I005_351(w_005_351, w_001_725, w_001_107);
  or2  I005_352(w_005_352, w_002_231, w_004_025);
  or2  I005_353(w_005_353, w_004_024, w_002_296);
  and2 I005_354(w_005_354, w_002_027, w_003_033);
  or2  I005_355(w_005_355, w_002_387, w_000_688);
  not1 I005_356(w_005_356, w_000_384);
  and2 I005_357(w_005_357, w_002_129, w_000_400);
  not1 I005_358(w_005_358, w_004_000);
  and2 I005_359(w_005_359, w_001_236, w_001_148);
  not1 I005_360(w_005_360, w_002_251);
  nand2 I005_361(w_005_361, w_003_195, w_003_174);
  or2  I005_362(w_005_362, w_000_214, w_002_042);
  and2 I005_363(w_005_363, w_002_444, w_001_518);
  and2 I005_364(w_005_364, w_000_000, w_002_260);
  not1 I005_365(w_005_365, w_001_768);
  not1 I005_366(w_005_366, w_004_005);
  and2 I005_367(w_005_367, w_003_130, w_004_011);
  not1 I005_368(w_005_368, w_002_338);
  nand2 I005_369(w_005_369, w_000_843, w_001_046);
  nand2 I005_371(w_005_371, w_003_180, w_001_238);
  nand2 I005_373(w_005_373, w_001_260, w_004_024);
  nand2 I005_374(w_005_374, w_000_674, w_002_291);
  and2 I005_375(w_005_375, w_001_269, w_000_685);
  nand2 I005_376(w_005_376, w_003_092, w_000_513);
  nand2 I005_377(w_005_377, w_001_103, w_001_032);
  not1 I005_378(w_005_378, w_000_168);
  nand2 I005_379(w_005_379, w_002_072, w_003_064);
  or2  I005_380(w_005_380, w_004_008, w_001_636);
  not1 I005_381(w_005_381, w_003_200);
  not1 I005_382(w_005_382, w_001_695);
  nand2 I005_384(w_005_384, w_002_415, w_000_895);
  not1 I005_385(w_005_385, w_000_017);
  not1 I005_386(w_005_386, w_004_004);
  nand2 I005_387(w_005_387, w_000_762, w_001_459);
  not1 I005_388(w_005_388, w_004_034);
  and2 I005_390(w_005_390, w_000_448, w_001_247);
  nand2 I005_391(w_005_391, w_000_085, w_003_189);
  and2 I005_392(w_005_392, w_003_141, w_001_000);
  nand2 I005_394(w_005_394, w_000_476, w_003_224);
  not1 I005_395(w_005_395, w_003_187);
  and2 I005_396(w_005_396, w_000_435, w_001_881);
  nand2 I005_397(w_005_397, w_000_480, w_001_155);
  not1 I005_399(w_005_399, w_000_896);
  or2  I005_400(w_005_400, w_004_020, w_001_032);
  or2  I005_401(w_005_401, w_003_182, w_003_035);
  nand2 I005_402(w_005_402, w_003_126, w_003_132);
  and2 I005_403(w_005_403, w_000_239, w_000_367);
  nand2 I005_404(w_005_404, w_001_522, w_002_048);
  or2  I005_405(w_005_405, w_001_465, w_004_025);
  or2  I005_407(w_005_407, w_001_174, w_003_085);
  or2  I005_408(w_005_408, w_002_234, w_003_160);
  or2  I005_409(w_005_409, w_000_604, w_004_022);
  nand2 I005_410(w_005_410, w_001_144, w_001_893);
  and2 I005_411(w_005_411, w_003_067, w_004_032);
  or2  I005_412(w_005_412, w_003_053, w_003_064);
  and2 I005_413(w_005_413, w_001_057, w_001_654);
  or2  I005_414(w_005_414, w_004_007, w_000_774);
  nand2 I005_415(w_005_415, w_000_084, w_000_629);
  not1 I005_416(w_005_416, w_001_885);
  not1 I005_417(w_005_417, w_002_130);
  not1 I005_418(w_005_418, w_003_002);
  nand2 I005_419(w_005_419, w_002_201, w_001_237);
  not1 I005_420(w_005_420, w_002_056);
  not1 I005_421(w_005_421, w_003_045);
  and2 I005_422(w_005_422, w_003_001, w_000_025);
  and2 I005_423(w_005_423, w_002_470, w_004_031);
  and2 I005_424(w_005_424, w_001_086, w_002_304);
  nand2 I005_425(w_005_425, w_003_014, w_000_897);
  nand2 I005_427(w_005_427, w_000_608, w_004_007);
  or2  I005_428(w_005_428, w_001_688, w_004_001);
  not1 I005_429(w_005_429, w_004_005);
  nand2 I005_431(w_005_431, w_004_005, w_001_794);
  or2  I005_433(w_005_433, w_000_823, w_002_462);
  and2 I005_436(w_005_436, w_004_027, w_001_094);
  not1 I005_440(w_005_440, w_000_072);
  not1 I005_441(w_005_441, w_004_011);
  and2 I005_443(w_005_443, w_000_294, w_001_047);
  nand2 I005_444(w_005_444, w_003_029, w_003_174);
  and2 I005_445(w_005_445, w_001_229, w_002_024);
  not1 I005_446(w_005_446, w_002_081);
  not1 I005_448(w_005_448, w_004_006);
  or2  I005_449(w_005_449, w_002_317, w_002_431);
  nand2 I005_450(w_005_450, w_004_038, w_003_072);
  nand2 I005_452(w_005_452, w_000_091, w_004_002);
  or2  I005_453(w_005_453, w_002_138, w_000_146);
  not1 I005_454(w_005_454, w_001_843);
  and2 I005_455(w_005_455, w_002_092, w_003_172);
  or2  I005_456(w_005_456, w_002_135, w_002_491);
  or2  I005_459(w_005_459, w_000_872, w_001_073);
  and2 I005_460(w_005_460, w_000_191, w_001_690);
  or2  I005_461(w_005_461, w_002_000, w_004_011);
  and2 I005_462(w_005_462, w_004_030, w_004_027);
  and2 I005_463(w_005_463, w_001_129, w_003_023);
  and2 I005_465(w_005_465, w_000_828, w_002_420);
  or2  I005_466(w_005_466, w_004_003, w_002_432);
  or2  I005_467(w_005_467, w_003_005, w_003_056);
  and2 I005_470(w_005_470, w_002_064, w_001_249);
  and2 I005_471(w_005_471, w_001_672, w_003_183);
  not1 I005_472(w_005_472, w_004_001);
  or2  I005_473(w_005_473, w_004_009, w_002_406);
  or2  I005_474(w_005_474, w_002_140, w_004_037);
  not1 I005_476(w_005_476, w_000_873);
  not1 I005_477(w_005_477, w_004_007);
  or2  I005_478(w_005_478, w_001_196, w_001_066);
  nand2 I005_480(w_005_480, w_001_598, w_000_815);
  or2  I005_482(w_005_482, w_004_026, w_001_893);
  and2 I005_483(w_005_483, w_001_767, w_001_006);
  or2  I005_485(w_005_485, w_004_030, w_001_216);
  not1 I005_486(w_005_486, w_004_012);
  not1 I005_490(w_005_490, w_003_185);
  or2  I005_493(w_005_493, w_002_431, w_004_007);
  and2 I005_495(w_005_495, w_004_014, w_001_288);
  and2 I005_496(w_005_496, w_003_217, w_004_011);
  or2  I005_497(w_005_497, w_004_033, w_003_200);
  or2  I005_499(w_005_499, w_002_340, w_004_002);
  or2  I005_502(w_005_502, w_000_852, w_000_761);
  nand2 I005_503(w_005_503, w_004_026, w_004_038);
  and2 I005_509(w_005_509, w_003_115, w_002_494);
  nand2 I005_511(w_005_511, w_001_432, w_000_844);
  or2  I005_512(w_005_512, w_001_762, w_004_031);
  or2  I005_515(w_005_515, w_000_782, w_002_340);
  and2 I005_516(w_005_516, w_004_021, w_004_027);
  and2 I005_517(w_005_517, w_001_388, w_004_038);
  and2 I005_518(w_005_518, w_000_065, w_001_001);
  or2  I005_521(w_005_521, w_004_019, w_002_486);
  and2 I005_524(w_005_524, w_004_011, w_001_031);
  or2  I005_525(w_005_525, w_002_033, w_001_205);
  nand2 I005_526(w_005_526, w_002_383, w_000_526);
  nand2 I005_531(w_005_531, w_004_034, w_003_095);
  and2 I005_532(w_005_532, w_001_480, w_002_325);
  not1 I005_537(w_005_537, w_004_008);
  or2  I005_539(w_005_539, w_002_088, w_003_099);
  or2  I005_542(w_005_542, w_004_028, w_004_026);
  not1 I005_544(w_005_544, w_004_036);
  not1 I005_545(w_005_545, w_002_423);
  and2 I005_547(w_005_547, w_004_010, w_001_606);
  not1 I005_548(w_005_548, w_001_757);
  or2  I005_549(w_005_549, w_000_166, w_000_859);
  nand2 I005_551(w_005_551, w_000_773, w_001_822);
  not1 I005_556(w_005_556, w_001_710);
  not1 I005_559(w_005_559, w_000_028);
  or2  I005_560(w_005_560, w_001_763, w_001_843);
  not1 I005_561(w_005_561, w_000_878);
  and2 I005_564(w_005_564, w_001_191, w_004_036);
  and2 I005_565(w_005_565, w_002_265, w_003_153);
  or2  I005_569(w_005_569, w_002_013, w_002_269);
  not1 I005_570(w_005_570, w_004_008);
  nand2 I005_574(w_005_574, w_000_272, w_001_479);
  nand2 I006_000(w_006_000, w_000_255, w_001_519);
  and2 I006_002(w_006_002, w_004_035, w_002_459);
  not1 I006_003(w_006_003, w_002_233);
  not1 I006_004(w_006_004, w_002_333);
  nand2 I006_005(w_006_005, w_005_329, w_003_172);
  nand2 I006_007(w_006_007, w_001_882, w_002_370);
  not1 I006_008(w_006_008, w_001_100);
  not1 I006_009(w_006_009, w_003_185);
  not1 I006_010(w_006_010, w_004_030);
  or2  I006_011(w_006_011, w_004_024, w_004_013);
  and2 I006_012(w_006_012, w_001_225, w_003_196);
  and2 I006_013(w_006_013, w_003_140, w_002_265);
  and2 I006_014(w_006_014, w_001_452, w_003_077);
  and2 I006_015(w_006_015, w_004_007, w_003_035);
  not1 I006_016(w_006_016, w_005_220);
  and2 I006_017(w_006_017, w_003_041, w_003_095);
  nand2 I006_018(w_006_018, w_002_185, w_001_533);
  not1 I006_020(w_006_020, w_005_565);
  not1 I006_021(w_006_021, w_004_018);
  and2 I006_022(w_006_022, w_001_293, w_002_297);
  or2  I006_023(w_006_023, w_003_139, w_004_036);
  nand2 I006_024(w_006_024, w_001_380, w_005_351);
  and2 I006_025(w_006_025, w_001_609, w_005_264);
  or2  I006_026(w_006_026, w_002_496, w_004_015);
  or2  I006_027(w_006_027, w_001_283, w_005_200);
  and2 I006_028(w_006_028, w_003_045, w_001_881);
  not1 I006_029(w_006_029, w_000_618);
  not1 I006_030(w_006_030, w_004_006);
  or2  I006_031(w_006_031, w_003_208, w_002_173);
  or2  I006_034(w_006_034, w_002_268, w_001_205);
  not1 I006_035(w_006_035, w_002_008);
  and2 I006_036(w_006_036, w_000_105, w_002_286);
  and2 I006_038(w_006_038, w_001_574, w_000_400);
  and2 I006_039(w_006_039, w_003_070, w_004_029);
  nand2 I006_040(w_006_040, w_005_448, w_002_341);
  nand2 I006_041(w_006_041, w_001_001, w_003_170);
  or2  I006_042(w_006_042, w_005_409, w_002_464);
  and2 I006_043(w_006_043, w_001_617, w_002_171);
  or2  I006_044(w_006_044, w_004_034, w_005_056);
  or2  I006_045(w_006_045, w_000_256, w_001_716);
  or2  I006_046(w_006_046, w_002_129, w_001_515);
  not1 I006_048(w_006_048, w_004_035);
  nand2 I006_050(w_006_050, w_005_116, w_003_212);
  not1 I006_051(w_006_051, w_000_777);
  or2  I006_052(w_006_052, w_002_290, w_005_136);
  or2  I006_053(w_006_053, w_000_357, w_004_013);
  nand2 I006_054(w_006_054, w_001_802, w_003_201);
  or2  I006_055(w_006_055, w_001_350, w_001_088);
  and2 I006_056(w_006_056, w_005_261, w_005_126);
  or2  I006_057(w_006_057, w_001_790, w_003_149);
  nand2 I006_058(w_006_058, w_004_021, w_001_006);
  and2 I006_059(w_006_059, w_003_056, w_005_499);
  or2  I006_060(w_006_060, w_002_174, w_005_281);
  or2  I006_061(w_006_061, w_002_307, w_005_161);
  not1 I006_062(w_006_062, w_004_020);
  nand2 I006_063(w_006_063, w_001_122, w_004_038);
  or2  I006_064(w_006_064, w_001_233, w_002_003);
  or2  I006_065(w_006_065, w_002_357, w_003_085);
  or2  I006_066(w_006_066, w_002_086, w_003_167);
  not1 I006_067(w_006_067, w_002_023);
  nand2 I006_068(w_006_068, w_003_180, w_003_224);
  nand2 I006_069(w_006_069, w_005_098, w_002_496);
  not1 I006_071(w_006_071, w_001_772);
  nand2 I006_073(w_006_073, w_001_716, w_004_037);
  not1 I006_074(w_006_074, w_005_110);
  or2  I006_075(w_006_075, w_002_367, w_002_448);
  and2 I006_076(w_006_076, w_005_121, w_000_754);
  or2  I006_078(w_006_078, w_000_438, w_001_325);
  and2 I006_079(w_006_079, w_001_457, w_003_050);
  or2  I006_080(w_006_080, w_002_440, w_005_431);
  nand2 I006_082(w_006_082, w_003_199, w_001_632);
  not1 I006_084(w_006_084, w_003_028);
  and2 I006_085(w_006_085, w_002_031, w_004_018);
  or2  I006_086(w_006_086, w_001_021, w_000_749);
  or2  I006_087(w_006_087, w_004_025, w_004_017);
  nand2 I006_088(w_006_088, w_001_088, w_003_181);
  or2  I006_089(w_006_089, w_004_001, w_000_554);
  nand2 I006_090(w_006_090, w_004_004, w_001_718);
  nand2 I006_091(w_006_091, w_001_226, w_005_449);
  nand2 I006_094(w_006_094, w_002_067, w_000_854);
  and2 I006_095(w_006_095, w_003_035, w_001_293);
  and2 I006_096(w_006_096, w_000_847, w_005_377);
  or2  I006_097(w_006_097, w_001_022, w_004_006);
  or2  I006_098(w_006_098, w_003_206, w_005_164);
  or2  I006_099(w_006_099, w_000_666, w_003_082);
  not1 I006_100(w_006_100, w_000_489);
  not1 I006_101(w_006_101, w_001_343);
  not1 I006_102(w_006_102, w_002_458);
  nand2 I006_103(w_006_103, w_002_312, w_005_336);
  nand2 I006_104(w_006_104, w_004_037, w_002_004);
  or2  I006_105(w_006_105, w_003_153, w_004_019);
  nand2 I006_106(w_006_106, w_000_903, w_005_490);
  nand2 I006_107(w_006_107, w_004_035, w_002_391);
  not1 I006_108(w_006_108, w_003_132);
  and2 I006_109(w_006_109, w_003_088, w_000_297);
  and2 I006_110(w_006_110, w_003_109, w_005_391);
  or2  I006_111(w_006_111, w_002_396, w_000_267);
  or2  I006_112(w_006_112, w_005_179, w_000_411);
  not1 I006_113(w_006_113, w_000_901);
  or2  I006_114(w_006_114, w_002_053, w_005_234);
  and2 I006_115(w_006_115, w_000_393, w_004_023);
  or2  I006_116(w_006_116, w_002_251, w_003_028);
  not1 I006_117(w_006_117, w_002_147);
  and2 I006_118(w_006_118, w_004_002, w_000_107);
  nand2 I006_119(w_006_119, w_003_213, w_003_012);
  nand2 I006_120(w_006_120, w_001_365, w_001_319);
  nand2 I006_121(w_006_121, w_000_128, w_001_871);
  or2  I006_122(w_006_122, w_005_323, w_004_016);
  and2 I006_123(w_006_123, w_001_270, w_003_076);
  nand2 I006_124(w_006_124, w_003_142, w_003_065);
  and2 I006_125(w_006_125, w_004_026, w_003_131);
  nand2 I006_126(w_006_126, w_001_631, w_005_358);
  not1 I006_127(w_006_127, w_000_010);
  nand2 I006_128(w_006_128, w_001_233, w_002_312);
  and2 I006_129(w_006_129, w_005_251, w_005_295);
  and2 I006_130(w_006_130, w_000_850, w_000_823);
  nand2 I006_131(w_006_131, w_003_014, w_005_081);
  nand2 I006_132(w_006_132, w_002_166, w_001_313);
  nand2 I006_133(w_006_133, w_004_023, w_000_336);
  nand2 I006_135(w_006_135, w_005_210, w_002_410);
  and2 I006_136(w_006_136, w_005_131, w_002_487);
  or2  I006_137(w_006_137, w_002_160, w_000_505);
  and2 I006_138(w_006_138, w_003_034, w_000_512);
  nand2 I006_139(w_006_139, w_005_177, w_002_489);
  or2  I006_140(w_006_140, w_002_323, w_003_059);
  not1 I006_141(w_006_141, w_000_027);
  nand2 I006_142(w_006_142, w_000_287, w_005_299);
  not1 I006_143(w_006_143, w_002_138);
  and2 I006_144(w_006_144, w_004_016, w_004_035);
  or2  I006_145(w_006_145, w_002_294, w_003_080);
  not1 I006_147(w_006_147, w_004_011);
  or2  I006_148(w_006_148, w_002_012, w_002_125);
  nand2 I006_149(w_006_149, w_002_262, w_003_216);
  or2  I006_150(w_006_150, w_003_078, w_005_063);
  or2  I006_153(w_006_153, w_003_059, w_003_196);
  or2  I006_154(w_006_154, w_002_010, w_005_195);
  not1 I006_155(w_006_155, w_001_745);
  or2  I006_156(w_006_156, w_001_007, w_000_875);
  and2 I006_157(w_006_157, w_003_180, w_005_280);
  or2  I006_158(w_006_158, w_003_124, w_005_436);
  not1 I006_159(w_006_159, w_000_786);
  and2 I006_160(w_006_160, w_003_071, w_001_635);
  not1 I006_161(w_006_161, w_001_100);
  or2  I006_162(w_006_162, w_003_145, w_000_364);
  and2 I006_163(w_006_163, w_002_226, w_003_137);
  and2 I006_164(w_006_164, w_000_904, w_002_417);
  and2 I006_165(w_006_165, w_003_166, w_005_226);
  not1 I006_166(w_006_166, w_005_012);
  not1 I006_167(w_006_167, w_002_236);
  not1 I006_168(w_006_168, w_003_081);
  nand2 I006_169(w_006_169, w_002_310, w_003_225);
  or2  I006_170(w_006_170, w_001_222, w_003_215);
  nand2 I006_171(w_006_171, w_002_482, w_001_192);
  not1 I006_172(w_006_172, w_001_328);
  nand2 I006_173(w_006_173, w_005_359, w_000_845);
  or2  I006_174(w_006_174, w_002_034, w_004_032);
  not1 I006_175(w_006_175, w_001_727);
  or2  I006_176(w_006_176, w_002_038, w_004_026);
  or2  I006_177(w_006_177, w_004_029, w_002_179);
  not1 I006_178(w_006_178, w_004_004);
  not1 I006_179(w_006_179, w_000_137);
  or2  I006_180(w_006_180, w_005_201, w_004_001);
  or2  I006_181(w_006_181, w_001_308, w_001_613);
  and2 I006_182(w_006_182, w_001_155, w_004_037);
  or2  I006_183(w_006_183, w_004_003, w_005_135);
  not1 I006_184(w_006_184, w_003_017);
  not1 I006_185(w_006_185, w_005_193);
  not1 I006_186(w_006_186, w_000_047);
  nand2 I006_187(w_006_187, w_004_018, w_002_156);
  and2 I006_188(w_006_188, w_003_023, w_004_002);
  and2 I006_189(w_006_189, w_005_249, w_000_511);
  and2 I006_191(w_006_191, w_000_745, w_005_158);
  nand2 I006_192(w_006_192, w_002_418, w_004_020);
  not1 I006_193(w_006_193, w_002_199);
  and2 I006_195(w_006_195, w_000_520, w_004_025);
  or2  I006_196(w_006_196, w_004_005, w_003_189);
  not1 I006_197(w_006_197, w_000_257);
  not1 I006_198(w_006_198, w_004_003);
  and2 I006_201(w_006_201, w_002_411, w_001_005);
  and2 I006_202(w_006_202, w_000_878, w_004_031);
  nand2 I006_203(w_006_203, w_000_090, w_004_010);
  or2  I006_205(w_006_205, w_001_098, w_002_377);
  not1 I006_206(w_006_206, w_004_011);
  and2 I006_207(w_006_207, w_002_161, w_000_905);
  not1 I006_208(w_006_208, w_000_906);
  not1 I006_209(w_006_209, w_000_830);
  or2  I006_210(w_006_210, w_004_005, w_001_056);
  nand2 I006_211(w_006_211, w_001_440, w_001_637);
  not1 I006_212(w_006_212, w_001_078);
  or2  I006_213(w_006_213, w_005_094, w_005_197);
  or2  I006_214(w_006_214, w_000_801, w_005_208);
  not1 I006_215(w_006_215, w_005_206);
  and2 I006_216(w_006_216, w_003_068, w_004_016);
  nand2 I006_218(w_006_218, w_004_038, w_002_259);
  nand2 I006_220(w_006_220, w_002_335, w_004_001);
  or2  I006_221(w_006_221, w_001_486, w_001_448);
  and2 I006_222(w_006_222, w_005_258, w_003_137);
  or2  I006_223(w_006_223, w_000_161, w_000_141);
  nand2 I006_224(w_006_224, w_005_188, w_005_413);
  nand2 I006_225(w_006_225, w_005_151, w_003_014);
  not1 I006_226(w_006_226, w_004_029);
  or2  I006_227(w_006_227, w_000_200, w_002_253);
  not1 I006_228(w_006_228, w_001_551);
  nand2 I006_229(w_006_229, w_000_161, w_000_667);
  nand2 I006_230(w_006_230, w_000_180, w_005_089);
  nand2 I006_231(w_006_231, w_004_037, w_002_412);
  not1 I006_232(w_006_232, w_005_062);
  nand2 I006_233(w_006_233, w_000_704, w_001_677);
  or2  I006_234(w_006_234, w_005_229, w_002_352);
  nand2 I006_235(w_006_235, w_003_076, w_000_122);
  nand2 I006_236(w_006_236, w_000_141, w_004_014);
  not1 I006_237(w_006_237, w_003_115);
  or2  I006_238(w_006_238, w_002_120, w_000_676);
  nand2 I006_239(w_006_239, w_003_090, w_002_325);
  not1 I006_240(w_006_240, w_002_354);
  and2 I006_241(w_006_241, w_001_081, w_000_384);
  or2  I006_242(w_006_242, w_003_138, w_005_071);
  or2  I006_243(w_006_243, w_004_018, w_002_089);
  nand2 I006_244(w_006_244, w_005_353, w_000_693);
  and2 I006_245(w_006_245, w_000_722, w_003_160);
  and2 I006_246(w_006_246, w_000_561, w_003_096);
  not1 I006_247(w_006_247, w_001_729);
  nand2 I006_248(w_006_248, w_005_113, w_004_003);
  nand2 I006_249(w_006_249, w_002_192, w_001_214);
  or2  I006_250(w_006_250, w_003_123, w_002_170);
  or2  I006_251(w_006_251, w_002_216, w_003_069);
  and2 I006_252(w_006_252, w_001_485, w_004_037);
  not1 I006_253(w_006_253, w_001_819);
  and2 I006_254(w_006_254, w_000_548, w_004_026);
  not1 I006_255(w_006_255, w_002_342);
  or2  I006_256(w_006_256, w_004_028, w_004_000);
  nand2 I006_257(w_006_257, w_005_304, w_001_036);
  and2 I006_258(w_006_258, w_001_750, w_000_038);
  not1 I006_259(w_006_259, w_001_523);
  not1 I006_260(w_006_260, w_004_024);
  not1 I006_261(w_006_261, w_003_156);
  and2 I006_262(w_006_262, w_001_042, w_002_307);
  nand2 I006_263(w_006_263, w_000_907, w_001_606);
  nand2 I006_264(w_006_264, w_004_000, w_005_425);
  and2 I006_265(w_006_265, w_003_060, w_001_353);
  and2 I006_266(w_006_266, w_002_243, w_003_037);
  or2  I006_267(w_006_267, w_001_607, w_003_098);
  not1 I006_268(w_006_268, w_002_391);
  and2 I006_270(w_006_270, w_003_066, w_003_071);
  or2  I006_271(w_006_271, w_002_074, w_001_697);
  and2 I006_272(w_006_272, w_002_402, w_002_216);
  or2  I006_273(w_006_273, w_003_104, w_001_236);
  nand2 I006_274(w_006_274, w_004_022, w_003_002);
  not1 I006_275(w_006_275, w_002_420);
  or2  I006_276(w_006_276, w_003_106, w_003_076);
  not1 I006_277(w_006_277, w_004_021);
  nand2 I006_278(w_006_278, w_005_252, w_004_018);
  and2 I006_279(w_006_279, w_001_123, w_005_060);
  and2 I006_280(w_006_280, w_002_091, w_001_177);
  nand2 I006_281(w_006_281, w_000_863, w_000_524);
  or2  I006_282(w_006_282, w_000_297, w_004_034);
  nand2 I006_283(w_006_283, w_005_377, w_002_400);
  not1 I006_284(w_006_284, w_005_423);
  not1 I006_285(w_006_285, w_004_027);
  not1 I006_286(w_006_286, w_003_066);
  nand2 I006_287(w_006_287, w_004_013, w_000_518);
  not1 I006_288(w_006_288, w_003_221);
  and2 I006_289(w_006_289, w_004_038, w_003_186);
  and2 I006_290(w_006_290, w_000_256, w_000_293);
  and2 I006_291(w_006_291, w_002_151, w_002_442);
  or2  I006_292(w_006_292, w_003_176, w_005_175);
  nand2 I006_293(w_006_293, w_000_721, w_000_036);
  and2 I006_294(w_006_294, w_000_554, w_004_002);
  nand2 I006_295(w_006_295, w_003_038, w_005_416);
  not1 I006_296(w_006_296, w_003_050);
  not1 I006_297(w_006_297, w_001_599);
  not1 I006_298(w_006_298, w_003_073);
  not1 I006_299(w_006_299, w_002_052);
  or2  I006_300(w_006_300, w_002_223, w_004_017);
  and2 I006_302(w_006_302, w_004_008, w_004_005);
  not1 I006_303(w_006_303, w_004_014);
  not1 I006_304(w_006_304, w_004_036);
  and2 I006_305(w_006_305, w_000_378, w_002_093);
  and2 I006_306(w_006_306, w_001_013, w_000_183);
  nand2 I006_307(w_006_307, w_000_758, w_003_128);
  nand2 I006_308(w_006_308, w_000_086, w_000_908);
  not1 I006_309(w_006_309, w_004_036);
  not1 I006_310(w_006_310, w_000_171);
  not1 I006_311(w_006_311, w_004_020);
  and2 I006_312(w_006_312, w_004_020, w_005_001);
  not1 I006_313(w_006_313, w_004_026);
  or2  I006_314(w_006_314, w_003_066, w_000_028);
  or2  I006_315(w_006_315, w_004_031, w_005_117);
  nand2 I006_316(w_006_316, w_005_281, w_000_501);
  not1 I006_317(w_006_317, w_005_156);
  not1 I006_318(w_006_318, w_002_196);
  not1 I006_319(w_006_319, w_001_723);
  and2 I006_320(w_006_320, w_005_177, w_001_269);
  and2 I006_321(w_006_321, w_003_050, w_005_102);
  not1 I006_322(w_006_322, w_000_255);
  and2 I006_323(w_006_323, w_003_210, w_001_765);
  nand2 I006_324(w_006_324, w_001_577, w_002_417);
  not1 I006_325(w_006_325, w_004_031);
  not1 I006_326(w_006_326, w_001_845);
  and2 I006_327(w_006_327, w_002_400, w_001_138);
  nand2 I006_328(w_006_328, w_003_114, w_002_447);
  nand2 I006_329(w_006_329, w_004_014, w_003_041);
  not1 I006_330(w_006_330, w_005_258);
  and2 I006_331(w_006_331, w_002_294, w_005_465);
  or2  I006_332(w_006_332, w_002_174, w_005_271);
  and2 I007_000(w_007_000, w_001_834, w_001_366);
  not1 I007_001(w_007_001, w_003_215);
  nand2 I007_002(w_007_002, w_006_130, w_005_306);
  not1 I007_004(w_007_004, w_000_043);
  not1 I007_005(w_007_005, w_003_102);
  or2  I007_007(w_007_007, w_001_103, w_002_299);
  and2 I007_010(w_007_010, w_000_136, w_003_168);
  not1 I007_011(w_007_011, w_002_254);
  or2  I007_012(w_007_012, w_001_547, w_006_239);
  nand2 I007_013(w_007_013, w_003_161, w_004_009);
  and2 I007_014(w_007_014, w_005_268, w_001_202);
  or2  I007_015(w_007_015, w_005_509, w_000_247);
  not1 I007_017(w_007_017, w_000_440);
  and2 I007_018(w_007_018, w_000_545, w_000_824);
  and2 I007_019(w_007_019, w_004_027, w_000_054);
  and2 I007_020(w_007_020, w_004_024, w_006_062);
  nand2 I007_021(w_007_021, w_005_375, w_001_791);
  and2 I007_023(w_007_023, w_001_678, w_002_390);
  nand2 I007_024(w_007_024, w_003_135, w_004_008);
  nand2 I007_026(w_007_026, w_001_053, w_001_046);
  and2 I007_027(w_007_027, w_000_775, w_002_483);
  and2 I007_029(w_007_029, w_005_394, w_006_054);
  and2 I007_030(w_007_030, w_001_063, w_000_499);
  or2  I007_031(w_007_031, w_002_283, w_005_299);
  not1 I007_032(w_007_032, w_001_010);
  or2  I007_033(w_007_033, w_002_063, w_005_329);
  not1 I007_035(w_007_035, w_001_403);
  nand2 I007_038(w_007_038, w_001_582, w_006_288);
  and2 I007_039(w_007_039, w_000_162, w_005_120);
  nand2 I007_040(w_007_040, w_005_110, w_002_030);
  not1 I007_041(w_007_041, w_005_061);
  and2 I007_042(w_007_042, w_005_011, w_000_618);
  not1 I007_043(w_007_043, w_006_029);
  or2  I007_044(w_007_044, w_002_419, w_005_388);
  nand2 I007_045(w_007_045, w_004_000, w_002_206);
  or2  I007_046(w_007_046, w_001_866, w_002_438);
  or2  I007_047(w_007_047, w_000_549, w_003_113);
  nand2 I007_048(w_007_048, w_006_193, w_006_162);
  not1 I007_049(w_007_049, w_006_133);
  and2 I007_050(w_007_050, w_003_168, w_003_116);
  not1 I007_052(w_007_052, w_000_738);
  nand2 I007_053(w_007_053, w_006_290, w_001_119);
  or2  I007_054(w_007_054, w_006_002, w_002_200);
  nand2 I007_055(w_007_055, w_006_060, w_001_714);
  nand2 I007_057(w_007_057, w_004_016, w_002_216);
  and2 I007_058(w_007_058, w_000_251, w_005_276);
  nand2 I007_060(w_007_060, w_006_244, w_005_224);
  nand2 I007_062(w_007_062, w_000_439, w_000_676);
  or2  I007_063(w_007_063, w_006_256, w_001_728);
  not1 I007_064(w_007_064, w_003_189);
  or2  I007_065(w_007_065, w_001_492, w_006_064);
  nand2 I007_067(w_007_067, w_001_612, w_003_027);
  not1 I007_068(w_007_068, w_000_713);
  or2  I007_069(w_007_069, w_001_152, w_001_046);
  or2  I007_070(w_007_070, w_005_320, w_003_035);
  and2 I007_072(w_007_072, w_005_271, w_001_195);
  not1 I007_073(w_007_073, w_000_454);
  not1 I007_074(w_007_074, w_003_053);
  or2  I007_075(w_007_075, w_005_033, w_000_499);
  nand2 I007_076(w_007_076, w_004_005, w_002_160);
  not1 I007_077(w_007_077, w_004_019);
  and2 I007_078(w_007_078, w_002_273, w_000_385);
  and2 I007_079(w_007_079, w_004_016, w_000_882);
  and2 I007_080(w_007_080, w_002_311, w_005_405);
  nand2 I007_081(w_007_081, w_000_289, w_004_017);
  not1 I007_082(w_007_082, w_003_111);
  or2  I007_083(w_007_083, w_005_185, w_003_158);
  or2  I007_085(w_007_085, w_003_131, w_004_017);
  or2  I007_088(w_007_088, w_001_639, w_002_067);
  and2 I007_089(w_007_089, w_003_066, w_006_225);
  nand2 I007_091(w_007_091, w_004_016, w_001_032);
  and2 I007_092(w_007_092, w_003_057, w_006_171);
  and2 I007_093(w_007_093, w_004_031, w_001_009);
  and2 I007_094(w_007_094, w_004_005, w_006_053);
  nand2 I007_095(w_007_095, w_001_018, w_004_000);
  and2 I007_097(w_007_097, w_004_006, w_002_160);
  not1 I007_098(w_007_098, w_001_604);
  nand2 I007_099(w_007_099, w_006_128, w_004_002);
  nand2 I007_100(w_007_100, w_005_296, w_006_161);
  or2  I007_101(w_007_101, w_003_096, w_004_013);
  not1 I007_103(w_007_103, w_004_018);
  not1 I007_105(w_007_105, w_002_235);
  nand2 I007_107(w_007_107, w_003_163, w_004_009);
  not1 I007_108(w_007_108, w_005_038);
  or2  I007_109(w_007_109, w_002_108, w_006_302);
  and2 I007_110(w_007_110, w_002_363, w_002_447);
  or2  I007_111(w_007_111, w_000_803, w_001_002);
  nand2 I007_113(w_007_113, w_002_068, w_002_465);
  nand2 I007_115(w_007_115, w_003_210, w_002_386);
  and2 I007_116(w_007_116, w_000_175, w_000_769);
  not1 I007_117(w_007_117, w_002_190);
  not1 I007_119(w_007_119, w_006_030);
  or2  I007_121(w_007_121, w_002_386, w_000_881);
  or2  I007_122(w_007_122, w_002_046, w_006_079);
  and2 I007_123(w_007_123, w_004_020, w_006_266);
  not1 I007_127(w_007_127, w_001_663);
  nand2 I007_128(w_007_128, w_004_010, w_004_025);
  nand2 I007_129(w_007_129, w_004_037, w_000_855);
  and2 I007_130(w_007_130, w_002_461, w_003_000);
  or2  I007_131(w_007_131, w_000_682, w_003_089);
  nand2 I007_132(w_007_132, w_001_115, w_000_396);
  nand2 I007_134(w_007_134, w_000_789, w_006_184);
  or2  I007_135(w_007_135, w_000_312, w_004_012);
  nand2 I007_136(w_007_136, w_006_126, w_006_170);
  not1 I007_137(w_007_137, w_003_209);
  or2  I007_138(w_007_138, w_006_298, w_005_286);
  or2  I007_139(w_007_139, w_006_034, w_006_298);
  not1 I007_140(w_007_140, w_000_749);
  and2 I007_142(w_007_142, w_004_028, w_005_397);
  and2 I007_143(w_007_143, w_003_086, w_003_111);
  nand2 I007_144(w_007_144, w_006_320, w_004_024);
  not1 I007_145(w_007_145, w_002_443);
  nand2 I007_147(w_007_147, w_003_075, w_000_909);
  not1 I007_148(w_007_148, w_004_004);
  not1 I007_149(w_007_149, w_001_282);
  not1 I007_150(w_007_150, w_003_158);
  nand2 I007_151(w_007_151, w_005_344, w_006_119);
  and2 I007_152(w_007_152, w_003_207, w_005_050);
  nand2 I007_153(w_007_153, w_000_434, w_003_055);
  or2  I007_155(w_007_155, w_006_263, w_003_054);
  nand2 I007_156(w_007_156, w_004_007, w_001_826);
  not1 I007_157(w_007_157, w_003_006);
  or2  I007_158(w_007_158, w_002_079, w_005_396);
  and2 I007_159(w_007_159, w_003_220, w_003_113);
  and2 I007_160(w_007_160, w_004_017, w_004_012);
  or2  I007_161(w_007_161, w_001_130, w_002_021);
  and2 I007_162(w_007_162, w_005_331, w_000_353);
  nand2 I007_163(w_007_163, w_001_179, w_006_046);
  or2  I007_164(w_007_164, w_003_117, w_001_729);
  nand2 I007_165(w_007_165, w_001_616, w_004_005);
  nand2 I007_166(w_007_166, w_003_160, w_004_029);
  nand2 I007_167(w_007_167, w_000_682, w_004_017);
  nand2 I007_168(w_007_168, w_003_014, w_003_189);
  nand2 I007_169(w_007_169, w_003_136, w_004_022);
  not1 I007_171(w_007_171, w_003_115);
  or2  I007_173(w_007_173, w_002_161, w_002_288);
  nand2 I007_175(w_007_175, w_003_194, w_006_332);
  and2 I007_177(w_007_177, w_000_614, w_002_207);
  and2 I007_179(w_007_179, w_001_071, w_001_761);
  or2  I007_182(w_007_182, w_001_006, w_005_220);
  nand2 I007_183(w_007_183, w_004_014, w_006_237);
  or2  I007_185(w_007_185, w_000_230, w_000_089);
  or2  I007_186(w_007_186, w_001_203, w_004_032);
  not1 I007_187(w_007_187, w_000_489);
  and2 I007_188(w_007_188, w_006_290, w_004_035);
  and2 I007_189(w_007_189, w_003_031, w_002_460);
  not1 I007_190(w_007_190, w_004_008);
  not1 I007_192(w_007_192, w_001_678);
  nand2 I007_193(w_007_193, w_005_331, w_003_183);
  or2  I007_194(w_007_194, w_005_282, w_004_018);
  not1 I007_195(w_007_195, w_003_048);
  and2 I007_196(w_007_196, w_003_037, w_001_798);
  and2 I007_198(w_007_198, w_006_162, w_005_503);
  not1 I007_199(w_007_199, w_004_025);
  or2  I007_200(w_007_200, w_003_060, w_006_175);
  or2  I007_201(w_007_201, w_004_006, w_004_000);
  or2  I007_202(w_007_202, w_005_164, w_003_095);
  or2  I007_203(w_007_203, w_002_199, w_004_019);
  not1 I007_204(w_007_204, w_002_421);
  not1 I007_205(w_007_205, w_006_250);
  not1 I007_207(w_007_207, w_003_066);
  and2 I007_208(w_007_208, w_004_029, w_006_131);
  or2  I007_209(w_007_209, w_006_170, w_000_899);
  and2 I007_210(w_007_210, w_005_357, w_005_446);
  nand2 I007_212(w_007_212, w_004_012, w_006_255);
  and2 I007_213(w_007_213, w_004_006, w_005_096);
  or2  I007_214(w_007_214, w_006_012, w_006_016);
  not1 I007_215(w_007_215, w_001_084);
  or2  I007_216(w_007_216, w_002_336, w_002_392);
  or2  I007_217(w_007_217, w_000_190, w_004_027);
  nand2 I007_218(w_007_218, w_002_227, w_002_431);
  or2  I007_219(w_007_219, w_006_039, w_002_316);
  and2 I007_220(w_007_220, w_005_339, w_004_007);
  and2 I007_221(w_007_221, w_003_115, w_004_027);
  nand2 I007_222(w_007_222, w_003_194, w_001_634);
  not1 I007_223(w_007_223, w_000_594);
  and2 I007_224(w_007_224, w_004_012, w_001_627);
  or2  I007_228(w_007_228, w_005_445, w_005_288);
  nand2 I007_229(w_007_229, w_004_031, w_004_021);
  and2 I007_230(w_007_230, w_005_118, w_002_087);
  or2  I007_232(w_007_232, w_006_034, w_005_482);
  not1 I007_233(w_007_233, w_005_147);
  not1 I007_234(w_007_234, w_002_029);
  not1 I007_235(w_007_235, w_000_479);
  or2  I007_236(w_007_236, w_004_034, w_002_345);
  and2 I007_237(w_007_237, w_003_179, w_000_910);
  or2  I007_238(w_007_238, w_003_134, w_001_118);
  or2  I007_239(w_007_239, w_002_275, w_001_136);
  and2 I007_240(w_007_240, w_004_014, w_004_003);
  not1 I007_243(w_007_243, w_004_009);
  nand2 I007_244(w_007_244, w_000_578, w_005_521);
  nand2 I007_245(w_007_245, w_006_007, w_005_179);
  and2 I007_246(w_007_246, w_006_048, w_006_254);
  or2  I007_247(w_007_247, w_003_085, w_002_492);
  not1 I007_248(w_007_248, w_001_570);
  and2 I007_249(w_007_249, w_006_314, w_001_158);
  nand2 I007_250(w_007_250, w_005_334, w_001_182);
  nand2 I007_251(w_007_251, w_004_017, w_003_035);
  nand2 I007_252(w_007_252, w_002_045, w_006_163);
  nand2 I007_253(w_007_253, w_005_175, w_000_066);
  nand2 I007_254(w_007_254, w_003_182, w_004_034);
  not1 I007_255(w_007_255, w_002_193);
  nand2 I007_256(w_007_256, w_003_026, w_006_296);
  or2  I007_257(w_007_257, w_000_144, w_000_270);
  nand2 I007_259(w_007_259, w_006_024, w_002_125);
  and2 I007_260(w_007_260, w_002_045, w_002_435);
  and2 I007_261(w_007_261, w_006_004, w_005_007);
  nand2 I007_262(w_007_262, w_006_040, w_006_227);
  not1 I007_264(w_007_264, w_006_191);
  nand2 I007_265(w_007_265, w_006_071, w_000_852);
  nand2 I007_266(w_007_266, w_000_330, w_004_033);
  or2  I007_267(w_007_267, w_006_198, w_004_029);
  not1 I007_268(w_007_268, w_001_857);
  not1 I007_269(w_007_269, w_005_230);
  not1 I007_272(w_007_272, w_002_378);
  nand2 I007_273(w_007_273, w_005_141, w_004_011);
  not1 I007_275(w_007_275, w_000_776);
  and2 I007_276(w_007_276, w_002_090, w_003_125);
  not1 I007_277(w_007_277, w_002_452);
  nand2 I007_278(w_007_278, w_006_209, w_004_014);
  or2  I007_280(w_007_280, w_001_308, w_005_293);
  or2  I007_281(w_007_281, w_005_539, w_000_549);
  not1 I007_282(w_007_282, w_001_325);
  not1 I007_283(w_007_283, w_003_040);
  nand2 I007_284(w_007_284, w_003_160, w_001_768);
  nand2 I007_286(w_007_286, w_004_016, w_003_160);
  not1 I007_287(w_007_287, w_005_273);
  nand2 I007_288(w_007_288, w_006_060, w_003_209);
  and2 I007_293(w_007_293, w_001_684, w_002_465);
  or2  I007_294(w_007_294, w_000_587, w_002_386);
  or2  I007_295(w_007_295, w_003_146, w_000_609);
  and2 I007_296(w_007_296, w_001_224, w_003_046);
  or2  I007_297(w_007_297, w_003_211, w_000_047);
  and2 I007_298(w_007_298, w_000_394, w_002_224);
  not1 I007_299(w_007_299, w_005_285);
  nand2 I007_301(w_007_301, w_004_016, w_003_065);
  not1 I007_302(w_007_302, w_005_315);
  nand2 I007_303(w_007_303, w_006_260, w_006_250);
  nand2 I007_304(w_007_304, w_001_277, w_006_187);
  and2 I007_306(w_007_306, w_004_010, w_000_075);
  and2 I007_307(w_007_307, w_006_087, w_002_130);
  not1 I007_308(w_007_308, w_006_164);
  or2  I007_309(w_007_309, w_002_387, w_002_333);
  or2  I007_310(w_007_310, w_006_099, w_000_236);
  or2  I007_311(w_007_311, w_006_108, w_004_029);
  and2 I007_313(w_007_313, w_000_849, w_000_120);
  not1 I007_314(w_007_314, w_002_100);
  or2  I007_315(w_007_315, w_006_264, w_002_342);
  or2  I007_316(w_007_316, w_002_028, w_000_779);
  or2  I007_317(w_007_317, w_000_015, w_000_912);
  or2  I007_318(w_007_318, w_005_084, w_001_484);
  not1 I007_319(w_007_319, w_005_035);
  not1 I007_321(w_007_321, w_001_029);
  nand2 I007_322(w_007_322, w_006_191, w_000_073);
  or2  I007_324(w_007_324, w_002_002, w_002_402);
  not1 I007_327(w_007_327, w_006_311);
  and2 I007_328(w_007_328, w_000_238, w_006_075);
  not1 I007_329(w_007_329, w_006_168);
  or2  I007_331(w_007_331, w_005_049, w_000_423);
  and2 I007_332(w_007_332, w_003_006, w_000_324);
  nand2 I007_333(w_007_333, w_006_016, w_000_223);
  and2 I007_335(w_007_335, w_002_117, w_002_274);
  and2 I007_336(w_007_336, w_006_010, w_002_258);
  not1 I007_337(w_007_337, w_000_777);
  and2 I007_338(w_007_338, w_005_201, w_000_914);
  or2  I007_340(w_007_340, w_000_221, w_006_187);
  nand2 I007_341(w_007_341, w_003_059, w_006_302);
  not1 I007_342(w_007_342, w_001_576);
  not1 I007_343(w_007_343, w_006_271);
  not1 I007_345(w_007_345, w_003_148);
  not1 I007_346(w_007_346, w_004_016);
  not1 I007_347(w_007_347, w_004_019);
  and2 I007_348(w_007_348, w_005_320, w_005_271);
  and2 I007_349(w_007_349, w_003_092, w_002_341);
  not1 I007_350(w_007_350, w_001_515);
  nand2 I007_351(w_007_351, w_006_255, w_001_188);
  nand2 I007_352(w_007_352, w_006_295, w_003_074);
  or2  I007_353(w_007_353, w_006_208, w_000_197);
  not1 I007_356(w_007_356, w_006_091);
  and2 I007_357(w_007_357, w_001_607, w_001_361);
  not1 I007_358(w_007_358, w_003_223);
  not1 I007_359(w_007_359, w_000_862);
  nand2 I007_360(w_007_360, w_003_041, w_005_450);
  nand2 I007_361(w_007_361, w_001_069, w_000_915);
  or2  I007_362(w_007_362, w_001_505, w_000_273);
  not1 I007_363(w_007_363, w_006_127);
  and2 I007_364(w_007_364, w_001_023, w_005_281);
  nand2 I007_365(w_007_365, w_005_070, w_001_074);
  and2 I007_366(w_007_366, w_006_270, w_000_504);
  nand2 I007_367(w_007_367, w_004_018, w_005_133);
  not1 I007_369(w_007_369, w_005_242);
  and2 I007_371(w_007_371, w_003_163, w_004_028);
  and2 I007_373(w_007_373, w_002_334, w_003_039);
  not1 I007_374(w_007_374, w_001_525);
  not1 I007_375(w_007_375, w_003_198);
  and2 I007_376(w_007_376, w_005_410, w_002_041);
  not1 I007_377(w_007_377, w_005_410);
  nand2 I007_378(w_007_378, w_002_305, w_003_210);
  or2  I007_381(w_007_381, w_001_306, w_005_266);
  or2  I007_383(w_007_383, w_006_156, w_002_056);
  nand2 I007_384(w_007_384, w_000_329, w_003_130);
  not1 I007_385(w_007_385, w_003_072);
  and2 I007_386(w_007_386, w_000_802, w_001_382);
  and2 I007_387(w_007_387, w_002_052, w_004_032);
  and2 I007_388(w_007_388, w_003_166, w_002_255);
  and2 I007_390(w_007_390, w_006_060, w_002_104);
  or2  I007_391(w_007_391, w_005_235, w_001_074);
  nand2 I007_392(w_007_392, w_001_472, w_005_431);
  not1 I007_393(w_007_393, w_005_269);
  and2 I007_394(w_007_394, w_001_847, w_003_032);
  and2 I007_395(w_007_395, w_003_137, w_004_029);
  or2  I007_398(w_007_398, w_002_304, w_001_277);
  and2 I007_399(w_007_399, w_006_061, w_005_150);
  not1 I007_400(w_007_400, w_000_561);
  or2  I007_401(w_007_401, w_001_048, w_006_163);
  not1 I007_402(w_007_402, w_001_480);
  not1 I007_403(w_007_403, w_002_449);
  nand2 I007_404(w_007_404, w_006_182, w_002_471);
  and2 I007_405(w_007_405, w_001_854, w_001_213);
  nand2 I007_406(w_007_406, w_001_341, w_006_273);
  and2 I007_407(w_007_407, w_000_603, w_006_103);
  and2 I007_408(w_007_408, w_000_400, w_004_006);
  nand2 I007_409(w_007_409, w_005_227, w_002_322);
  nand2 I007_411(w_007_411, w_002_017, w_003_223);
  nand2 I007_413(w_007_413, w_000_917, w_002_179);
  or2  I007_414(w_007_414, w_006_114, w_004_016);
  or2  I007_415(w_007_415, w_001_700, w_004_036);
  nand2 I007_416(w_007_416, w_004_009, w_000_386);
  or2  I007_417(w_007_417, w_000_142, w_003_033);
  nand2 I007_418(w_007_418, w_006_150, w_002_009);
  and2 I007_419(w_007_419, w_003_120, w_003_008);
  nand2 I007_420(w_007_420, w_000_632, w_003_046);
  or2  I007_421(w_007_421, w_004_027, w_005_056);
  nand2 I007_422(w_007_422, w_001_366, w_004_029);
  and2 I007_423(w_007_423, w_003_065, w_004_008);
  or2  I007_425(w_007_425, w_002_162, w_000_891);
  nand2 I007_426(w_007_426, w_000_211, w_005_359);
  not1 I007_427(w_007_427, w_000_622);
  and2 I007_428(w_007_428, w_003_031, w_004_020);
  or2  I007_430(w_007_430, w_006_104, w_003_152);
  not1 I007_431(w_007_431, w_005_075);
  nand2 I007_432(w_007_432, w_000_164, w_004_016);
  nand2 I007_433(w_007_433, w_004_034, w_000_123);
  not1 I007_435(w_007_435, w_002_129);
  not1 I007_436(w_007_436, w_005_526);
  nand2 I007_437(w_007_437, w_000_675, w_001_755);
  not1 I007_438(w_007_438, w_001_457);
  not1 I007_446(w_007_446, w_000_873);
  and2 I007_447(w_007_447, w_000_449, w_001_658);
  not1 I007_448(w_007_448, w_001_275);
  or2  I007_450(w_007_450, w_003_210, w_001_088);
  nand2 I007_451(w_007_451, w_000_310, w_002_093);
  not1 I007_454(w_007_454, w_006_031);
  and2 I007_456(w_007_456, w_004_017, w_003_043);
  or2  I007_459(w_007_459, w_001_035, w_006_292);
  nand2 I007_460(w_007_460, w_005_012, w_001_719);
  and2 I007_463(w_007_463, w_000_531, w_005_110);
  and2 I007_464(w_007_464, w_003_013, w_002_483);
  not1 I007_472(w_007_472, w_000_918);
  and2 I007_475(w_007_475, w_002_428, w_001_767);
  or2  I007_476(w_007_476, w_002_275, w_006_034);
  or2  I007_484(w_007_484, w_002_154, w_001_478);
  not1 I007_485(w_007_485, w_000_370);
  not1 I007_487(w_007_487, w_000_865);
  and2 I007_488(w_007_488, w_006_310, w_000_741);
  nand2 I007_489(w_007_489, w_001_481, w_004_028);
  and2 I007_491(w_007_491, w_003_030, w_002_189);
  not1 I007_495(w_007_495, w_002_153);
  and2 I007_497(w_007_497, w_000_431, w_001_671);
  not1 I007_499(w_007_499, w_003_225);
  nand2 I007_500(w_007_500, w_004_013, w_000_592);
  not1 I007_501(w_007_501, w_001_026);
  or2  I007_504(w_007_504, w_000_584, w_001_098);
  not1 I007_507(w_007_507, w_003_116);
  or2  I007_509(w_007_509, w_006_288, w_002_434);
  nand2 I007_511(w_007_511, w_002_172, w_004_019);
  and2 I007_512(w_007_512, w_002_224, w_005_349);
  and2 I007_513(w_007_513, w_001_393, w_004_001);
  or2  I007_515(w_007_515, w_005_063, w_005_006);
  not1 I007_517(w_007_517, w_001_726);
  nand2 I007_524(w_007_524, w_006_233, w_002_046);
  and2 I007_526(w_007_526, w_001_852, w_003_038);
  and2 I007_532(w_007_532, w_001_723, w_005_354);
  nand2 I007_535(w_007_535, w_000_301, w_005_521);
  and2 I007_537(w_007_537, w_001_524, w_005_282);
  and2 I007_538(w_007_538, w_004_002, w_005_029);
  nand2 I007_539(w_007_539, w_001_071, w_006_168);
  not1 I007_540(w_007_540, w_001_469);
  or2  I007_543(w_007_543, w_005_242, w_003_073);
  nand2 I007_546(w_007_546, w_002_146, w_005_284);
  and2 I007_549(w_007_549, w_003_158, w_001_259);
  not1 I007_551(w_007_551, w_001_395);
  or2  I007_552(w_007_552, w_001_245, w_005_086);
  and2 I007_553(w_007_553, w_005_233, w_006_243);
  nand2 I007_554(w_007_554, w_006_287, w_003_128);
  nand2 I007_556(w_007_556, w_005_411, w_000_686);
  not1 I007_558(w_007_558, w_001_638);
  nand2 I007_559(w_007_559, w_004_037, w_003_073);
  and2 I008_001(w_008_001, w_007_149, w_003_172);
  nand2 I008_002(w_008_002, w_004_022, w_005_128);
  not1 I008_004(w_008_004, w_007_108);
  and2 I008_006(w_008_006, w_004_024, w_004_021);
  and2 I008_007(w_008_007, w_003_149, w_004_026);
  not1 I008_010(w_008_010, w_002_140);
  or2  I008_012(w_008_012, w_001_001, w_002_149);
  or2  I008_013(w_008_013, w_003_055, w_001_081);
  not1 I008_015(w_008_015, w_006_064);
  not1 I008_016(w_008_016, w_006_263);
  or2  I008_017(w_008_017, w_004_010, w_004_019);
  and2 I008_018(w_008_018, w_003_086, w_005_063);
  nand2 I008_021(w_008_021, w_001_395, w_005_195);
  and2 I008_022(w_008_022, w_000_042, w_006_286);
  and2 I008_023(w_008_023, w_005_549, w_001_753);
  nand2 I008_024(w_008_024, w_006_319, w_003_195);
  nand2 I008_025(w_008_025, w_001_039, w_004_027);
  not1 I008_026(w_008_026, w_007_556);
  not1 I008_028(w_008_028, w_005_163);
  and2 I008_030(w_008_030, w_004_027, w_005_385);
  and2 I008_033(w_008_033, w_000_191, w_003_137);
  nand2 I008_034(w_008_034, w_001_019, w_007_559);
  or2  I008_035(w_008_035, w_005_074, w_007_195);
  or2  I008_036(w_008_036, w_000_031, w_001_613);
  and2 I008_037(w_008_037, w_007_156, w_004_011);
  or2  I008_038(w_008_038, w_003_001, w_002_244);
  or2  I008_043(w_008_043, w_003_167, w_001_362);
  nand2 I008_044(w_008_044, w_005_036, w_005_281);
  or2  I008_046(w_008_046, w_002_455, w_002_445);
  and2 I008_049(w_008_049, w_002_110, w_001_685);
  or2  I008_050(w_008_050, w_002_047, w_001_711);
  and2 I008_051(w_008_051, w_006_253, w_007_213);
  not1 I008_053(w_008_053, w_007_134);
  and2 I008_054(w_008_054, w_007_213, w_001_441);
  nand2 I008_056(w_008_056, w_004_019, w_000_854);
  or2  I008_061(w_008_061, w_004_006, w_004_016);
  not1 I008_064(w_008_064, w_004_034);
  nand2 I008_067(w_008_067, w_002_467, w_001_755);
  and2 I008_069(w_008_069, w_005_086, w_001_151);
  nand2 I008_071(w_008_071, w_001_155, w_007_188);
  not1 I008_072(w_008_072, w_001_589);
  or2  I008_073(w_008_073, w_007_203, w_005_495);
  not1 I008_074(w_008_074, w_007_252);
  or2  I008_077(w_008_077, w_003_135, w_005_329);
  nand2 I008_078(w_008_078, w_006_059, w_002_080);
  not1 I008_079(w_008_079, w_003_167);
  and2 I008_084(w_008_084, w_004_001, w_002_451);
  or2  I008_086(w_008_086, w_003_002, w_004_036);
  not1 I008_088(w_008_088, w_001_103);
  or2  I008_090(w_008_090, w_006_148, w_000_283);
  and2 I008_092(w_008_092, w_000_302, w_005_135);
  nand2 I008_096(w_008_096, w_005_352, w_001_827);
  not1 I008_097(w_008_097, w_001_462);
  and2 I008_100(w_008_100, w_002_305, w_006_321);
  or2  I008_102(w_008_102, w_000_194, w_006_241);
  and2 I008_104(w_008_104, w_000_628, w_007_161);
  not1 I008_107(w_008_107, w_006_060);
  or2  I008_108(w_008_108, w_001_647, w_004_016);
  and2 I008_109(w_008_109, w_005_288, w_006_246);
  nand2 I008_116(w_008_116, w_005_287, w_003_111);
  not1 I008_118(w_008_118, w_001_890);
  or2  I008_122(w_008_122, w_006_235, w_005_123);
  nand2 I008_126(w_008_126, w_006_035, w_000_079);
  nand2 I008_129(w_008_129, w_006_239, w_007_222);
  nand2 I008_130(w_008_130, w_000_657, w_004_033);
  and2 I008_131(w_008_131, w_007_540, w_002_367);
  or2  I008_133(w_008_133, w_007_392, w_006_182);
  and2 I008_134(w_008_134, w_005_254, w_004_025);
  nand2 I008_135(w_008_135, w_006_018, w_007_284);
  and2 I008_138(w_008_138, w_004_025, w_002_491);
  and2 I008_142(w_008_142, w_003_060, w_007_431);
  or2  I008_143(w_008_143, w_005_043, w_002_435);
  nand2 I008_145(w_008_145, w_004_023, w_001_408);
  nand2 I008_147(w_008_147, w_003_042, w_000_747);
  and2 I008_149(w_008_149, w_003_143, w_001_409);
  nand2 I008_154(w_008_154, w_001_050, w_003_052);
  not1 I008_155(w_008_155, w_000_090);
  not1 I008_156(w_008_156, w_000_314);
  and2 I008_158(w_008_158, w_003_058, w_004_008);
  not1 I008_161(w_008_161, w_004_001);
  and2 I008_163(w_008_163, w_001_423, w_001_684);
  not1 I008_167(w_008_167, w_003_068);
  or2  I008_168(w_008_168, w_007_155, w_004_006);
  nand2 I008_169(w_008_169, w_004_020, w_003_045);
  not1 I008_170(w_008_170, w_004_003);
  or2  I008_172(w_008_172, w_000_878, w_005_217);
  and2 I008_174(w_008_174, w_003_062, w_001_370);
  and2 I008_176(w_008_176, w_003_003, w_007_240);
  not1 I008_178(w_008_178, w_004_036);
  and2 I008_179(w_008_179, w_001_063, w_001_559);
  not1 I008_182(w_008_182, w_002_350);
  or2  I008_184(w_008_184, w_004_004, w_005_005);
  nand2 I008_186(w_008_186, w_001_349, w_005_482);
  not1 I008_187(w_008_187, w_004_007);
  and2 I008_188(w_008_188, w_007_367, w_004_005);
  nand2 I008_191(w_008_191, w_003_024, w_005_190);
  nand2 I008_192(w_008_192, w_006_255, w_007_192);
  not1 I008_194(w_008_194, w_003_160);
  or2  I008_200(w_008_200, w_005_128, w_005_200);
  or2  I008_202(w_008_202, w_005_149, w_005_570);
  and2 I008_209(w_008_209, w_007_336, w_006_251);
  not1 I008_210(w_008_210, w_002_298);
  and2 I008_211(w_008_211, w_000_586, w_005_119);
  or2  I008_213(w_008_213, w_004_022, w_000_370);
  nand2 I008_215(w_008_215, w_003_092, w_007_099);
  nand2 I008_216(w_008_216, w_006_243, w_005_121);
  not1 I008_217(w_008_217, w_005_337);
  and2 I008_218(w_008_218, w_002_456, w_004_010);
  or2  I008_220(w_008_220, w_007_233, w_006_218);
  not1 I008_222(w_008_222, w_005_467);
  or2  I008_225(w_008_225, w_006_137, w_006_144);
  and2 I008_226(w_008_226, w_004_007, w_005_196);
  nand2 I008_227(w_008_227, w_004_032, w_006_223);
  or2  I008_230(w_008_230, w_006_212, w_006_319);
  nand2 I008_231(w_008_231, w_003_093, w_000_209);
  or2  I008_232(w_008_232, w_000_662, w_004_013);
  nand2 I008_234(w_008_234, w_001_406, w_004_006);
  and2 I008_235(w_008_235, w_001_540, w_006_048);
  not1 I008_236(w_008_236, w_007_336);
  and2 I008_237(w_008_237, w_006_234, w_000_529);
  not1 I008_241(w_008_241, w_000_845);
  nand2 I008_242(w_008_242, w_002_385, w_001_732);
  nand2 I008_244(w_008_244, w_004_008, w_000_917);
  or2  I008_246(w_008_246, w_006_307, w_006_069);
  nand2 I008_247(w_008_247, w_002_344, w_002_362);
  or2  I008_251(w_008_251, w_000_443, w_007_060);
  or2  I008_252(w_008_252, w_004_037, w_000_098);
  or2  I008_253(w_008_253, w_000_596, w_005_107);
  not1 I008_254(w_008_254, w_002_125);
  and2 I008_257(w_008_257, w_005_049, w_001_077);
  and2 I008_259(w_008_259, w_001_110, w_001_233);
  not1 I008_260(w_008_260, w_006_249);
  and2 I008_261(w_008_261, w_000_890, w_003_116);
  not1 I008_263(w_008_263, w_003_065);
  not1 I008_264(w_008_264, w_001_367);
  or2  I008_267(w_008_267, w_007_367, w_003_007);
  and2 I008_268(w_008_268, w_003_023, w_005_051);
  and2 I008_269(w_008_269, w_000_609, w_006_281);
  nand2 I008_271(w_008_271, w_003_072, w_003_012);
  nand2 I008_272(w_008_272, w_007_422, w_005_213);
  and2 I008_275(w_008_275, w_003_118, w_004_026);
  and2 I008_276(w_008_276, w_002_372, w_004_029);
  nand2 I008_277(w_008_277, w_004_009, w_006_224);
  and2 I008_278(w_008_278, w_001_688, w_007_160);
  not1 I008_279(w_008_279, w_004_002);
  nand2 I008_280(w_008_280, w_001_459, w_004_022);
  or2  I008_281(w_008_281, w_002_443, w_005_086);
  and2 I008_282(w_008_282, w_001_584, w_004_006);
  not1 I008_283(w_008_283, w_000_191);
  nand2 I008_285(w_008_285, w_000_909, w_007_032);
  nand2 I008_288(w_008_288, w_002_161, w_007_076);
  or2  I008_289(w_008_289, w_003_042, w_000_060);
  not1 I008_294(w_008_294, w_007_031);
  not1 I008_297(w_008_297, w_001_894);
  nand2 I008_299(w_008_299, w_000_865, w_005_094);
  not1 I008_300(w_008_300, w_000_372);
  not1 I008_302(w_008_302, w_001_737);
  not1 I008_303(w_008_303, w_004_024);
  or2  I008_304(w_008_304, w_001_658, w_007_395);
  and2 I008_305(w_008_305, w_001_012, w_007_215);
  or2  I008_306(w_008_306, w_007_230, w_005_088);
  not1 I008_310(w_008_310, w_002_190);
  or2  I008_314(w_008_314, w_000_703, w_004_013);
  or2  I008_318(w_008_318, w_004_035, w_000_610);
  not1 I008_319(w_008_319, w_001_453);
  not1 I008_325(w_008_325, w_005_265);
  and2 I008_326(w_008_326, w_007_085, w_006_325);
  or2  I008_327(w_008_327, w_005_212, w_004_009);
  or2  I008_328(w_008_328, w_003_040, w_004_002);
  nand2 I008_331(w_008_331, w_002_028, w_000_829);
  not1 I008_332(w_008_332, w_006_283);
  nand2 I008_333(w_008_333, w_006_210, w_006_073);
  and2 I008_335(w_008_335, w_003_160, w_003_063);
  nand2 I008_340(w_008_340, w_006_091, w_000_170);
  not1 I008_343(w_008_343, w_003_107);
  nand2 I008_344(w_008_344, w_007_421, w_005_228);
  or2  I008_346(w_008_346, w_005_319, w_002_324);
  or2  I008_347(w_008_347, w_005_415, w_003_154);
  and2 I008_348(w_008_348, w_001_080, w_007_067);
  and2 I008_349(w_008_349, w_002_219, w_002_035);
  and2 I008_354(w_008_354, w_005_035, w_004_017);
  and2 I008_355(w_008_355, w_003_159, w_000_029);
  not1 I008_356(w_008_356, w_002_416);
  and2 I008_358(w_008_358, w_004_012, w_004_019);
  and2 I008_361(w_008_361, w_005_154, w_005_300);
  and2 I008_365(w_008_365, w_004_010, w_007_363);
  or2  I008_373(w_008_373, w_000_655, w_002_254);
  nand2 I008_374(w_008_374, w_001_276, w_002_254);
  nand2 I008_377(w_008_377, w_005_460, w_002_001);
  and2 I008_379(w_008_379, w_002_413, w_003_212);
  and2 I008_383(w_008_383, w_005_102, w_000_071);
  not1 I008_384(w_008_384, w_007_540);
  or2  I008_386(w_008_386, w_000_675, w_000_558);
  or2  I008_387(w_008_387, w_004_017, w_005_274);
  not1 I008_388(w_008_388, w_001_762);
  not1 I008_389(w_008_389, w_006_082);
  not1 I008_392(w_008_392, w_003_047);
  nand2 I008_396(w_008_396, w_004_032, w_002_340);
  nand2 I008_397(w_008_397, w_000_525, w_004_003);
  and2 I008_398(w_008_398, w_001_324, w_002_097);
  not1 I008_400(w_008_400, w_007_105);
  nand2 I008_401(w_008_401, w_003_130, w_006_292);
  or2  I008_405(w_008_405, w_003_152, w_007_476);
  not1 I008_406(w_008_406, w_005_425);
  or2  I008_407(w_008_407, w_004_023, w_004_027);
  and2 I008_408(w_008_408, w_002_120, w_007_286);
  and2 I008_409(w_008_409, w_000_662, w_003_037);
  not1 I008_411(w_008_411, w_004_022);
  not1 I008_414(w_008_414, w_000_655);
  or2  I008_423(w_008_423, w_001_674, w_001_701);
  nand2 I008_425(w_008_425, w_007_416, w_007_374);
  and2 I008_428(w_008_428, w_004_022, w_005_075);
  or2  I008_432(w_008_432, w_005_064, w_005_078);
  not1 I008_434(w_008_434, w_000_071);
  and2 I008_435(w_008_435, w_003_164, w_004_031);
  nand2 I008_437(w_008_437, w_003_130, w_002_030);
  and2 I008_442(w_008_442, w_000_361, w_001_710);
  and2 I008_446(w_008_446, w_007_384, w_007_358);
  not1 I008_447(w_008_447, w_006_257);
  not1 I008_448(w_008_448, w_005_072);
  nand2 I008_450(w_008_450, w_000_697, w_005_261);
  nand2 I008_458(w_008_458, w_000_754, w_004_003);
  and2 I008_459(w_008_459, w_007_205, w_004_012);
  and2 I008_461(w_008_461, w_006_056, w_001_783);
  or2  I008_462(w_008_462, w_004_036, w_005_400);
  not1 I008_466(w_008_466, w_005_160);
  and2 I008_473(w_008_473, w_007_248, w_004_001);
  or2  I008_474(w_008_474, w_004_037, w_002_013);
  or2  I008_477(w_008_477, w_004_011, w_005_309);
  and2 I008_478(w_008_478, w_007_322, w_004_015);
  not1 I008_480(w_008_480, w_000_745);
  nand2 I008_482(w_008_482, w_001_787, w_000_660);
  and2 I008_484(w_008_484, w_001_577, w_001_085);
  not1 I008_485(w_008_485, w_000_320);
  not1 I008_486(w_008_486, w_006_237);
  not1 I008_487(w_008_487, w_002_218);
  not1 I008_488(w_008_488, w_004_023);
  nand2 I008_490(w_008_490, w_000_576, w_002_462);
  and2 I008_491(w_008_491, w_005_376, w_007_338);
  nand2 I008_494(w_008_494, w_003_225, w_005_496);
  nand2 I008_496(w_008_496, w_006_132, w_003_202);
  not1 I008_497(w_008_497, w_007_077);
  nand2 I008_499(w_008_499, w_006_331, w_005_157);
  or2  I008_501(w_008_501, w_002_015, w_003_098);
  or2  I008_503(w_008_503, w_002_175, w_007_072);
  and2 I008_505(w_008_505, w_001_403, w_005_034);
  not1 I008_510(w_008_510, w_005_195);
  nand2 I008_514(w_008_514, w_007_517, w_001_562);
  or2  I008_515(w_008_515, w_006_317, w_000_268);
  and2 I008_517(w_008_517, w_007_284, w_003_157);
  not1 I008_520(w_008_520, w_002_061);
  or2  I008_527(w_008_527, w_003_108, w_000_820);
  not1 I008_528(w_008_528, w_005_213);
  and2 I008_529(w_008_529, w_005_117, w_007_031);
  nand2 I008_534(w_008_534, w_000_516, w_007_108);
  or2  I008_542(w_008_542, w_003_009, w_006_156);
  nand2 I008_545(w_008_545, w_007_321, w_007_129);
  and2 I008_548(w_008_548, w_003_011, w_003_183);
  or2  I008_553(w_008_553, w_000_422, w_000_786);
  not1 I008_555(w_008_555, w_005_176);
  and2 I008_557(w_008_557, w_001_462, w_001_199);
  nand2 I008_559(w_008_559, w_004_015, w_007_152);
  nand2 I008_560(w_008_560, w_007_366, w_003_223);
  not1 I008_562(w_008_562, w_006_311);
  and2 I008_565(w_008_565, w_003_036, w_007_265);
  nand2 I008_566(w_008_566, w_004_018, w_004_017);
  nand2 I008_567(w_008_567, w_004_027, w_006_307);
  and2 I008_568(w_008_568, w_007_337, w_007_109);
  nand2 I008_574(w_008_574, w_006_136, w_004_026);
  nand2 I008_575(w_008_575, w_007_299, w_001_155);
  or2  I008_578(w_008_578, w_003_200, w_005_171);
  or2  I008_581(w_008_581, w_006_218, w_005_363);
  or2  I008_582(w_008_582, w_004_027, w_002_045);
  and2 I008_585(w_008_585, w_003_139, w_001_414);
  not1 I008_586(w_008_586, w_003_186);
  nand2 I008_588(w_008_588, w_005_243, w_000_136);
  or2  I008_591(w_008_591, w_003_188, w_001_230);
  or2  I008_595(w_008_595, w_005_371, w_000_796);
  not1 I008_596(w_008_596, w_005_219);
  nand2 I008_597(w_008_597, w_000_820, w_004_011);
  and2 I008_598(w_008_598, w_006_220, w_003_195);
  not1 I008_599(w_008_599, w_000_703);
  not1 I008_600(w_008_600, w_005_142);
  or2  I008_601(w_008_601, w_001_684, w_006_162);
  not1 I008_604(w_008_604, w_002_473);
  nand2 I008_608(w_008_608, w_003_122, w_005_000);
  not1 I008_609(w_008_609, w_007_262);
  not1 I008_610(w_008_610, w_003_089);
  and2 I008_611(w_008_611, w_000_924, w_000_874);
  or2  I008_613(w_008_613, w_004_009, w_007_298);
  nand2 I008_615(w_008_615, w_002_171, w_000_362);
  or2  I008_616(w_008_616, w_000_184, w_004_001);
  or2  I008_619(w_008_619, w_000_873, w_002_139);
  nand2 I008_620(w_008_620, w_002_437, w_004_000);
  nand2 I008_621(w_008_621, w_003_213, w_002_341);
  and2 I008_629(w_008_629, w_006_046, w_001_014);
  and2 I008_631(w_008_631, w_001_428, w_000_357);
  and2 I008_632(w_008_632, w_001_217, w_005_556);
  nand2 I008_633(w_008_633, w_001_858, w_003_167);
  not1 I008_636(w_008_636, w_006_020);
  not1 I008_638(w_008_638, w_001_184);
  and2 I008_642(w_008_642, w_000_176, w_002_232);
  or2  I008_645(w_008_645, w_001_322, w_006_188);
  or2  I008_646(w_008_646, w_000_275, w_005_311);
  nand2 I008_647(w_008_647, w_002_327, w_007_273);
  not1 I008_651(w_008_651, w_002_310);
  or2  I008_652(w_008_652, w_001_681, w_002_031);
  and2 I008_654(w_008_654, w_003_019, w_005_390);
  and2 I008_655(w_008_655, w_007_136, w_005_316);
  or2  I008_656(w_008_656, w_001_030, w_005_057);
  nand2 I008_658(w_008_658, w_003_046, w_001_061);
  or2  I008_661(w_008_661, w_005_124, w_001_580);
  nand2 I008_662(w_008_662, w_006_138, w_000_447);
  nand2 I008_665(w_008_665, w_000_397, w_003_200);
  or2  I008_666(w_008_666, w_003_211, w_007_411);
  or2  I008_668(w_008_668, w_003_000, w_004_017);
  nand2 I008_669(w_008_669, w_002_439, w_000_835);
  not1 I008_670(w_008_670, w_000_926);
  nand2 I008_671(w_008_671, w_007_335, w_003_212);
  and2 I008_672(w_008_672, w_006_228, w_005_265);
  and2 I008_674(w_008_674, w_001_663, w_001_380);
  nand2 I008_675(w_008_675, w_006_318, w_006_078);
  or2  I008_676(w_008_676, w_006_265, w_003_128);
  nand2 I008_677(w_008_677, w_003_170, w_002_446);
  not1 I008_678(w_008_678, w_006_178);
  and2 I008_679(w_008_679, w_003_009, w_001_095);
  or2  I008_680(w_008_680, w_003_062, w_005_062);
  or2  I008_681(w_008_681, w_007_017, w_004_038);
  or2  I008_682(w_008_682, w_002_445, w_003_065);
  or2  I008_684(w_008_684, w_005_015, w_003_175);
  nand2 I008_685(w_008_685, w_007_047, w_000_417);
  not1 I008_689(w_008_689, w_000_758);
  or2  I008_690(w_008_690, w_004_015, w_007_233);
  and2 I008_692(w_008_692, w_003_067, w_003_092);
  or2  I008_694(w_008_694, w_004_034, w_004_022);
  and2 I008_702(w_008_702, w_004_015, w_005_018);
  and2 I008_703(w_008_703, w_004_000, w_005_066);
  or2  I008_704(w_008_704, w_002_351, w_004_005);
  or2  I008_706(w_008_706, w_005_223, w_003_154);
  not1 I008_707(w_008_707, w_007_132);
  and2 I008_708(w_008_708, w_007_278, w_000_499);
  nand2 I008_712(w_008_712, w_001_456, w_005_350);
  and2 I008_714(w_008_714, w_001_382, w_002_186);
  or2  I008_717(w_008_717, w_003_215, w_002_460);
  and2 I008_718(w_008_718, w_003_169, w_003_092);
  not1 I008_720(w_008_720, w_005_480);
  or2  I008_722(w_008_722, w_004_023, w_000_726);
  nand2 I008_727(w_008_727, w_003_038, w_001_827);
  nand2 I008_734(w_008_734, w_007_310, w_000_175);
  and2 I008_735(w_008_735, w_007_472, w_004_007);
  nand2 I008_737(w_008_737, w_001_076, w_005_061);
  not1 I008_739(w_008_739, w_004_038);
  or2  I008_746(w_008_746, w_002_151, w_002_099);
  and2 I008_747(w_008_747, w_005_363, w_004_037);
  not1 I008_748(w_008_748, w_001_080);
  not1 I008_749(w_008_749, w_005_532);
  not1 I008_750(w_008_750, w_003_139);
  or2  I008_756(w_008_756, w_003_030, w_007_391);
  or2  I008_758(w_008_758, w_003_147, w_006_121);
  and2 I008_759(w_008_759, w_002_306, w_002_005);
  nand2 I008_760(w_008_760, w_006_202, w_004_037);
  nand2 I008_761(w_008_761, w_001_751, w_002_472);
  nand2 I008_764(w_008_764, w_003_189, w_001_734);
  or2  I008_765(w_008_765, w_007_208, w_005_250);
  not1 I008_768(w_008_768, w_003_059);
  and2 I008_769(w_008_769, w_003_083, w_003_150);
  and2 I008_770(w_008_770, w_001_761, w_003_059);
  and2 I008_771(w_008_771, w_006_172, w_001_508);
  not1 I008_772(w_008_772, w_001_716);
  nand2 I008_773(w_008_773, w_002_085, w_002_331);
  not1 I008_779(w_008_779, w_002_409);
  or2  I008_780(w_008_780, w_004_038, w_005_308);
  or2  I008_785(w_008_785, w_000_766, w_003_050);
  or2  I008_790(w_008_790, w_003_040, w_004_027);
  nand2 I008_792(w_008_792, w_006_130, w_003_005);
  nand2 I008_793(w_008_793, w_005_084, w_004_002);
  and2 I008_794(w_008_794, w_006_007, w_007_099);
  nand2 I008_795(w_008_795, w_002_261, w_006_263);
  not1 I008_803(w_008_803, w_005_375);
  not1 I008_804(w_008_804, w_005_088);
  or2  I008_806(w_008_806, w_000_484, w_000_837);
  not1 I008_808(w_008_808, w_004_027);
  not1 I008_810(w_008_810, w_006_104);
  not1 I008_813(w_008_813, w_004_011);
  nand2 I008_814(w_008_814, w_001_486, w_005_033);
  not1 I008_815(w_008_815, w_005_296);
  or2  I008_820(w_008_820, w_006_255, w_001_296);
  or2  I008_822(w_008_822, w_006_243, w_006_084);
  and2 I008_824(w_008_824, w_005_386, w_005_098);
  not1 I008_826(w_008_826, w_004_028);
  nand2 I008_827(w_008_827, w_005_062, w_000_296);
  and2 I008_828(w_008_828, w_001_669, w_005_009);
  and2 I008_829(w_008_829, w_004_022, w_001_068);
  and2 I008_830(w_008_830, w_002_496, w_000_551);
  not1 I008_832(w_008_832, w_006_225);
  not1 I008_835(w_008_835, w_001_023);
  and2 I008_836(w_008_836, w_001_039, w_004_012);
  or2  I008_837(w_008_837, w_001_030, w_003_009);
  not1 I008_840(w_008_840, w_002_026);
  not1 I008_848(w_008_848, w_004_018);
  or2  I008_850(w_008_850, w_001_436, w_005_515);
  not1 I008_853(w_008_853, w_004_028);
  not1 I008_857(w_008_857, w_000_583);
  not1 I008_861(w_008_861, w_001_234);
  not1 I008_862(w_008_862, w_007_074);
  nand2 I008_863(w_008_863, w_000_210, w_006_203);
  or2  I008_864(w_008_864, w_004_025, w_007_103);
  or2  I008_866(w_008_866, w_006_321, w_003_112);
  or2  I008_874(w_008_874, w_001_083, w_006_128);
  and2 I008_877(w_008_877, w_005_260, w_004_008);
  nand2 I008_878(w_008_878, w_002_360, w_007_554);
  and2 I008_879(w_008_879, w_007_040, w_005_399);
  not1 I008_880(w_008_880, w_005_322);
  and2 I008_881(w_008_881, w_006_303, w_006_095);
  not1 I008_882(w_008_882, w_006_052);
  and2 I008_884(w_008_884, w_005_142, w_000_932);
  or2  I008_885(w_008_885, w_003_208, w_000_325);
  and2 I008_886(w_008_886, w_000_717, w_001_366);
  nand2 I008_888(w_008_888, w_006_116, w_001_716);
  not1 I008_889(w_008_889, w_003_201);
  not1 I008_890(w_008_890, w_003_156);
  not1 I008_891(w_008_891, w_001_524);
  nand2 I008_892(w_008_892, w_005_525, w_006_002);
  not1 I008_893(w_008_893, w_003_172);
  not1 I008_894(w_008_894, w_000_688);
  and2 I008_896(w_008_896, w_004_009, w_001_845);
  not1 I008_897(w_008_897, w_007_064);
  not1 I008_898(w_008_898, w_005_189);
  and2 I008_899(w_008_899, w_007_245, w_001_642);
  not1 I008_900(w_008_900, w_006_088);
  not1 I008_906(w_008_906, w_001_092);
  or2  I008_908(w_008_908, w_000_934, w_005_419);
  nand2 I008_910(w_008_910, w_007_450, w_003_100);
  not1 I008_912(w_008_912, w_005_201);
  nand2 I008_914(w_008_914, w_005_164, w_005_317);
  or2  I008_917(w_008_917, w_007_430, w_004_035);
  not1 I008_918(w_008_918, w_005_197);
  nand2 I008_919(w_008_919, w_002_014, w_000_794);
  not1 I008_920(w_008_920, w_006_246);
  nand2 I008_921(w_008_921, w_005_459, w_004_004);
  and2 I008_922(w_008_922, w_002_178, w_003_012);
  or2  I008_923(w_008_923, w_007_024, w_001_603);
  nand2 I008_925(w_008_925, w_002_049, w_002_323);
  nand2 I008_926(w_008_926, w_002_469, w_006_177);
  nand2 I008_927(w_008_927, w_005_335, w_003_011);
  not1 I008_930(w_008_930, w_003_073);
  nand2 I008_931(w_008_931, w_004_018, w_004_017);
  or2  I008_933(w_008_933, w_006_174, w_007_543);
  or2  I008_935(w_008_935, w_005_539, w_001_881);
  nand2 I008_936(w_008_936, w_007_303, w_005_366);
  not1 I008_939(w_008_939, w_006_288);
  nand2 I008_941(w_008_941, w_002_215, w_005_559);
  nand2 I008_943(w_008_943, w_005_107, w_004_009);
  not1 I008_947(w_008_947, w_001_722);
  or2  I008_949(w_008_949, w_000_907, w_001_430);
  nand2 I008_951(w_008_951, w_004_011, w_007_318);
  and2 I008_952(w_008_952, w_000_572, w_000_863);
  and2 I008_953(w_008_953, w_002_144, w_003_063);
  nand2 I008_955(w_008_955, w_007_239, w_006_319);
  nand2 I008_959(w_008_959, w_005_476, w_007_023);
  not1 I009_000(w_009_000, w_000_387);
  and2 I009_001(w_009_001, w_002_434, w_003_067);
  not1 I009_002(w_009_002, w_008_874);
  nand2 I009_003(w_009_003, w_007_384, w_003_032);
  not1 I009_004(w_009_004, w_002_217);
  nand2 I009_005(w_009_005, w_004_014, w_003_197);
  or2  I009_006(w_009_006, w_003_099, w_008_143);
  and2 I009_007(w_009_007, w_007_381, w_005_109);
  or2  I009_008(w_009_008, w_007_393, w_006_195);
  nand2 I009_009(w_009_009, w_005_402, w_001_479);
  nand2 I009_010(w_009_010, w_005_388, w_007_171);
  and2 I009_011(w_009_011, w_005_178, w_003_084);
  or2  I009_012(w_009_012, w_002_217, w_002_254);
  and2 I009_013(w_009_013, w_000_936, w_000_112);
  or2  I009_014(w_009_014, w_003_121, w_005_121);
  or2  I009_015(w_009_015, w_001_276, w_000_157);
  nand2 I009_016(w_009_016, w_006_238, w_001_050);
  nand2 I009_017(w_009_017, w_005_328, w_002_461);
  and2 I009_018(w_009_018, w_006_248, w_004_030);
  nand2 I009_019(w_009_019, w_002_179, w_000_602);
  or2  I009_020(w_009_020, w_000_152, w_000_432);
  not1 I009_021(w_009_021, w_008_638);
  not1 I009_022(w_009_022, w_007_147);
  or2  I009_023(w_009_023, w_004_012, w_003_091);
  not1 I009_024(w_009_024, w_008_645);
  and2 I009_025(w_009_025, w_006_313, w_000_781);
  nand2 I009_026(w_009_026, w_006_303, w_005_275);
  and2 I009_027(w_009_027, w_006_325, w_007_399);
  not1 I009_028(w_009_028, w_001_585);
  or2  I009_029(w_009_029, w_004_020, w_006_007);
  and2 I009_030(w_009_030, w_002_059, w_006_325);
  or2  I009_031(w_009_031, w_003_184, w_004_008);
  or2  I009_032(w_009_032, w_002_150, w_003_119);
  or2  I009_033(w_009_033, w_000_647, w_005_512);
  nand2 I009_034(w_009_034, w_002_471, w_002_262);
  or2  I009_035(w_009_035, w_008_620, w_006_265);
  and2 I009_036(w_009_036, w_007_045, w_003_051);
  and2 I009_037(w_009_037, w_004_006, w_006_142);
  not1 I009_038(w_009_038, w_006_118);
  not1 I009_039(w_009_039, w_001_268);
  nand2 I009_040(w_009_040, w_001_267, w_007_099);
  not1 I009_041(w_009_041, w_000_482);
  nand2 I009_042(w_009_042, w_002_243, w_007_156);
  and2 I009_043(w_009_043, w_002_198, w_007_526);
  nand2 I009_044(w_009_044, w_000_474, w_008_769);
  not1 I009_045(w_009_045, w_006_069);
  nand2 I009_046(w_009_046, w_008_349, w_005_456);
  and2 I009_047(w_009_047, w_004_022, w_001_247);
  not1 I009_048(w_009_048, w_001_082);
  not1 I009_049(w_009_049, w_001_325);
  and2 I009_050(w_009_050, w_000_169, w_007_013);
  not1 I009_051(w_009_051, w_006_309);
  and2 I009_052(w_009_052, w_005_310, w_002_315);
  nand2 I009_053(w_009_053, w_007_402, w_004_004);
  and2 I009_054(w_009_054, w_000_679, w_002_474);
  and2 I009_055(w_009_055, w_001_306, w_004_010);
  and2 I009_056(w_009_056, w_005_072, w_002_454);
  or2  I009_057(w_009_057, w_000_028, w_006_306);
  or2  I009_058(w_009_058, w_003_003, w_001_074);
  and2 I009_059(w_009_059, w_006_101, w_007_408);
  not1 I009_060(w_009_060, w_005_216);
  not1 I009_061(w_009_061, w_007_188);
  not1 I009_062(w_009_062, w_006_181);
  nand2 I009_063(w_009_063, w_007_499, w_003_113);
  and2 I009_064(w_009_064, w_004_009, w_005_135);
  or2  I009_065(w_009_065, w_001_176, w_006_213);
  not1 I009_066(w_009_066, w_000_776);
  nand2 I009_067(w_009_067, w_000_937, w_002_089);
  not1 I009_068(w_009_068, w_008_283);
  nand2 I010_002(w_010_002, w_009_025, w_001_165);
  or2  I010_003(w_010_003, w_005_240, w_004_000);
  not1 I010_004(w_010_004, w_006_298);
  not1 I010_005(w_010_005, w_006_225);
  or2  I010_006(w_010_006, w_004_005, w_001_832);
  and2 I010_007(w_010_007, w_009_051, w_004_021);
  or2  I010_008(w_010_008, w_005_032, w_009_009);
  and2 I010_009(w_010_009, w_008_448, w_005_230);
  or2  I010_010(w_010_010, w_002_122, w_001_109);
  nand2 I010_011(w_010_011, w_008_425, w_009_044);
  and2 I010_012(w_010_012, w_001_612, w_008_414);
  and2 I010_013(w_010_013, w_004_020, w_004_001);
  or2  I010_014(w_010_014, w_009_037, w_006_162);
  and2 I010_015(w_010_015, w_000_117, w_002_127);
  not1 I010_016(w_010_016, w_009_011);
  nand2 I010_017(w_010_017, w_003_089, w_002_195);
  not1 I010_018(w_010_018, w_003_063);
  not1 I010_020(w_010_020, w_003_019);
  nand2 I010_021(w_010_021, w_006_017, w_007_250);
  not1 I010_023(w_010_023, w_000_479);
  not1 I010_025(w_010_025, w_000_444);
  not1 I010_027(w_010_027, w_003_137);
  or2  I010_029(w_010_029, w_009_004, w_007_089);
  or2  I010_031(w_010_031, w_002_157, w_000_022);
  or2  I010_033(w_010_033, w_004_016, w_003_139);
  or2  I010_034(w_010_034, w_004_005, w_001_094);
  nand2 I010_035(w_010_035, w_004_010, w_002_453);
  and2 I010_037(w_010_037, w_009_043, w_009_034);
  not1 I010_039(w_010_039, w_005_305);
  not1 I010_040(w_010_040, w_009_019);
  and2 I010_042(w_010_042, w_009_024, w_006_309);
  and2 I010_043(w_010_043, w_005_395, w_002_039);
  not1 I010_044(w_010_044, w_002_419);
  and2 I010_047(w_010_047, w_002_054, w_007_447);
  not1 I010_049(w_010_049, w_009_040);
  not1 I010_050(w_010_050, w_007_348);
  and2 I010_052(w_010_052, w_006_188, w_002_475);
  or2  I010_053(w_010_053, w_007_301, w_001_043);
  and2 I010_054(w_010_054, w_004_035, w_006_031);
  or2  I010_057(w_010_057, w_002_270, w_009_026);
  nand2 I010_058(w_010_058, w_007_079, w_006_309);
  nand2 I010_059(w_010_059, w_002_163, w_002_189);
  or2  I010_060(w_010_060, w_009_065, w_004_003);
  and2 I010_061(w_010_061, w_000_389, w_008_277);
  not1 I010_063(w_010_063, w_008_935);
  not1 I010_065(w_010_065, w_004_017);
  and2 I010_067(w_010_067, w_008_396, w_003_066);
  not1 I010_070(w_010_070, w_006_094);
  or2  I010_072(w_010_072, w_004_027, w_007_427);
  not1 I010_073(w_010_073, w_006_144);
  and2 I010_074(w_010_074, w_007_321, w_006_025);
  and2 I010_077(w_010_077, w_001_066, w_009_003);
  or2  I010_078(w_010_078, w_009_008, w_004_010);
  not1 I010_079(w_010_079, w_008_326);
  or2  I010_080(w_010_080, w_007_144, w_000_574);
  and2 I010_081(w_010_081, w_009_048, w_001_215);
  and2 I010_082(w_010_082, w_008_072, w_008_084);
  not1 I010_084(w_010_084, w_006_278);
  and2 I010_085(w_010_085, w_001_065, w_007_167);
  nand2 I010_086(w_010_086, w_000_281, w_000_656);
  nand2 I010_087(w_010_087, w_007_152, w_005_414);
  and2 I010_088(w_010_088, w_004_026, w_009_037);
  not1 I010_090(w_010_090, w_002_225);
  or2  I010_091(w_010_091, w_000_521, w_005_269);
  nand2 I010_092(w_010_092, w_002_073, w_008_484);
  and2 I010_094(w_010_094, w_006_196, w_001_623);
  nand2 I010_095(w_010_095, w_002_074, w_003_208);
  or2  I010_097(w_010_097, w_005_480, w_008_328);
  or2  I010_099(w_010_099, w_007_183, w_009_025);
  or2  I010_103(w_010_103, w_007_360, w_008_933);
  nand2 I010_107(w_010_107, w_000_548, w_007_024);
  or2  I010_109(w_010_109, w_005_400, w_005_028);
  or2  I010_110(w_010_110, w_008_952, w_008_680);
  nand2 I010_111(w_010_111, w_003_150, w_008_002);
  or2  I010_113(w_010_113, w_003_001, w_003_030);
  not1 I010_114(w_010_114, w_004_002);
  nand2 I010_115(w_010_115, w_001_053, w_000_498);
  not1 I010_116(w_010_116, w_006_121);
  nand2 I010_117(w_010_117, w_004_016, w_000_616);
  or2  I010_118(w_010_118, w_003_088, w_004_033);
  or2  I010_120(w_010_120, w_006_099, w_003_068);
  not1 I010_121(w_010_121, w_007_149);
  or2  I010_122(w_010_122, w_000_554, w_005_394);
  and2 I010_123(w_010_123, w_003_197, w_002_421);
  and2 I010_125(w_010_125, w_000_056, w_008_194);
  and2 I010_127(w_010_127, w_005_373, w_008_682);
  or2  I010_128(w_010_128, w_005_152, w_004_001);
  and2 I010_130(w_010_130, w_007_002, w_006_323);
  not1 I010_132(w_010_132, w_006_182);
  nand2 I010_134(w_010_134, w_000_010, w_000_412);
  not1 I010_136(w_010_136, w_004_025);
  not1 I010_137(w_010_137, w_005_023);
  nand2 I010_139(w_010_139, w_002_194, w_006_247);
  nand2 I010_140(w_010_140, w_008_758, w_000_380);
  or2  I010_141(w_010_141, w_000_390, w_009_056);
  not1 I010_143(w_010_143, w_003_204);
  nand2 I010_144(w_010_144, w_000_843, w_002_175);
  nand2 I010_145(w_010_145, w_003_092, w_009_019);
  and2 I010_146(w_010_146, w_001_677, w_000_650);
  and2 I010_147(w_010_147, w_008_408, w_004_003);
  not1 I010_148(w_010_148, w_004_018);
  or2  I010_152(w_010_152, w_002_280, w_004_033);
  and2 I010_155(w_010_155, w_006_241, w_000_044);
  and2 I010_156(w_010_156, w_003_110, w_008_478);
  and2 I010_157(w_010_157, w_000_475, w_006_211);
  and2 I010_158(w_010_158, w_007_419, w_000_293);
  and2 I010_159(w_010_159, w_004_033, w_000_193);
  not1 I010_160(w_010_160, w_008_411);
  and2 I010_161(w_010_161, w_008_281, w_005_424);
  nand2 I010_162(w_010_162, w_007_261, w_009_021);
  nand2 I010_163(w_010_163, w_009_016, w_003_016);
  and2 I010_164(w_010_164, w_000_119, w_008_529);
  nand2 I010_165(w_010_165, w_000_822, w_007_425);
  or2  I010_166(w_010_166, w_008_178, w_003_130);
  nand2 I010_170(w_010_170, w_004_005, w_007_456);
  nand2 I010_171(w_010_171, w_005_410, w_008_056);
  and2 I010_176(w_010_176, w_002_138, w_008_071);
  not1 I010_177(w_010_177, w_008_147);
  nand2 I010_178(w_010_178, w_006_222, w_008_884);
  and2 I010_181(w_010_181, w_009_050, w_005_246);
  and2 I010_184(w_010_184, w_008_600, w_007_376);
  and2 I010_190(w_010_190, w_000_716, w_001_101);
  not1 I010_192(w_010_192, w_002_189);
  and2 I010_193(w_010_193, w_001_147, w_002_165);
  and2 I010_196(w_010_196, w_007_202, w_009_056);
  nand2 I010_197(w_010_197, w_009_055, w_004_029);
  nand2 I010_198(w_010_198, w_004_029, w_004_028);
  not1 I010_200(w_010_200, w_008_707);
  or2  I010_204(w_010_204, w_003_065, w_005_367);
  and2 I010_205(w_010_205, w_000_440, w_000_122);
  and2 I010_208(w_010_208, w_008_170, w_008_898);
  and2 I010_210(w_010_210, w_004_022, w_006_023);
  and2 I010_211(w_010_211, w_001_086, w_000_493);
  and2 I010_212(w_010_212, w_003_064, w_002_127);
  and2 I010_218(w_010_218, w_001_469, w_003_075);
  or2  I010_220(w_010_220, w_004_006, w_008_088);
  nand2 I010_222(w_010_222, w_000_345, w_002_277);
  and2 I010_223(w_010_223, w_004_020, w_007_253);
  or2  I010_225(w_010_225, w_006_023, w_007_014);
  or2  I010_226(w_010_226, w_003_167, w_004_008);
  nand2 I010_229(w_010_229, w_007_162, w_000_806);
  and2 I010_232(w_010_232, w_004_006, w_007_048);
  not1 I010_234(w_010_234, w_006_156);
  not1 I010_236(w_010_236, w_003_073);
  not1 I010_240(w_010_240, w_004_024);
  and2 I010_246(w_010_246, w_006_129, w_004_006);
  or2  I010_247(w_010_247, w_000_652, w_004_024);
  not1 I010_249(w_010_249, w_001_388);
  nand2 I010_251(w_010_251, w_002_243, w_009_005);
  not1 I010_253(w_010_253, w_004_022);
  or2  I010_255(w_010_255, w_000_482, w_001_717);
  or2  I010_256(w_010_256, w_004_028, w_003_111);
  and2 I010_257(w_010_257, w_008_202, w_000_592);
  not1 I010_259(w_010_259, w_003_133);
  and2 I010_260(w_010_260, w_007_004, w_004_027);
  or2  I010_261(w_010_261, w_002_133, w_000_938);
  nand2 I010_264(w_010_264, w_008_672, w_001_250);
  or2  I010_265(w_010_265, w_002_123, w_005_270);
  not1 I010_267(w_010_267, w_008_013);
  and2 I010_269(w_010_269, w_005_357, w_000_402);
  not1 I010_272(w_010_272, w_003_026);
  or2  I010_278(w_010_278, w_005_294, w_004_031);
  nand2 I010_279(w_010_279, w_007_454, w_009_008);
  not1 I010_280(w_010_280, w_004_035);
  or2  I010_281(w_010_281, w_007_269, w_009_051);
  and2 I010_294(w_010_294, w_007_185, w_008_749);
  nand2 I010_295(w_010_295, w_002_028, w_002_265);
  nand2 I010_296(w_010_296, w_004_013, w_006_017);
  or2  I010_297(w_010_297, w_001_134, w_003_076);
  not1 I010_298(w_010_298, w_002_150);
  or2  I010_302(w_010_302, w_001_206, w_002_017);
  nand2 I010_304(w_010_304, w_000_853, w_007_108);
  and2 I010_307(w_010_307, w_001_853, w_003_183);
  or2  I010_310(w_010_310, w_004_038, w_005_278);
  nand2 I010_311(w_010_311, w_007_067, w_004_031);
  nand2 I010_312(w_010_312, w_009_038, w_005_559);
  or2  I010_313(w_010_313, w_000_492, w_006_307);
  not1 I010_315(w_010_315, w_000_240);
  or2  I010_316(w_010_316, w_002_402, w_002_267);
  not1 I010_321(w_010_321, w_007_094);
  not1 I010_323(w_010_323, w_007_183);
  nand2 I010_326(w_010_326, w_007_121, w_007_127);
  nand2 I010_329(w_010_329, w_004_003, w_002_086);
  or2  I010_330(w_010_330, w_001_270, w_004_000);
  not1 I010_332(w_010_332, w_002_161);
  and2 I010_334(w_010_334, w_005_049, w_004_031);
  and2 I010_335(w_010_335, w_005_144, w_003_195);
  not1 I010_338(w_010_338, w_000_399);
  nand2 I010_339(w_010_339, w_003_214, w_001_186);
  nand2 I010_340(w_010_340, w_003_142, w_008_952);
  or2  I010_344(w_010_344, w_002_079, w_007_233);
  and2 I010_346(w_010_346, w_000_864, w_004_003);
  not1 I010_349(w_010_349, w_003_185);
  not1 I010_353(w_010_353, w_007_148);
  or2  I010_358(w_010_358, w_006_276, w_001_260);
  and2 I010_359(w_010_359, w_001_176, w_002_427);
  not1 I010_365(w_010_365, w_009_060);
  and2 I010_366(w_010_366, w_005_288, w_006_009);
  not1 I010_367(w_010_367, w_005_244);
  nand2 I010_370(w_010_370, w_008_534, w_001_880);
  nand2 I010_374(w_010_374, w_000_324, w_009_024);
  nand2 I010_376(w_010_376, w_004_008, w_009_015);
  or2  I010_377(w_010_377, w_009_039, w_002_303);
  not1 I010_378(w_010_378, w_006_237);
  not1 I010_379(w_010_379, w_005_455);
  or2  I010_381(w_010_381, w_001_243, w_006_206);
  or2  I010_385(w_010_385, w_004_022, w_000_509);
  and2 I010_387(w_010_387, w_005_040, w_008_501);
  or2  I010_388(w_010_388, w_004_019, w_002_115);
  nand2 I010_389(w_010_389, w_000_058, w_000_909);
  nand2 I010_391(w_010_391, w_003_091, w_004_031);
  and2 I010_392(w_010_392, w_007_101, w_009_045);
  and2 I010_396(w_010_396, w_002_248, w_001_085);
  or2  I010_397(w_010_397, w_001_527, w_002_339);
  nand2 I010_401(w_010_401, w_009_038, w_002_184);
  and2 I010_403(w_010_403, w_005_138, w_001_848);
  or2  I010_404(w_010_404, w_003_008, w_002_061);
  or2  I010_406(w_010_406, w_001_748, w_007_332);
  not1 I010_407(w_010_407, w_003_168);
  nand2 I010_409(w_010_409, w_001_410, w_003_011);
  nand2 I010_413(w_010_413, w_007_342, w_002_442);
  or2  I010_414(w_010_414, w_007_352, w_000_631);
  or2  I010_415(w_010_415, w_008_237, w_000_579);
  nand2 I010_416(w_010_416, w_005_168, w_007_432);
  not1 I010_417(w_010_417, w_005_100);
  not1 I010_420(w_010_420, w_003_063);
  or2  I010_424(w_010_424, w_006_038, w_009_062);
  and2 I010_426(w_010_426, w_008_168, w_009_008);
  not1 I010_430(w_010_430, w_009_005);
  nand2 I010_432(w_010_432, w_000_430, w_008_661);
  nand2 I010_436(w_010_436, w_000_238, w_009_001);
  not1 I010_438(w_010_438, w_008_401);
  nand2 I010_440(w_010_440, w_004_023, w_009_049);
  or2  I010_445(w_010_445, w_005_203, w_003_034);
  nand2 I010_446(w_010_446, w_002_402, w_007_253);
  and2 I010_448(w_010_448, w_004_009, w_003_006);
  and2 I010_449(w_010_449, w_008_574, w_008_023);
  and2 I010_450(w_010_450, w_002_066, w_005_297);
  or2  I010_452(w_010_452, w_006_008, w_001_725);
  or2  I010_453(w_010_453, w_009_004, w_003_094);
  or2  I010_456(w_010_456, w_000_803, w_008_485);
  not1 I010_459(w_010_459, w_005_194);
  not1 I010_461(w_010_461, w_003_220);
  and2 I010_463(w_010_463, w_008_926, w_008_264);
  or2  I010_465(w_010_465, w_004_004, w_007_248);
  nand2 I010_466(w_010_466, w_008_021, w_001_133);
  or2  I010_467(w_010_467, w_008_450, w_000_453);
  and2 I010_468(w_010_468, w_005_129, w_003_018);
  or2  I010_473(w_010_473, w_009_068, w_004_011);
  not1 I010_474(w_010_474, w_004_007);
  and2 I010_475(w_010_475, w_009_059, w_006_157);
  nand2 I010_479(w_010_479, w_005_355, w_008_241);
  nand2 I010_480(w_010_480, w_007_310, w_005_302);
  and2 I010_484(w_010_484, w_001_665, w_005_119);
  and2 I010_486(w_010_486, w_002_302, w_000_299);
  or2  I010_488(w_010_488, w_006_321, w_005_188);
  and2 I010_491(w_010_491, w_002_032, w_008_026);
  or2  I010_492(w_010_492, w_008_088, w_007_188);
  or2  I010_494(w_010_494, w_009_045, w_004_033);
  nand2 I010_499(w_010_499, w_009_022, w_001_692);
  or2  I010_501(w_010_501, w_002_267, w_008_793);
  and2 I010_504(w_010_504, w_003_161, w_001_342);
  nand2 I010_506(w_010_506, w_007_264, w_004_036);
  not1 I010_507(w_010_507, w_004_036);
  or2  I010_511(w_010_511, w_003_088, w_000_186);
  nand2 I010_514(w_010_514, w_006_244, w_009_024);
  not1 I010_518(w_010_518, w_004_019);
  or2  I010_519(w_010_519, w_004_018, w_001_410);
  or2  I010_520(w_010_520, w_004_028, w_008_271);
  not1 I010_522(w_010_522, w_006_214);
  and2 I010_523(w_010_523, w_006_307, w_006_191);
  not1 I010_525(w_010_525, w_002_143);
  not1 I010_526(w_010_526, w_005_418);
  and2 I010_528(w_010_528, w_004_017, w_003_092);
  or2  I010_530(w_010_530, w_007_039, w_003_110);
  and2 I010_531(w_010_531, w_008_227, w_006_109);
  nand2 I010_536(w_010_536, w_008_910, w_004_007);
  and2 I010_539(w_010_539, w_009_029, w_000_684);
  nand2 I010_540(w_010_540, w_001_500, w_008_943);
  or2  I010_542(w_010_542, w_009_044, w_003_069);
  not1 I010_543(w_010_543, w_005_302);
  and2 I010_547(w_010_547, w_003_041, w_002_069);
  or2  I010_548(w_010_548, w_007_358, w_003_205);
  nand2 I010_549(w_010_549, w_003_046, w_004_000);
  nand2 I010_550(w_010_550, w_009_030, w_005_074);
  not1 I010_551(w_010_551, w_003_118);
  not1 I010_557(w_010_557, w_003_197);
  not1 I010_562(w_010_562, w_006_091);
  not1 I010_565(w_010_565, w_008_237);
  and2 I010_567(w_010_567, w_007_043, w_002_026);
  nand2 I010_570(w_010_570, w_008_289, w_002_412);
  and2 I010_571(w_010_571, w_003_102, w_002_476);
  not1 I010_573(w_010_573, w_001_305);
  or2  I010_575(w_010_575, w_009_005, w_000_553);
  nand2 I010_576(w_010_576, w_006_023, w_003_208);
  not1 I010_579(w_010_579, w_002_397);
  and2 I010_580(w_010_580, w_005_200, w_009_039);
  not1 I010_583(w_010_583, w_003_052);
  and2 I010_586(w_010_586, w_005_403, w_004_034);
  and2 I010_588(w_010_588, w_007_186, w_001_861);
  not1 I010_590(w_010_590, w_005_293);
  or2  I010_591(w_010_591, w_009_067, w_008_025);
  not1 I010_592(w_010_592, w_009_017);
  and2 I010_595(w_010_595, w_005_425, w_000_553);
  nand2 I010_596(w_010_596, w_003_064, w_004_035);
  not1 I010_597(w_010_597, w_006_317);
  nand2 I010_598(w_010_598, w_009_051, w_002_167);
  not1 I010_599(w_010_599, w_000_267);
  or2  I010_601(w_010_601, w_001_813, w_005_238);
  and2 I010_606(w_010_606, w_008_133, w_000_093);
  not1 I010_607(w_010_607, w_007_165);
  nand2 I010_609(w_010_609, w_003_208, w_005_537);
  or2  I010_612(w_010_612, w_005_371, w_003_047);
  and2 I010_613(w_010_613, w_003_041, w_006_244);
  and2 I010_614(w_010_614, w_003_084, w_006_009);
  nand2 I010_615(w_010_615, w_003_198, w_009_051);
  and2 I010_618(w_010_618, w_006_207, w_001_559);
  or2  I010_622(w_010_622, w_007_393, w_009_001);
  nand2 I010_623(w_010_623, w_008_735, w_006_294);
  and2 I010_624(w_010_624, w_006_306, w_003_211);
  or2  I010_626(w_010_626, w_001_564, w_006_159);
  and2 I010_627(w_010_627, w_008_864, w_005_001);
  nand2 I010_628(w_010_628, w_000_826, w_005_417);
  not1 I010_632(w_010_632, w_006_015);
  not1 I010_633(w_010_633, w_006_016);
  not1 I010_637(w_010_637, w_006_182);
  and2 I010_640(w_010_640, w_008_354, w_004_020);
  and2 I010_641(w_010_641, w_006_138, w_008_021);
  or2  I010_642(w_010_642, w_007_353, w_008_242);
  not1 I010_643(w_010_643, w_009_034);
  and2 I010_645(w_010_645, w_001_794, w_009_008);
  or2  I010_646(w_010_646, w_004_036, w_005_288);
  nand2 I010_649(w_010_649, w_009_066, w_004_037);
  or2  I010_650(w_010_650, w_005_428, w_004_014);
  not1 I010_652(w_010_652, w_001_507);
  or2  I010_653(w_010_653, w_005_204, w_006_074);
  not1 I010_654(w_010_654, w_001_519);
  not1 I010_657(w_010_657, w_005_106);
  not1 I010_659(w_010_659, w_000_438);
  and2 I010_665(w_010_665, w_000_579, w_004_037);
  or2  I010_667(w_010_667, w_001_503, w_004_008);
  or2  I010_670(w_010_670, w_006_094, w_003_022);
  or2  I010_680(w_010_680, w_006_147, w_001_184);
  or2  I010_683(w_010_683, w_008_857, w_001_805);
  nand2 I010_685(w_010_685, w_003_089, w_008_314);
  or2  I010_688(w_010_688, w_004_000, w_002_452);
  nand2 I010_689(w_010_689, w_005_232, w_003_210);
  not1 I010_693(w_010_693, w_006_327);
  and2 I010_694(w_010_694, w_004_034, w_009_042);
  nand2 I010_697(w_010_697, w_005_327, w_008_727);
  and2 I010_698(w_010_698, w_007_385, w_006_208);
  not1 I010_699(w_010_699, w_008_348);
  nand2 I010_703(w_010_703, w_008_028, w_008_023);
  or2  I010_706(w_010_706, w_002_179, w_001_470);
  or2  I010_707(w_010_707, w_000_816, w_003_087);
  nand2 I010_708(w_010_708, w_005_203, w_009_050);
  or2  I010_712(w_010_712, w_002_297, w_007_254);
  nand2 I010_714(w_010_714, w_000_245, w_008_090);
  and2 I010_715(w_010_715, w_005_293, w_009_052);
  nand2 I010_716(w_010_716, w_009_032, w_007_448);
  or2  I010_717(w_010_717, w_005_323, w_003_031);
  or2  I010_718(w_010_718, w_004_001, w_007_556);
  or2  I010_719(w_010_719, w_006_163, w_006_273);
  and2 I010_729(w_010_729, w_005_217, w_000_244);
  and2 I010_730(w_010_730, w_006_158, w_003_224);
  and2 I010_734(w_010_734, w_004_016, w_008_734);
  nand2 I010_736(w_010_736, w_006_287, w_006_071);
  not1 I010_738(w_010_738, w_008_889);
  nand2 I010_740(w_010_740, w_006_255, w_005_471);
  nand2 I010_741(w_010_741, w_005_205, w_000_020);
  not1 I010_744(w_010_744, w_008_477);
  not1 I010_746(w_010_746, w_009_059);
  or2  I010_747(w_010_747, w_005_073, w_009_011);
  or2  I010_749(w_010_749, w_002_423, w_006_150);
  or2  I010_751(w_010_751, w_001_239, w_009_002);
  nand2 I010_754(w_010_754, w_001_506, w_008_365);
  nand2 I010_756(w_010_756, w_003_026, w_007_335);
  or2  I010_757(w_010_757, w_002_159, w_004_003);
  and2 I010_760(w_010_760, w_009_012, w_006_327);
  or2  I010_766(w_010_766, w_009_027, w_004_032);
  and2 I010_767(w_010_767, w_004_018, w_002_016);
  and2 I010_768(w_010_768, w_008_892, w_009_025);
  and2 I010_771(w_010_771, w_003_007, w_001_645);
  or2  I010_772(w_010_772, w_006_050, w_006_102);
  nand2 I010_773(w_010_773, w_000_943, w_007_364);
  not1 I010_776(w_010_776, w_009_006);
  and2 I010_777(w_010_777, w_003_214, w_004_015);
  or2  I010_779(w_010_779, w_002_182, w_000_343);
  or2  I010_780(w_010_780, w_007_267, w_000_019);
  not1 I010_781(w_010_781, w_007_000);
  and2 I010_785(w_010_785, w_005_038, w_007_331);
  nand2 I010_790(w_010_790, w_009_004, w_007_110);
  nand2 I010_793(w_010_793, w_002_074, w_009_003);
  nand2 I010_795(w_010_795, w_006_003, w_000_142);
  or2  I010_798(w_010_798, w_008_261, w_003_065);
  not1 I010_802(w_010_802, w_002_312);
  and2 I010_804(w_010_804, w_002_496, w_000_060);
  and2 I010_805(w_010_805, w_000_673, w_001_327);
  or2  I010_806(w_010_806, w_004_009, w_003_024);
  and2 I010_807(w_010_807, w_003_035, w_000_354);
  and2 I010_809(w_010_809, w_002_114, w_009_047);
  or2  I010_810(w_010_810, w_007_139, w_007_417);
  nand2 I010_812(w_010_812, w_007_345, w_006_029);
  not1 I010_813(w_010_813, w_004_028);
  and2 I010_815(w_010_815, w_005_532, w_006_042);
  nand2 I010_817(w_010_817, w_002_385, w_009_042);
  nand2 I010_819(w_010_819, w_003_171, w_007_268);
  or2  I010_820(w_010_820, w_001_765, w_006_282);
  or2  I010_821(w_010_821, w_002_328, w_005_137);
  or2  I010_822(w_010_822, w_001_197, w_001_218);
  not1 I010_825(w_010_825, w_006_241);
  not1 I010_827(w_010_827, w_002_107);
  not1 I010_831(w_010_831, w_001_099);
  or2  I010_833(w_010_833, w_007_433, w_009_001);
  nand2 I010_834(w_010_834, w_006_169, w_001_087);
  or2  I011_000(w_011_000, w_005_099, w_007_491);
  not1 I011_001(w_011_001, w_006_167);
  or2  I011_003(w_011_003, w_002_358, w_003_042);
  nand2 I011_004(w_011_004, w_007_151, w_010_166);
  and2 I011_006(w_011_006, w_003_118, w_004_020);
  nand2 I011_007(w_011_007, w_010_330, w_003_034);
  not1 I011_008(w_011_008, w_001_497);
  not1 I011_009(w_011_009, w_003_174);
  and2 I011_010(w_011_010, w_005_483, w_004_025);
  not1 I011_011(w_011_011, w_009_051);
  not1 I011_013(w_011_013, w_008_681);
  not1 I011_014(w_011_014, w_003_049);
  nand2 I011_016(w_011_016, w_007_095, w_003_114);
  not1 I011_017(w_011_017, w_009_050);
  nand2 I011_018(w_011_018, w_008_446, w_003_014);
  and2 I011_020(w_011_020, w_004_004, w_001_411);
  nand2 I011_022(w_011_022, w_001_861, w_004_030);
  and2 I011_023(w_011_023, w_000_895, w_001_046);
  or2  I011_025(w_011_025, w_007_033, w_001_534);
  nand2 I011_026(w_011_026, w_009_020, w_008_409);
  nand2 I011_029(w_011_029, w_007_053, w_002_462);
  and2 I011_030(w_011_030, w_001_358, w_008_077);
  and2 I011_031(w_011_031, w_006_038, w_008_300);
  or2  I011_032(w_011_032, w_006_263, w_006_213);
  or2  I011_033(w_011_033, w_005_119, w_008_188);
  nand2 I011_034(w_011_034, w_004_024, w_006_141);
  nand2 I011_037(w_011_037, w_006_267, w_000_691);
  or2  I011_039(w_011_039, w_001_672, w_000_331);
  and2 I011_040(w_011_040, w_005_322, w_004_024);
  not1 I011_041(w_011_041, w_001_293);
  not1 I011_042(w_011_042, w_010_806);
  or2  I011_043(w_011_043, w_004_006, w_009_010);
  nand2 I011_044(w_011_044, w_002_182, w_006_020);
  and2 I011_045(w_011_045, w_005_173, w_009_027);
  not1 I011_046(w_011_046, w_008_534);
  not1 I011_047(w_011_047, w_007_186);
  or2  I011_049(w_011_049, w_002_305, w_004_014);
  and2 I011_050(w_011_050, w_007_386, w_004_017);
  and2 I011_053(w_011_053, w_004_006, w_009_005);
  and2 I011_056(w_011_056, w_008_001, w_000_944);
  not1 I011_057(w_011_057, w_007_374);
  or2  I011_058(w_011_058, w_007_280, w_000_596);
  and2 I011_059(w_011_059, w_008_632, w_004_012);
  or2  I011_062(w_011_062, w_006_046, w_009_040);
  nand2 I011_063(w_011_063, w_009_035, w_002_264);
  and2 I011_064(w_011_064, w_005_109, w_009_065);
  or2  I011_065(w_011_065, w_004_005, w_008_325);
  or2  I011_066(w_011_066, w_008_104, w_009_063);
  nand2 I011_067(w_011_067, w_002_086, w_003_210);
  nand2 I011_068(w_011_068, w_005_019, w_008_056);
  or2  I011_069(w_011_069, w_009_063, w_000_278);
  nand2 I011_071(w_011_071, w_005_119, w_001_803);
  not1 I011_072(w_011_072, w_007_128);
  nand2 I011_075(w_011_075, w_002_004, w_006_279);
  or2  I011_078(w_011_078, w_002_462, w_006_247);
  nand2 I011_079(w_011_079, w_002_393, w_009_037);
  and2 I011_082(w_011_082, w_008_619, w_009_037);
  and2 I011_084(w_011_084, w_008_235, w_006_132);
  or2  I011_087(w_011_087, w_003_066, w_009_038);
  nand2 I011_088(w_011_088, w_005_251, w_006_183);
  not1 I011_090(w_011_090, w_000_483);
  nand2 I011_091(w_011_091, w_007_159, w_003_213);
  and2 I011_092(w_011_092, w_007_324, w_003_102);
  and2 I011_093(w_011_093, w_005_511, w_007_365);
  and2 I011_094(w_011_094, w_008_109, w_004_026);
  nand2 I011_096(w_011_096, w_009_027, w_005_303);
  nand2 I011_097(w_011_097, w_002_185, w_000_667);
  or2  I011_101(w_011_101, w_003_123, w_008_836);
  nand2 I011_102(w_011_102, w_010_140, w_007_336);
  nand2 I011_103(w_011_103, w_006_285, w_002_221);
  and2 I011_106(w_011_106, w_002_014, w_009_048);
  not1 I011_107(w_011_107, w_001_347);
  and2 I011_109(w_011_109, w_006_249, w_009_049);
  not1 I011_110(w_011_110, w_004_013);
  nand2 I011_111(w_011_111, w_008_473, w_010_184);
  not1 I011_112(w_011_112, w_007_202);
  nand2 I011_114(w_011_114, w_006_195, w_008_656);
  or2  I011_118(w_011_118, w_010_059, w_000_151);
  nand2 I011_120(w_011_120, w_006_290, w_006_319);
  not1 I011_121(w_011_121, w_001_180);
  not1 I011_122(w_011_122, w_005_176);
  and2 I011_125(w_011_125, w_002_222, w_001_514);
  not1 I011_126(w_011_126, w_000_161);
  and2 I011_127(w_011_127, w_002_184, w_003_155);
  or2  I011_129(w_011_129, w_009_048, w_009_055);
  nand2 I011_130(w_011_130, w_005_305, w_006_268);
  nand2 I011_131(w_011_131, w_010_192, w_004_020);
  not1 I011_133(w_011_133, w_003_212);
  nand2 I011_135(w_011_135, w_008_585, w_005_441);
  not1 I011_136(w_011_136, w_001_565);
  or2  I011_137(w_011_137, w_006_222, w_003_032);
  not1 I011_138(w_011_138, w_002_128);
  nand2 I011_140(w_011_140, w_003_012, w_005_416);
  and2 I011_141(w_011_141, w_010_615, w_008_651);
  not1 I011_142(w_011_142, w_005_014);
  nand2 I011_143(w_011_143, w_009_065, w_008_921);
  and2 I011_144(w_011_144, w_001_143, w_003_007);
  and2 I011_146(w_011_146, w_003_083, w_005_103);
  not1 I011_150(w_011_150, w_003_090);
  or2  I011_153(w_011_153, w_010_729, w_009_053);
  and2 I011_154(w_011_154, w_001_100, w_000_945);
  not1 I011_155(w_011_155, w_010_624);
  and2 I011_156(w_011_156, w_003_115, w_008_033);
  not1 I011_157(w_011_157, w_003_087);
  nand2 I011_158(w_011_158, w_003_210, w_006_062);
  not1 I011_159(w_011_159, w_007_426);
  and2 I011_160(w_011_160, w_009_001, w_004_019);
  or2  I011_161(w_011_161, w_005_047, w_009_035);
  or2  I011_162(w_011_162, w_002_358, w_003_046);
  and2 I011_163(w_011_163, w_006_192, w_005_058);
  not1 I011_164(w_011_164, w_007_161);
  or2  I011_167(w_011_167, w_009_053, w_008_900);
  or2  I011_168(w_011_168, w_006_311, w_000_730);
  and2 I011_170(w_011_170, w_010_164, w_009_005);
  or2  I011_171(w_011_171, w_002_260, w_006_091);
  not1 I011_172(w_011_172, w_004_005);
  nand2 I011_173(w_011_173, w_009_038, w_003_119);
  nand2 I011_175(w_011_175, w_009_039, w_002_217);
  or2  I011_176(w_011_176, w_005_246, w_002_100);
  not1 I011_177(w_011_177, w_010_526);
  nand2 I011_178(w_011_178, w_001_786, w_009_048);
  or2  I011_180(w_011_180, w_002_494, w_009_068);
  not1 I011_182(w_011_182, w_000_785);
  nand2 I011_183(w_011_183, w_003_031, w_001_195);
  nand2 I011_186(w_011_186, w_007_504, w_007_280);
  and2 I011_187(w_011_187, w_006_126, w_004_029);
  or2  I011_190(w_011_190, w_001_096, w_000_426);
  not1 I011_191(w_011_191, w_007_107);
  or2  I011_192(w_011_192, w_000_181, w_007_517);
  and2 I011_193(w_011_193, w_004_022, w_006_118);
  nand2 I011_195(w_011_195, w_006_295, w_001_884);
  nand2 I011_198(w_011_198, w_009_054, w_001_818);
  not1 I011_200(w_011_200, w_010_685);
  or2  I011_201(w_011_201, w_003_137, w_002_253);
  or2  I011_203(w_011_203, w_006_062, w_001_656);
  or2  I011_205(w_011_205, w_007_121, w_001_591);
  and2 I011_206(w_011_206, w_010_417, w_004_027);
  not1 I011_209(w_011_209, w_006_220);
  not1 I011_211(w_011_211, w_006_232);
  or2  I011_212(w_011_212, w_002_463, w_008_908);
  or2  I011_213(w_011_213, w_000_264, w_002_365);
  nand2 I011_216(w_011_216, w_006_025, w_001_783);
  or2  I011_217(w_011_217, w_009_032, w_010_140);
  not1 I011_221(w_011_221, w_002_350);
  or2  I011_222(w_011_222, w_007_349, w_010_050);
  and2 I011_223(w_011_223, w_003_145, w_001_319);
  not1 I011_224(w_011_224, w_008_669);
  not1 I011_225(w_011_225, w_010_080);
  nand2 I011_226(w_011_226, w_001_084, w_005_477);
  or2  I011_227(w_011_227, w_000_558, w_006_186);
  or2  I011_229(w_011_229, w_001_176, w_009_001);
  or2  I011_231(w_011_231, w_004_001, w_010_365);
  or2  I011_232(w_011_232, w_007_075, w_009_037);
  and2 I011_233(w_011_233, w_003_135, w_006_236);
  nand2 I011_236(w_011_236, w_010_067, w_001_878);
  and2 I011_239(w_011_239, w_009_060, w_006_096);
  not1 I011_240(w_011_240, w_002_453);
  or2  I011_241(w_011_241, w_000_119, w_001_551);
  and2 I011_242(w_011_242, w_005_139, w_010_754);
  not1 I011_243(w_011_243, w_000_947);
  and2 I011_245(w_011_245, w_003_101, w_007_306);
  and2 I011_246(w_011_246, w_000_566, w_005_036);
  not1 I011_247(w_011_247, w_008_202);
  or2  I011_250(w_011_250, w_001_335, w_000_598);
  or2  I011_251(w_011_251, w_003_166, w_006_021);
  not1 I011_253(w_011_253, w_010_776);
  or2  I011_254(w_011_254, w_003_007, w_001_493);
  and2 I011_257(w_011_257, w_003_155, w_001_010);
  or2  I011_258(w_011_258, w_005_281, w_006_004);
  nand2 I011_259(w_011_259, w_006_263, w_007_327);
  not1 I011_260(w_011_260, w_001_066);
  or2  I011_261(w_011_261, w_002_061, w_006_169);
  nand2 I011_262(w_011_262, w_009_027, w_006_171);
  not1 I011_263(w_011_263, w_009_057);
  not1 I011_264(w_011_264, w_010_335);
  nand2 I011_265(w_011_265, w_004_030, w_007_488);
  or2  I011_266(w_011_266, w_006_099, w_001_539);
  and2 I011_267(w_011_267, w_004_012, w_003_136);
  not1 I011_268(w_011_268, w_006_273);
  or2  I011_269(w_011_269, w_010_432, w_001_729);
  or2  I011_271(w_011_271, w_001_035, w_004_034);
  nand2 I011_272(w_011_272, w_000_263, w_008_191);
  not1 I011_273(w_011_273, w_009_041);
  not1 I011_274(w_011_274, w_001_328);
  and2 I011_276(w_011_276, w_002_456, w_003_098);
  or2  I011_277(w_011_277, w_004_003, w_005_074);
  or2  I011_278(w_011_278, w_006_018, w_008_015);
  or2  I011_280(w_011_280, w_005_378, w_002_232);
  not1 I011_281(w_011_281, w_010_145);
  or2  I011_282(w_011_282, w_010_654, w_001_353);
  not1 I011_283(w_011_283, w_004_014);
  not1 I011_287(w_011_287, w_000_535);
  not1 I011_288(w_011_288, w_002_145);
  and2 I011_291(w_011_291, w_010_632, w_005_396);
  or2  I011_292(w_011_292, w_000_786, w_006_122);
  or2  I011_295(w_011_295, w_004_038, w_010_459);
  or2  I011_297(w_011_297, w_004_025, w_000_762);
  and2 I011_299(w_011_299, w_009_013, w_004_033);
  and2 I011_304(w_011_304, w_008_074, w_003_153);
  or2  I011_305(w_011_305, w_003_074, w_008_033);
  and2 I011_306(w_011_306, w_007_403, w_005_227);
  or2  I011_308(w_011_308, w_009_061, w_005_392);
  nand2 I011_309(w_011_309, w_008_383, w_004_004);
  nand2 I011_310(w_011_310, w_002_250, w_010_567);
  nand2 I011_312(w_011_312, w_001_816, w_007_100);
  and2 I011_314(w_011_314, w_009_054, w_006_182);
  and2 I011_315(w_011_315, w_000_393, w_007_451);
  and2 I011_317(w_011_317, w_004_020, w_010_592);
  or2  I011_318(w_011_318, w_009_012, w_010_107);
  and2 I011_322(w_011_322, w_004_023, w_004_032);
  and2 I011_327(w_011_327, w_006_318, w_003_029);
  or2  I011_335(w_011_335, w_010_583, w_006_319);
  not1 I011_336(w_011_336, w_004_012);
  and2 I011_337(w_011_337, w_010_155, w_004_021);
  nand2 I011_339(w_011_339, w_001_069, w_004_037);
  not1 I011_340(w_011_340, w_008_006);
  nand2 I011_343(w_011_343, w_005_097, w_001_387);
  and2 I011_347(w_011_347, w_007_210, w_002_009);
  nand2 I011_349(w_011_349, w_004_034, w_008_654);
  and2 I011_351(w_011_351, w_004_030, w_001_279);
  and2 I011_353(w_011_353, w_007_404, w_003_040);
  or2  I011_355(w_011_355, w_001_119, w_009_041);
  not1 I011_356(w_011_356, w_000_240);
  nand2 I011_359(w_011_359, w_000_105, w_008_303);
  or2  I011_360(w_011_360, w_002_059, w_000_066);
  or2  I011_361(w_011_361, w_003_061, w_004_025);
  or2  I011_367(w_011_367, w_000_114, w_010_321);
  not1 I011_369(w_011_369, w_002_406);
  nand2 I011_370(w_011_370, w_010_063, w_008_269);
  not1 I011_371(w_011_371, w_005_058);
  not1 I011_372(w_011_372, w_003_047);
  or2  I011_373(w_011_373, w_001_566, w_010_014);
  not1 I011_374(w_011_374, w_010_297);
  or2  I011_376(w_011_376, w_003_017, w_006_045);
  and2 I011_380(w_011_380, w_005_191, w_004_017);
  and2 I011_387(w_011_387, w_002_185, w_010_256);
  and2 I011_394(w_011_394, w_010_599, w_000_140);
  or2  I011_395(w_011_395, w_003_036, w_000_456);
  or2  I011_396(w_011_396, w_002_302, w_007_275);
  nand2 I011_398(w_011_398, w_010_315, w_004_015);
  and2 I011_399(w_011_399, w_006_005, w_003_009);
  or2  I011_402(w_011_402, w_009_053, w_000_231);
  and2 I011_403(w_011_403, w_006_069, w_001_000);
  or2  I011_406(w_011_406, w_000_596, w_009_067);
  not1 I011_407(w_011_407, w_002_012);
  nand2 I011_409(w_011_409, w_006_176, w_006_240);
  nand2 I011_412(w_011_412, w_004_037, w_005_216);
  and2 I011_415(w_011_415, w_003_054, w_006_265);
  nand2 I011_419(w_011_419, w_009_019, w_000_228);
  not1 I011_420(w_011_420, w_003_083);
  and2 I011_422(w_011_422, w_003_131, w_007_237);
  nand2 I011_423(w_011_423, w_010_781, w_004_016);
  not1 I011_426(w_011_426, w_003_177);
  not1 I011_430(w_011_430, w_006_281);
  and2 I011_433(w_011_433, w_003_097, w_009_004);
  or2  I011_434(w_011_434, w_000_824, w_007_026);
  or2  I011_437(w_011_437, w_005_149, w_009_039);
  nand2 I011_449(w_011_449, w_009_050, w_007_142);
  not1 I011_456(w_011_456, w_002_267);
  nand2 I011_457(w_011_457, w_006_261, w_009_048);
  nand2 I011_458(w_011_458, w_004_032, w_006_016);
  or2  I011_459(w_011_459, w_002_250, w_003_175);
  not1 I011_460(w_011_460, w_005_471);
  or2  I011_463(w_011_463, w_004_013, w_007_072);
  or2  I011_464(w_011_464, w_005_472, w_000_105);
  not1 I011_467(w_011_467, w_001_312);
  and2 I011_474(w_011_474, w_002_125, w_000_289);
  nand2 I011_476(w_011_476, w_003_176, w_006_120);
  and2 I011_477(w_011_477, w_008_621, w_006_197);
  or2  I011_478(w_011_478, w_004_022, w_004_033);
  and2 I011_485(w_011_485, w_009_063, w_003_157);
  not1 I011_486(w_011_486, w_006_254);
  and2 I011_492(w_011_492, w_006_290, w_009_004);
  nand2 I011_495(w_011_495, w_001_667, w_003_043);
  nand2 I011_496(w_011_496, w_000_608, w_004_019);
  or2  I011_500(w_011_500, w_004_001, w_006_155);
  and2 I011_501(w_011_501, w_006_067, w_000_421);
  and2 I011_502(w_011_502, w_002_361, w_001_446);
  nand2 I011_503(w_011_503, w_002_243, w_005_446);
  not1 I011_504(w_011_504, w_003_137);
  not1 I011_505(w_011_505, w_008_064);
  and2 I011_510(w_011_510, w_009_020, w_000_930);
  nand2 I011_511(w_011_511, w_007_353, w_006_142);
  not1 I011_513(w_011_513, w_009_023);
  not1 I011_514(w_011_514, w_006_231);
  nand2 I011_520(w_011_520, w_005_288, w_003_086);
  nand2 I011_523(w_011_523, w_001_896, w_000_470);
  and2 I011_525(w_011_525, w_005_518, w_010_575);
  or2  I011_526(w_011_526, w_001_548, w_005_482);
  or2  I011_530(w_011_530, w_007_097, w_007_343);
  or2  I011_534(w_011_534, w_004_028, w_006_116);
  or2  I011_535(w_011_535, w_004_038, w_005_420);
  and2 I011_537(w_011_537, w_005_069, w_008_078);
  and2 I011_540(w_011_540, w_004_026, w_002_019);
  not1 I011_543(w_011_543, w_002_041);
  not1 I011_546(w_011_546, w_009_065);
  not1 I011_548(w_011_548, w_002_106);
  and2 I011_553(w_011_553, w_004_000, w_007_088);
  nand2 I011_556(w_011_556, w_004_003, w_006_014);
  nand2 I011_558(w_011_558, w_002_247, w_010_633);
  not1 I011_560(w_011_560, w_006_021);
  nand2 I011_564(w_011_564, w_000_949, w_006_201);
  and2 I011_565(w_011_565, w_004_012, w_007_135);
  or2  I011_566(w_011_566, w_009_051, w_005_419);
  and2 I011_568(w_011_568, w_002_176, w_006_178);
  and2 I011_569(w_011_569, w_001_652, w_007_267);
  or2  I011_577(w_011_577, w_005_080, w_006_256);
  not1 I011_578(w_011_578, w_000_950);
  or2  I011_581(w_011_581, w_009_040, w_003_105);
  not1 I011_583(w_011_583, w_007_360);
  nand2 I011_584(w_011_584, w_010_091, w_003_068);
  nand2 I011_587(w_011_587, w_003_160, w_003_003);
  or2  I011_596(w_011_596, w_009_002, w_004_007);
  or2  I011_601(w_011_601, w_009_055, w_008_578);
  nand2 I011_603(w_011_603, w_010_511, w_000_386);
  and2 I011_604(w_011_604, w_002_003, w_000_494);
  nand2 I011_606(w_011_606, w_004_035, w_006_137);
  and2 I011_607(w_011_607, w_004_003, w_003_176);
  nand2 I011_608(w_011_608, w_006_182, w_007_214);
  nand2 I011_610(w_011_610, w_004_018, w_002_348);
  nand2 I011_615(w_011_615, w_001_868, w_008_790);
  not1 I011_618(w_011_618, w_008_884);
  nand2 I011_619(w_011_619, w_005_030, w_003_215);
  and2 I011_622(w_011_622, w_010_637, w_009_059);
  not1 I011_624(w_011_624, w_005_102);
  and2 I011_628(w_011_628, w_000_466, w_000_633);
  not1 I011_631(w_011_631, w_010_085);
  or2  I011_635(w_011_635, w_007_237, w_007_127);
  and2 I011_637(w_011_637, w_004_016, w_005_176);
  nand2 I011_644(w_011_644, w_006_189, w_003_132);
  or2  I011_645(w_011_645, w_000_302, w_010_302);
  and2 I011_646(w_011_646, w_000_374, w_008_158);
  and2 I011_648(w_011_648, w_008_832, w_010_344);
  and2 I011_649(w_011_649, w_004_002, w_010_650);
  not1 I011_650(w_011_650, w_008_528);
  not1 I011_652(w_011_652, w_010_519);
  nand2 I011_655(w_011_655, w_008_947, w_006_221);
  nand2 I011_656(w_011_656, w_004_017, w_003_136);
  nand2 I011_657(w_011_657, w_001_521, w_010_087);
  and2 I011_659(w_011_659, w_003_087, w_001_796);
  and2 I011_661(w_011_661, w_010_643, w_003_103);
  and2 I011_662(w_011_662, w_007_261, w_009_063);
  or2  I011_666(w_011_666, w_007_196, w_009_043);
  nand2 I011_667(w_011_667, w_005_031, w_005_313);
  nand2 I011_669(w_011_669, w_003_136, w_002_350);
  not1 I011_673(w_011_673, w_009_057);
  or2  I011_675(w_011_675, w_004_008, w_003_009);
  and2 I011_678(w_011_678, w_003_130, w_003_210);
  and2 I011_679(w_011_679, w_003_136, w_006_126);
  not1 I012_002(w_012_002, w_007_092);
  not1 I012_003(w_012_003, w_009_055);
  nand2 I012_006(w_012_006, w_010_501, w_006_230);
  nand2 I012_007(w_012_007, w_001_663, w_008_890);
  nand2 I012_008(w_012_008, w_001_201, w_002_373);
  and2 I012_010(w_012_010, w_002_334, w_010_438);
  nand2 I012_011(w_012_011, w_011_094, w_011_211);
  and2 I012_012(w_012_012, w_002_253, w_005_262);
  nand2 I012_017(w_012_017, w_005_047, w_002_329);
  or2  I012_018(w_012_018, w_005_346, w_008_804);
  and2 I012_022(w_012_022, w_008_891, w_003_075);
  nand2 I012_023(w_012_023, w_003_037, w_002_118);
  or2  I012_025(w_012_025, w_007_030, w_007_558);
  and2 I012_026(w_012_026, w_001_854, w_008_484);
  and2 I012_027(w_012_027, w_002_116, w_007_252);
  not1 I012_028(w_012_028, w_011_540);
  or2  I012_030(w_012_030, w_010_683, w_011_322);
  nand2 I012_037(w_012_037, w_000_694, w_001_548);
  and2 I012_038(w_012_038, w_001_316, w_001_464);
  not1 I012_039(w_012_039, w_010_785);
  not1 I012_040(w_012_040, w_003_038);
  nand2 I012_042(w_012_042, w_003_108, w_001_125);
  not1 I012_043(w_012_043, w_000_086);
  not1 I012_044(w_012_044, w_011_040);
  not1 I012_045(w_012_045, w_009_060);
  and2 I012_048(w_012_048, w_011_367, w_007_319);
  or2  I012_050(w_012_050, w_004_005, w_011_351);
  nand2 I012_054(w_012_054, w_006_318, w_011_205);
  or2  I012_055(w_012_055, w_007_117, w_007_145);
  nand2 I012_056(w_012_056, w_005_545, w_003_008);
  and2 I012_057(w_012_057, w_004_023, w_001_635);
  nand2 I012_058(w_012_058, w_009_039, w_003_087);
  or2  I012_061(w_012_061, w_002_321, w_002_492);
  and2 I012_062(w_012_062, w_006_287, w_001_101);
  nand2 I012_063(w_012_063, w_010_777, w_008_343);
  nand2 I012_066(w_012_066, w_008_559, w_003_036);
  not1 I012_068(w_012_068, w_006_169);
  or2  I012_069(w_012_069, w_007_062, w_000_317);
  and2 I012_070(w_012_070, w_000_661, w_009_039);
  or2  I012_071(w_012_071, w_002_130, w_005_007);
  and2 I012_072(w_012_072, w_006_137, w_004_013);
  or2  I012_076(w_012_076, w_006_058, w_002_497);
  not1 I012_077(w_012_077, w_003_159);
  nand2 I012_080(w_012_080, w_008_447, w_009_011);
  nand2 I012_083(w_012_083, w_000_092, w_001_300);
  or2  I012_084(w_012_084, w_005_381, w_002_305);
  and2 I012_085(w_012_085, w_009_032, w_003_059);
  or2  I012_086(w_012_086, w_006_245, w_008_615);
  nand2 I012_088(w_012_088, w_011_046, w_011_000);
  nand2 I012_089(w_012_089, w_006_106, w_007_403);
  nand2 I012_091(w_012_091, w_011_566, w_003_132);
  and2 I012_092(w_012_092, w_010_222, w_009_065);
  nand2 I012_093(w_012_093, w_010_232, w_007_324);
  nand2 I012_096(w_012_096, w_011_637, w_001_559);
  and2 I012_098(w_012_098, w_003_035, w_004_029);
  or2  I012_099(w_012_099, w_001_022, w_004_000);
  not1 I012_101(w_012_101, w_000_483);
  nand2 I012_102(w_012_102, w_004_032, w_003_144);
  or2  I012_104(w_012_104, w_008_936, w_009_055);
  nand2 I012_105(w_012_105, w_005_054, w_008_919);
  or2  I012_106(w_012_106, w_005_270, w_000_032);
  not1 I012_107(w_012_107, w_001_868);
  and2 I012_108(w_012_108, w_001_704, w_008_149);
  and2 I012_109(w_012_109, w_011_190, w_008_282);
  nand2 I012_110(w_012_110, w_008_668, w_008_033);
  nand2 I012_112(w_012_112, w_000_952, w_000_925);
  or2  I012_113(w_012_113, w_000_310, w_011_217);
  not1 I012_114(w_012_114, w_007_111);
  not1 I012_115(w_012_115, w_003_172);
  nand2 I012_116(w_012_116, w_003_044, w_007_049);
  nand2 I012_117(w_012_117, w_007_277, w_003_060);
  and2 I012_121(w_012_121, w_003_137, w_006_274);
  or2  I012_124(w_012_124, w_000_191, w_008_096);
  not1 I012_126(w_012_126, w_008_714);
  nand2 I012_127(w_012_127, w_004_029, w_000_685);
  not1 I012_128(w_012_128, w_002_031);
  or2  I012_130(w_012_130, w_009_016, w_010_548);
  nand2 I012_133(w_012_133, w_007_209, w_002_049);
  and2 I012_134(w_012_134, w_002_233, w_002_056);
  not1 I012_136(w_012_136, w_004_012);
  and2 I012_137(w_012_137, w_001_082, w_010_249);
  nand2 I012_138(w_012_138, w_000_341, w_005_107);
  or2  I012_139(w_012_139, w_004_021, w_004_020);
  not1 I012_142(w_012_142, w_006_143);
  not1 I012_143(w_012_143, w_011_240);
  or2  I012_149(w_012_149, w_008_278, w_007_143);
  not1 I012_151(w_012_151, w_007_232);
  or2  I012_154(w_012_154, w_000_528, w_009_002);
  and2 I012_155(w_012_155, w_001_033, w_000_349);
  and2 I012_157(w_012_157, w_001_885, w_000_465);
  and2 I012_158(w_012_158, w_011_049, w_010_536);
  or2  I012_159(w_012_159, w_003_224, w_009_044);
  nand2 I012_161(w_012_161, w_008_828, w_009_042);
  or2  I012_162(w_012_162, w_009_064, w_000_656);
  not1 I012_163(w_012_163, w_001_189);
  and2 I012_165(w_012_165, w_005_365, w_005_166);
  or2  I012_166(w_012_166, w_002_494, w_008_188);
  nand2 I012_167(w_012_167, w_004_016, w_010_820);
  not1 I012_169(w_012_169, w_005_045);
  and2 I012_170(w_012_170, w_010_586, w_007_243);
  or2  I012_171(w_012_171, w_003_071, w_002_314);
  and2 I012_172(w_012_172, w_011_553, w_001_342);
  or2  I012_173(w_012_173, w_002_384, w_001_202);
  not1 I012_174(w_012_174, w_011_374);
  and2 I012_177(w_012_177, w_004_025, w_005_012);
  nand2 I012_178(w_012_178, w_011_399, w_008_655);
  or2  I012_179(w_012_179, w_009_004, w_002_453);
  nand2 I012_182(w_012_182, w_010_316, w_000_295);
  or2  I012_183(w_012_183, w_004_008, w_009_030);
  not1 I012_184(w_012_184, w_008_285);
  or2  I012_185(w_012_185, w_004_019, w_006_065);
  or2  I012_186(w_012_186, w_001_349, w_005_356);
  not1 I012_188(w_012_188, w_004_000);
  nand2 I012_190(w_012_190, w_010_549, w_000_953);
  nand2 I012_191(w_012_191, w_001_241, w_000_061);
  not1 I012_192(w_012_192, w_011_459);
  nand2 I012_193(w_012_193, w_000_161, w_000_596);
  not1 I012_195(w_012_195, w_011_190);
  or2  I012_197(w_012_197, w_002_147, w_005_382);
  not1 I012_199(w_012_199, w_011_607);
  or2  I012_203(w_012_203, w_004_000, w_005_265);
  nand2 I012_204(w_012_204, w_008_485, w_008_017);
  and2 I012_206(w_012_206, w_001_146, w_010_015);
  nand2 I012_207(w_012_207, w_004_019, w_003_021);
  nand2 I012_209(w_012_209, w_007_140, w_001_345);
  nand2 I012_211(w_012_211, w_006_011, w_002_140);
  not1 I012_212(w_012_212, w_002_199);
  or2  I012_216(w_012_216, w_010_707, w_000_307);
  and2 I012_217(w_012_217, w_005_064, w_004_025);
  or2  I012_218(w_012_218, w_008_038, w_011_056);
  nand2 I012_220(w_012_220, w_011_209, w_003_063);
  and2 I012_221(w_012_221, w_003_023, w_002_371);
  not1 I012_223(w_012_223, w_004_006);
  not1 I012_224(w_012_224, w_000_124);
  not1 I012_226(w_012_226, w_006_101);
  not1 I012_231(w_012_231, w_000_081);
  not1 I012_236(w_012_236, w_007_500);
  and2 I012_237(w_012_237, w_000_226, w_002_181);
  or2  I012_238(w_012_238, w_002_116, w_005_409);
  and2 I012_242(w_012_242, w_002_451, w_007_373);
  not1 I012_244(w_012_244, w_011_587);
  and2 I012_245(w_012_245, w_004_025, w_003_083);
  and2 I012_246(w_012_246, w_004_030, w_009_056);
  or2  I012_248(w_012_248, w_006_137, w_001_040);
  nand2 I012_249(w_012_249, w_008_414, w_006_042);
  and2 I012_252(w_012_252, w_009_029, w_008_770);
  and2 I012_253(w_012_253, w_007_201, w_010_094);
  not1 I012_256(w_012_256, w_007_257);
  not1 I012_257(w_012_257, w_011_282);
  nand2 I012_260(w_012_260, w_003_191, w_011_239);
  and2 I012_262(w_012_262, w_010_385, w_000_543);
  and2 I012_263(w_012_263, w_007_153, w_006_203);
  and2 I012_265(w_012_265, w_000_309, w_007_026);
  nand2 I012_266(w_012_266, w_011_064, w_002_162);
  and2 I012_268(w_012_268, w_001_024, w_004_011);
  or2  I012_269(w_012_269, w_005_178, w_001_280);
  nand2 I012_270(w_012_270, w_011_154, w_011_501);
  or2  I012_271(w_012_271, w_003_014, w_010_776);
  nand2 I012_272(w_012_272, w_009_016, w_002_238);
  nand2 I012_273(w_012_273, w_009_043, w_009_019);
  or2  I012_275(w_012_275, w_003_087, w_011_492);
  and2 I012_276(w_012_276, w_011_500, w_011_666);
  and2 I012_279(w_012_279, w_001_469, w_003_046);
  nand2 I012_280(w_012_280, w_005_283, w_009_058);
  or2  I012_281(w_012_281, w_002_271, w_002_055);
  nand2 I012_284(w_012_284, w_005_117, w_007_020);
  or2  I012_287(w_012_287, w_007_119, w_002_210);
  and2 I012_288(w_012_288, w_009_056, w_010_334);
  or2  I012_289(w_012_289, w_004_030, w_006_108);
  not1 I012_290(w_012_290, w_006_211);
  not1 I012_297(w_012_297, w_000_254);
  or2  I012_299(w_012_299, w_009_063, w_003_100);
  not1 I012_300(w_012_300, w_008_102);
  nand2 I012_301(w_012_301, w_002_321, w_004_006);
  nand2 I012_303(w_012_303, w_010_296, w_010_706);
  and2 I012_304(w_012_304, w_009_044, w_009_035);
  and2 I012_306(w_012_306, w_010_821, w_008_192);
  and2 I012_307(w_012_307, w_008_294, w_007_166);
  or2  I012_308(w_012_308, w_003_131, w_004_021);
  nand2 I012_312(w_012_312, w_005_094, w_004_010);
  not1 I012_314(w_012_314, w_010_031);
  or2  I012_316(w_012_316, w_010_659, w_010_366);
  or2  I012_317(w_012_317, w_000_873, w_002_263);
  not1 I012_318(w_012_318, w_000_886);
  and2 I012_321(w_012_321, w_005_145, w_002_205);
  nand2 I012_322(w_012_322, w_003_029, w_000_770);
  and2 I012_323(w_012_323, w_010_488, w_009_015);
  not1 I012_324(w_012_324, w_003_006);
  and2 I012_325(w_012_325, w_008_344, w_001_267);
  or2  I012_327(w_012_327, w_001_279, w_006_313);
  nand2 I012_329(w_012_329, w_009_013, w_003_111);
  not1 I012_330(w_012_330, w_001_051);
  and2 I012_331(w_012_331, w_004_024, w_003_132);
  not1 I012_332(w_012_332, w_003_154);
  nand2 I012_336(w_012_336, w_004_030, w_002_261);
  not1 I012_337(w_012_337, w_008_810);
  not1 I012_338(w_012_338, w_004_031);
  not1 I012_339(w_012_339, w_011_126);
  or2  I012_341(w_012_341, w_003_051, w_002_228);
  not1 I012_343(w_012_343, w_009_061);
  not1 I012_344(w_012_344, w_009_038);
  or2  I012_345(w_012_345, w_007_337, w_008_462);
  nand2 I012_349(w_012_349, w_011_163, w_006_094);
  nand2 I012_350(w_012_350, w_010_353, w_008_633);
  and2 I012_352(w_012_352, w_009_023, w_002_349);
  or2  I012_357(w_012_357, w_004_026, w_004_032);
  and2 I012_359(w_012_359, w_005_443, w_003_146);
  or2  I012_361(w_012_361, w_004_004, w_008_931);
  nand2 I012_365(w_012_365, w_007_038, w_000_288);
  or2  I012_367(w_012_367, w_009_011, w_005_049);
  not1 I012_369(w_012_369, w_002_209);
  nand2 I012_371(w_012_371, w_002_138, w_007_053);
  not1 I012_373(w_012_373, w_002_277);
  or2  I012_374(w_012_374, w_010_037, w_007_216);
  not1 I012_375(w_012_375, w_001_653);
  nand2 I012_378(w_012_378, w_011_183, w_005_317);
  and2 I012_382(w_012_382, w_006_005, w_000_954);
  nand2 I012_383(w_012_383, w_005_305, w_006_022);
  not1 I012_384(w_012_384, w_002_036);
  not1 I012_385(w_012_385, w_011_170);
  or2  I012_387(w_012_387, w_005_436, w_010_260);
  nand2 I012_388(w_012_388, w_009_001, w_008_829);
  nand2 I012_389(w_012_389, w_003_117, w_009_043);
  or2  I012_392(w_012_392, w_000_931, w_000_367);
  or2  I012_395(w_012_395, w_000_241, w_010_809);
  or2  I012_396(w_012_396, w_005_379, w_010_815);
  and2 I012_397(w_012_397, w_002_487, w_003_015);
  nand2 I012_399(w_012_399, w_004_011, w_008_591);
  and2 I012_400(w_012_400, w_007_253, w_005_132);
  or2  I012_403(w_012_403, w_008_795, w_001_027);
  or2  I012_405(w_012_405, w_001_052, w_005_186);
  and2 I012_406(w_012_406, w_009_020, w_009_052);
  and2 I012_409(w_012_409, w_001_293, w_001_274);
  and2 I012_410(w_012_410, w_007_093, w_007_239);
  nand2 I012_411(w_012_411, w_001_528, w_008_814);
  nand2 I012_413(w_012_413, w_010_312, w_006_067);
  not1 I012_414(w_012_414, w_004_012);
  or2  I012_415(w_012_415, w_000_793, w_001_261);
  not1 I012_416(w_012_416, w_003_083);
  nand2 I012_419(w_012_419, w_002_184, w_009_018);
  not1 I012_420(w_012_420, w_000_085);
  not1 I012_422(w_012_422, w_011_212);
  nand2 I012_423(w_012_423, w_004_031, w_000_406);
  nand2 I012_424(w_012_424, w_006_327, w_010_123);
  nand2 I012_425(w_012_425, w_007_002, w_004_012);
  or2  I012_426(w_012_426, w_010_547, w_010_718);
  or2  I012_427(w_012_427, w_002_305, w_006_031);
  not1 I012_428(w_012_428, w_003_014);
  or2  I012_429(w_012_429, w_002_260, w_008_251);
  not1 I012_431(w_012_431, w_003_196);
  or2  I012_432(w_012_432, w_010_148, w_009_016);
  or2  I012_434(w_012_434, w_006_242, w_011_457);
  and2 I012_435(w_012_435, w_009_011, w_007_387);
  and2 I012_436(w_012_436, w_009_026, w_004_028);
  or2  I012_437(w_012_437, w_000_013, w_009_030);
  nand2 I012_438(w_012_438, w_000_633, w_004_025);
  not1 I012_439(w_012_439, w_002_323);
  not1 I012_441(w_012_441, w_005_461);
  not1 I012_442(w_012_442, w_002_024);
  and2 I012_446(w_012_446, w_006_014, w_006_290);
  and2 I012_447(w_012_447, w_000_226, w_005_564);
  or2  I012_451(w_012_451, w_006_247, w_004_025);
  and2 I012_453(w_012_453, w_004_018, w_000_204);
  and2 I012_456(w_012_456, w_008_242, w_011_505);
  nand2 I012_458(w_012_458, w_011_016, w_004_017);
  not1 I012_459(w_012_459, w_001_150);
  not1 I012_460(w_012_460, w_009_012);
  nand2 I012_462(w_012_462, w_003_041, w_003_187);
  not1 I012_463(w_012_463, w_000_118);
  and2 I012_465(w_012_465, w_000_513, w_006_160);
  nand2 I012_469(w_012_469, w_005_387, w_010_246);
  or2  I012_470(w_012_470, w_002_218, w_000_521);
  not1 I012_471(w_012_471, w_004_035);
  nand2 I012_472(w_012_472, w_002_251, w_007_359);
  not1 I012_474(w_012_474, w_001_770);
  nand2 I012_477(w_012_477, w_000_078, w_009_011);
  not1 I012_478(w_012_478, w_010_614);
  not1 I012_488(w_012_488, w_000_023);
  not1 I012_491(w_012_491, w_005_201);
  and2 I012_493(w_012_493, w_002_157, w_004_037);
  nand2 I012_494(w_012_494, w_011_161, w_006_237);
  or2  I012_500(w_012_500, w_001_420, w_005_103);
  and2 I012_504(w_012_504, w_002_417, w_003_094);
  and2 I012_511(w_012_511, w_002_186, w_003_030);
  nand2 I012_516(w_012_516, w_011_112, w_000_538);
  nand2 I012_519(w_012_519, w_009_032, w_008_878);
  not1 I012_523(w_012_523, w_003_011);
  not1 I012_524(w_012_524, w_009_064);
  or2  I012_525(w_012_525, w_005_270, w_007_392);
  and2 I012_531(w_012_531, w_008_553, w_006_144);
  and2 I012_533(w_012_533, w_009_057, w_007_183);
  or2  I012_535(w_012_535, w_011_103, w_005_233);
  and2 I012_538(w_012_538, w_001_093, w_007_246);
  and2 I012_539(w_012_539, w_002_397, w_000_928);
  not1 I012_543(w_012_543, w_002_485);
  or2  I012_544(w_012_544, w_007_243, w_000_300);
  or2  I012_551(w_012_551, w_002_433, w_001_771);
  or2  I013_002(w_013_002, w_011_666, w_005_010);
  not1 I013_003(w_013_003, w_004_026);
  and2 I013_004(w_013_004, w_003_115, w_007_234);
  or2  I013_005(w_013_005, w_002_358, w_007_553);
  not1 I013_006(w_013_006, w_004_006);
  nand2 I013_009(w_013_009, w_003_156, w_007_089);
  nand2 I013_010(w_013_010, w_003_091, w_002_494);
  nand2 I013_011(w_013_011, w_007_413, w_000_096);
  not1 I013_012(w_013_012, w_004_016);
  and2 I013_013(w_013_013, w_000_438, w_012_551);
  nand2 I013_014(w_013_014, w_000_955, w_005_466);
  not1 I013_016(w_013_016, w_000_388);
  or2  I013_017(w_013_017, w_005_283, w_004_000);
  nand2 I013_019(w_013_019, w_010_599, w_001_854);
  nand2 I013_020(w_013_020, w_001_644, w_004_013);
  or2  I013_022(w_013_022, w_005_353, w_012_089);
  nand2 I013_025(w_013_025, w_009_053, w_011_040);
  nand2 I013_026(w_013_026, w_012_246, w_008_704);
  not1 I013_028(w_013_028, w_008_935);
  or2  I013_029(w_013_029, w_006_104, w_009_002);
  nand2 I013_030(w_013_030, w_003_072, w_001_558);
  or2  I013_031(w_013_031, w_008_671, w_002_281);
  not1 I013_032(w_013_032, w_001_046);
  and2 I013_033(w_013_033, w_012_155, w_003_195);
  not1 I013_034(w_013_034, w_006_085);
  nand2 I013_035(w_013_035, w_005_149, w_000_743);
  not1 I013_037(w_013_037, w_011_062);
  not1 I013_039(w_013_039, w_006_160);
  not1 I013_042(w_013_042, w_000_165);
  not1 I013_044(w_013_044, w_005_196);
  and2 I013_045(w_013_045, w_007_073, w_012_524);
  not1 I013_047(w_013_047, w_010_397);
  not1 I013_048(w_013_048, w_006_094);
  nand2 I013_050(w_013_050, w_009_029, w_011_010);
  and2 I013_052(w_013_052, w_000_444, w_004_016);
  and2 I013_054(w_013_054, w_005_225, w_001_068);
  not1 I013_057(w_013_057, w_009_001);
  not1 I013_058(w_013_058, w_007_175);
  nand2 I013_060(w_013_060, w_011_127, w_010_420);
  or2  I013_064(w_013_064, w_003_014, w_009_057);
  not1 I013_065(w_013_065, w_005_067);
  not1 I013_067(w_013_067, w_000_112);
  not1 I013_073(w_013_073, w_002_189);
  or2  I013_074(w_013_074, w_007_495, w_006_327);
  not1 I013_075(w_013_075, w_001_141);
  nand2 I013_077(w_013_077, w_012_199, w_012_011);
  and2 I013_078(w_013_078, w_000_929, w_005_256);
  or2  I013_079(w_013_079, w_003_046, w_006_167);
  and2 I013_080(w_013_080, w_011_187, w_009_009);
  not1 I013_081(w_013_081, w_004_018);
  or2  I013_086(w_013_086, w_007_264, w_006_241);
  nand2 I013_090(w_013_090, w_005_277, w_010_005);
  not1 I013_096(w_013_096, w_002_469);
  not1 I013_097(w_013_097, w_004_001);
  not1 I013_098(w_013_098, w_006_319);
  and2 I013_099(w_013_099, w_002_206, w_008_568);
  not1 I013_100(w_013_100, w_010_810);
  and2 I013_102(w_013_102, w_000_425, w_000_238);
  or2  I013_104(w_013_104, w_007_349, w_008_340);
  not1 I013_105(w_013_105, w_004_008);
  nand2 I013_106(w_013_106, w_010_279, w_002_066);
  not1 I013_107(w_013_107, w_007_460);
  not1 I013_108(w_013_108, w_009_011);
  not1 I013_112(w_013_112, w_004_024);
  and2 I013_114(w_013_114, w_005_094, w_011_525);
  and2 I013_116(w_013_116, w_005_308, w_003_170);
  or2  I013_119(w_013_119, w_003_059, w_001_031);
  nand2 I013_120(w_013_120, w_001_031, w_010_029);
  not1 I013_121(w_013_121, w_008_906);
  not1 I013_123(w_013_123, w_002_300);
  not1 I013_126(w_013_126, w_011_510);
  and2 I013_127(w_013_127, w_004_038, w_006_222);
  and2 I013_128(w_013_128, w_006_035, w_010_210);
  and2 I013_129(w_013_129, w_004_017, w_011_223);
  and2 I013_133(w_013_133, w_005_108, w_008_213);
  or2  I013_136(w_013_136, w_010_613, w_000_066);
  nand2 I013_139(w_013_139, w_000_444, w_007_415);
  or2  I013_140(w_013_140, w_001_659, w_010_023);
  or2  I013_142(w_013_142, w_009_025, w_012_383);
  not1 I013_143(w_013_143, w_001_884);
  not1 I013_146(w_013_146, w_008_257);
  or2  I013_147(w_013_147, w_001_670, w_010_609);
  and2 I013_148(w_013_148, w_010_090, w_001_259);
  or2  I013_150(w_013_150, w_007_223, w_004_000);
  not1 I013_152(w_013_152, w_006_174);
  or2  I013_154(w_013_154, w_012_516, w_003_075);
  and2 I013_157(w_013_157, w_009_024, w_002_246);
  not1 I013_158(w_013_158, w_002_137);
  or2  I013_159(w_013_159, w_003_089, w_005_287);
  nand2 I013_160(w_013_160, w_009_031, w_008_299);
  nand2 I013_161(w_013_161, w_008_815, w_002_153);
  or2  I013_164(w_013_164, w_010_157, w_006_133);
  not1 I013_165(w_013_165, w_008_386);
  not1 I013_167(w_013_167, w_008_662);
  nand2 I013_170(w_013_170, w_012_442, w_002_320);
  nand2 I013_171(w_013_171, w_001_078, w_009_009);
  not1 I013_172(w_013_172, w_006_035);
  or2  I013_174(w_013_174, w_001_777, w_002_122);
  and2 I013_175(w_013_175, w_007_422, w_008_888);
  or2  I013_176(w_013_176, w_000_686, w_002_327);
  not1 I013_177(w_013_177, w_004_016);
  not1 I013_178(w_013_178, w_003_105);
  not1 I013_180(w_013_180, w_005_232);
  and2 I013_181(w_013_181, w_005_473, w_005_407);
  nand2 I013_184(w_013_184, w_012_127, w_008_143);
  or2  I013_186(w_013_186, w_007_132, w_007_023);
  not1 I013_187(w_013_187, w_001_167);
  not1 I013_188(w_013_188, w_009_020);
  not1 I013_189(w_013_189, w_006_188);
  not1 I013_191(w_013_191, w_000_260);
  nand2 I013_192(w_013_192, w_006_059, w_007_293);
  nand2 I013_194(w_013_194, w_011_163, w_000_593);
  nand2 I013_197(w_013_197, w_008_785, w_010_802);
  and2 I013_198(w_013_198, w_010_414, w_001_670);
  or2  I013_202(w_013_202, w_010_719, w_006_080);
  not1 I013_203(w_013_203, w_009_047);
  or2  I013_204(w_013_204, w_000_949, w_008_331);
  or2  I013_207(w_013_207, w_002_119, w_008_333);
  not1 I013_208(w_013_208, w_000_399);
  nand2 I013_209(w_013_209, w_011_596, w_000_891);
  or2  I013_210(w_013_210, w_002_204, w_011_399);
  nand2 I013_213(w_013_213, w_000_956, w_011_406);
  nand2 I013_219(w_013_219, w_001_074, w_000_300);
  nand2 I013_220(w_013_220, w_000_706, w_008_720);
  or2  I013_223(w_013_223, w_004_031, w_011_500);
  nand2 I013_224(w_013_224, w_012_428, w_002_416);
  and2 I013_228(w_013_228, w_006_166, w_012_260);
  nand2 I013_233(w_013_233, w_006_177, w_003_053);
  not1 I013_235(w_013_235, w_008_374);
  or2  I013_237(w_013_237, w_012_337, w_008_069);
  and2 I013_238(w_013_238, w_005_545, w_011_335);
  nand2 I013_239(w_013_239, w_000_894, w_008_814);
  or2  I013_240(w_013_240, w_000_671, w_000_476);
  or2  I013_241(w_013_241, w_002_167, w_004_021);
  nand2 I013_242(w_013_242, w_007_388, w_008_682);
  nand2 I013_243(w_013_243, w_009_064, w_011_615);
  or2  I013_244(w_013_244, w_003_084, w_004_022);
  not1 I013_249(w_013_249, w_001_694);
  nand2 I013_251(w_013_251, w_005_132, w_011_046);
  not1 I013_252(w_013_252, w_011_045);
  and2 I013_253(w_013_253, w_010_211, w_003_097);
  nand2 I013_254(w_013_254, w_009_061, w_008_599);
  or2  I013_258(w_013_258, w_009_063, w_001_686);
  not1 I013_259(w_013_259, w_001_083);
  not1 I013_260(w_013_260, w_011_646);
  or2  I013_261(w_013_261, w_008_694, w_010_039);
  or2  I013_263(w_013_263, w_006_088, w_011_403);
  not1 I013_264(w_013_264, w_002_081);
  or2  I013_265(w_013_265, w_009_037, w_005_101);
  or2  I013_267(w_013_267, w_003_041, w_002_341);
  not1 I013_268(w_013_268, w_010_387);
  nand2 I013_271(w_013_271, w_009_030, w_005_142);
  and2 I013_272(w_013_272, w_003_122, w_011_644);
  not1 I013_273(w_013_273, w_010_820);
  and2 I013_274(w_013_274, w_001_213, w_012_488);
  or2  I013_276(w_013_276, w_003_128, w_004_016);
  nand2 I013_277(w_013_277, w_002_260, w_004_012);
  not1 I013_278(w_013_278, w_011_020);
  not1 I013_279(w_013_279, w_001_501);
  and2 I013_280(w_013_280, w_000_648, w_006_202);
  and2 I013_281(w_013_281, w_009_058, w_004_008);
  and2 I013_282(w_013_282, w_002_054, w_005_342);
  or2  I013_285(w_013_285, w_006_201, w_011_091);
  nand2 I013_286(w_013_286, w_007_135, w_003_014);
  not1 I013_288(w_013_288, w_003_055);
  or2  I013_290(w_013_290, w_008_923, w_011_114);
  not1 I013_291(w_013_291, w_010_166);
  and2 I013_292(w_013_292, w_010_223, w_000_912);
  nand2 I013_297(w_013_297, w_012_477, w_003_191);
  nand2 I013_298(w_013_298, w_002_357, w_004_036);
  or2  I013_299(w_013_299, w_006_062, w_012_104);
  nand2 I013_300(w_013_300, w_011_661, w_005_102);
  and2 I013_301(w_013_301, w_010_779, w_000_384);
  and2 I013_302(w_013_302, w_005_515, w_005_394);
  or2  I013_303(w_013_303, w_010_790, w_011_269);
  and2 I013_305(w_013_305, w_007_192, w_011_495);
  nand2 I013_307(w_013_307, w_007_164, w_000_754);
  or2  I013_308(w_013_308, w_005_065, w_008_356);
  nand2 I013_309(w_013_309, w_004_003, w_011_032);
  and2 I013_310(w_013_310, w_002_070, w_004_007);
  and2 I013_311(w_013_311, w_010_232, w_005_298);
  nand2 I013_312(w_013_312, w_009_009, w_012_121);
  and2 I013_313(w_013_313, w_009_003, w_000_458);
  or2  I013_315(w_013_315, w_001_856, w_003_119);
  or2  I013_316(w_013_316, w_004_035, w_007_340);
  and2 I013_317(w_013_317, w_003_077, w_007_192);
  not1 I013_319(w_013_319, w_011_661);
  or2  I013_320(w_013_320, w_000_120, w_010_825);
  and2 I013_321(w_013_321, w_011_548, w_006_164);
  nand2 I013_324(w_013_324, w_002_423, w_003_220);
  not1 I013_325(w_013_325, w_004_006);
  or2  I013_326(w_013_326, w_005_420, w_004_037);
  nand2 I013_327(w_013_327, w_001_644, w_012_431);
  and2 I013_328(w_013_328, w_008_147, w_006_201);
  or2  I013_329(w_013_329, w_006_297, w_007_311);
  and2 I013_330(w_013_330, w_000_480, w_000_120);
  or2  I013_333(w_013_333, w_002_408, w_010_807);
  not1 I013_335(w_013_335, w_009_045);
  or2  I013_338(w_013_338, w_008_739, w_000_532);
  nand2 I013_339(w_013_339, w_011_010, w_003_117);
  or2  I013_350(w_013_350, w_005_207, w_008_033);
  and2 I013_353(w_013_353, w_004_006, w_009_014);
  or2  I013_355(w_013_355, w_011_339, w_012_414);
  and2 I013_357(w_013_357, w_009_019, w_008_015);
  nand2 I013_362(w_013_362, w_012_017, w_003_057);
  or2  I013_363(w_013_363, w_003_015, w_009_058);
  not1 I013_365(w_013_365, w_000_414);
  not1 I013_368(w_013_368, w_003_193);
  and2 I013_370(w_013_370, w_003_060, w_003_202);
  and2 I013_372(w_013_372, w_004_004, w_002_151);
  and2 I013_373(w_013_373, w_001_184, w_004_025);
  and2 I013_375(w_013_375, w_006_107, w_006_225);
  and2 I013_376(w_013_376, w_000_721, w_008_813);
  not1 I013_377(w_013_377, w_006_066);
  not1 I013_379(w_013_379, w_005_049);
  not1 I013_381(w_013_381, w_000_833);
  or2  I013_382(w_013_382, w_006_109, w_005_110);
  not1 I013_384(w_013_384, w_002_088);
  and2 I013_386(w_013_386, w_000_055, w_012_493);
  not1 I013_387(w_013_387, w_007_094);
  or2  I013_389(w_013_389, w_001_784, w_003_005);
  and2 I013_391(w_013_391, w_011_478, w_012_003);
  not1 I013_392(w_013_392, w_011_464);
  not1 I013_396(w_013_396, w_010_703);
  nand2 I013_399(w_013_399, w_010_812, w_005_202);
  or2  I013_404(w_013_404, w_001_691, w_012_465);
  not1 I013_405(w_013_405, w_002_034);
  nand2 I013_406(w_013_406, w_006_176, w_009_046);
  and2 I013_407(w_013_407, w_003_043, w_009_010);
  and2 I013_409(w_013_409, w_005_386, w_003_171);
  and2 I013_412(w_013_412, w_001_425, w_007_329);
  not1 I013_415(w_013_415, w_001_798);
  not1 I013_416(w_013_416, w_007_511);
  or2  I013_417(w_013_417, w_000_758, w_012_345);
  and2 I013_418(w_013_418, w_000_370, w_000_958);
  not1 I013_419(w_013_419, w_011_371);
  not1 I013_420(w_013_420, w_012_395);
  nand2 I013_421(w_013_421, w_007_092, w_012_397);
  or2  I013_422(w_013_422, w_005_109, w_004_006);
  and2 I013_423(w_013_423, w_007_232, w_010_080);
  or2  I013_424(w_013_424, w_012_027, w_006_170);
  and2 I013_426(w_013_426, w_011_264, w_000_550);
  or2  I013_428(w_013_428, w_003_050, w_002_226);
  not1 I013_430(w_013_430, w_012_085);
  or2  I013_431(w_013_431, w_007_265, w_011_069);
  not1 I013_433(w_013_433, w_000_267);
  not1 I013_434(w_013_434, w_009_022);
  not1 I013_437(w_013_437, w_003_108);
  not1 I013_441(w_013_441, w_001_351);
  or2  I013_442(w_013_442, w_008_672, w_006_051);
  nand2 I013_444(w_013_444, w_000_008, w_007_105);
  and2 I013_445(w_013_445, w_005_258, w_011_037);
  or2  I013_446(w_013_446, w_011_343, w_001_804);
  nand2 I013_448(w_013_448, w_003_047, w_004_003);
  not1 I013_449(w_013_449, w_001_051);
  and2 I013_450(w_013_450, w_011_622, w_011_569);
  nand2 I013_451(w_013_451, w_008_026, w_004_009);
  and2 I013_452(w_013_452, w_002_117, w_008_611);
  and2 I013_453(w_013_453, w_009_008, w_010_160);
  and2 I013_455(w_013_455, w_005_228, w_003_132);
  or2  I013_457(w_013_457, w_010_456, w_003_063);
  nand2 I013_458(w_013_458, w_012_084, w_006_197);
  nand2 I013_459(w_013_459, w_011_678, w_000_596);
  or2  I013_462(w_013_462, w_003_167, w_004_015);
  or2  I013_463(w_013_463, w_000_774, w_011_195);
  and2 I013_465(w_013_465, w_003_175, w_009_042);
  nand2 I013_466(w_013_466, w_006_227, w_004_008);
  not1 I013_469(w_013_469, w_001_771);
  and2 I013_470(w_013_470, w_001_318, w_004_000);
  or2  I013_471(w_013_471, w_009_035, w_003_189);
  and2 I013_475(w_013_475, w_001_567, w_003_087);
  not1 I013_477(w_013_477, w_009_000);
  nand2 I013_478(w_013_478, w_008_491, w_010_528);
  nand2 I013_479(w_013_479, w_011_014, w_008_959);
  or2  I013_480(w_013_480, w_002_222, w_002_375);
  nand2 I013_481(w_013_481, w_005_245, w_002_478);
  not1 I013_485(w_013_485, w_009_010);
  or2  I013_486(w_013_486, w_009_051, w_000_286);
  and2 I013_487(w_013_487, w_004_002, w_003_169);
  and2 I013_488(w_013_488, w_008_092, w_007_042);
  not1 I014_000(w_014_000, w_013_326);
  nand2 I014_006(w_014_006, w_004_031, w_011_120);
  or2  I014_008(w_014_008, w_009_030, w_005_010);
  or2  I014_010(w_014_010, w_003_024, w_003_161);
  and2 I014_013(w_014_013, w_002_015, w_009_015);
  nand2 I014_017(w_014_017, w_006_264, w_000_919);
  and2 I014_020(w_014_020, w_010_504, w_000_610);
  and2 I014_021(w_014_021, w_011_628, w_005_314);
  not1 I014_024(w_014_024, w_006_282);
  not1 I014_025(w_014_025, w_000_683);
  not1 I014_026(w_014_026, w_008_955);
  not1 I014_030(w_014_030, w_004_037);
  or2  I014_031(w_014_031, w_008_545, w_000_937);
  nand2 I014_032(w_014_032, w_009_025, w_003_025);
  nand2 I014_033(w_014_033, w_001_803, w_005_090);
  nand2 I014_034(w_014_034, w_004_027, w_005_315);
  not1 I014_035(w_014_035, w_010_379);
  or2  I014_036(w_014_036, w_001_406, w_010_359);
  nand2 I014_039(w_014_039, w_011_065, w_013_368);
  and2 I014_040(w_014_040, w_004_016, w_012_436);
  or2  I014_042(w_014_042, w_011_387, w_004_003);
  or2  I014_043(w_014_043, w_013_338, w_001_010);
  and2 I014_046(w_014_046, w_010_416, w_007_050);
  and2 I014_051(w_014_051, w_003_191, w_006_234);
  and2 I014_052(w_014_052, w_001_107, w_013_243);
  nand2 I014_053(w_014_053, w_004_034, w_012_287);
  nand2 I014_054(w_014_054, w_013_165, w_009_020);
  or2  I014_055(w_014_055, w_010_120, w_010_111);
  or2  I014_056(w_014_056, w_008_348, w_004_014);
  nand2 I014_057(w_014_057, w_011_501, w_008_053);
  or2  I014_058(w_014_058, w_008_100, w_005_485);
  not1 I014_060(w_014_060, w_011_433);
  and2 I014_061(w_014_061, w_005_299, w_003_049);
  and2 I014_063(w_014_063, w_005_444, w_011_610);
  or2  I014_064(w_014_064, w_005_088, w_010_114);
  not1 I014_069(w_014_069, w_001_824);
  not1 I014_070(w_014_070, w_005_268);
  or2  I014_071(w_014_071, w_007_005, w_008_885);
  nand2 I014_072(w_014_072, w_006_000, w_001_725);
  nand2 I014_073(w_014_073, w_005_569, w_011_373);
  nand2 I014_076(w_014_076, w_000_122, w_006_056);
  nand2 I014_078(w_014_078, w_002_349, w_010_132);
  not1 I014_080(w_014_080, w_000_646);
  nand2 I014_085(w_014_085, w_004_002, w_013_299);
  or2  I014_086(w_014_086, w_000_220, w_004_006);
  not1 I014_087(w_014_087, w_011_114);
  or2  I014_088(w_014_088, w_007_157, w_009_011);
  nand2 I014_091(w_014_091, w_001_405, w_010_349);
  not1 I014_092(w_014_092, w_009_000);
  nand2 I014_093(w_014_093, w_007_220, w_011_314);
  and2 I014_095(w_014_095, w_000_937, w_013_139);
  or2  I014_097(w_014_097, w_007_187, w_006_314);
  nand2 I014_098(w_014_098, w_003_178, w_006_327);
  or2  I014_099(w_014_099, w_009_033, w_004_005);
  or2  I014_101(w_014_101, w_002_416, w_000_960);
  or2  I014_104(w_014_104, w_006_171, w_013_328);
  and2 I014_109(w_014_109, w_013_424, w_000_357);
  or2  I014_111(w_014_111, w_003_065, w_006_165);
  or2  I014_115(w_014_115, w_013_029, w_001_807);
  nand2 I014_116(w_014_116, w_009_048, w_007_122);
  not1 I014_119(w_014_119, w_009_048);
  not1 I014_123(w_014_123, w_006_008);
  nand2 I014_124(w_014_124, w_006_277, w_009_036);
  and2 I014_125(w_014_125, w_008_756, w_008_034);
  or2  I014_127(w_014_127, w_010_204, w_006_021);
  and2 I014_128(w_014_128, w_010_313, w_008_747);
  nand2 I014_130(w_014_130, w_012_186, w_005_474);
  or2  I014_131(w_014_131, w_010_751, w_010_637);
  or2  I014_135(w_014_135, w_010_047, w_011_058);
  not1 I014_136(w_014_136, w_011_177);
  and2 I014_137(w_014_137, w_000_332, w_001_602);
  or2  I014_139(w_014_139, w_006_073, w_007_095);
  and2 I014_140(w_014_140, w_007_129, w_012_426);
  or2  I014_141(w_014_141, w_000_726, w_004_001);
  or2  I014_142(w_014_142, w_000_176, w_013_120);
  nand2 I014_143(w_014_143, w_000_721, w_001_825);
  nand2 I014_145(w_014_145, w_011_216, w_010_081);
  not1 I014_147(w_014_147, w_008_596);
  nand2 I014_150(w_014_150, w_003_158, w_001_561);
  not1 I014_152(w_014_152, w_004_019);
  and2 I014_155(w_014_155, w_007_432, w_011_243);
  or2  I014_157(w_014_157, w_001_024, w_004_002);
  or2  I014_158(w_014_158, w_003_004, w_006_165);
  not1 I014_159(w_014_159, w_008_670);
  or2  I014_160(w_014_160, w_007_501, w_005_561);
  nand2 I014_161(w_014_161, w_002_237, w_009_041);
  nand2 I014_162(w_014_162, w_000_145, w_009_003);
  nand2 I014_163(w_014_163, w_006_221, w_004_014);
  not1 I014_164(w_014_164, w_006_209);
  and2 I014_165(w_014_165, w_009_063, w_008_138);
  and2 I014_167(w_014_167, w_008_662, w_001_553);
  or2  I014_168(w_014_168, w_001_288, w_008_824);
  nand2 I014_169(w_014_169, w_007_409, w_002_122);
  and2 I014_179(w_014_179, w_007_220, w_010_267);
  nand2 I014_180(w_014_180, w_001_590, w_010_760);
  nand2 I014_181(w_014_181, w_012_163, w_007_435);
  not1 I014_183(w_014_183, w_006_287);
  not1 I014_184(w_014_184, w_005_402);
  not1 I014_186(w_014_186, w_003_134);
  and2 I014_188(w_014_188, w_001_066, w_007_081);
  nand2 I014_190(w_014_190, w_007_089, w_012_272);
  nand2 I014_191(w_014_191, w_012_218, w_004_027);
  or2  I014_192(w_014_192, w_008_585, w_013_175);
  and2 I014_198(w_014_198, w_010_424, w_005_057);
  or2  I014_201(w_014_201, w_006_182, w_002_175);
  or2  I014_210(w_014_210, w_001_094, w_004_029);
  nand2 I014_213(w_014_213, w_005_285, w_010_074);
  and2 I014_217(w_014_217, w_002_030, w_013_210);
  nand2 I014_218(w_014_218, w_013_240, w_005_093);
  and2 I014_219(w_014_219, w_004_004, w_009_053);
  not1 I014_220(w_014_220, w_004_031);
  not1 I014_221(w_014_221, w_004_003);
  and2 I014_222(w_014_222, w_011_603, w_012_352);
  and2 I014_223(w_014_223, w_009_035, w_003_225);
  or2  I014_225(w_014_225, w_013_273, w_012_037);
  not1 I014_226(w_014_226, w_005_403);
  nand2 I014_228(w_014_228, w_012_399, w_009_063);
  nand2 I014_230(w_014_230, w_013_376, w_000_032);
  nand2 I014_235(w_014_235, w_006_284, w_010_171);
  or2  I014_236(w_014_236, w_011_523, w_002_088);
  nand2 I014_237(w_014_237, w_000_473, w_002_162);
  not1 I014_240(w_014_240, w_013_160);
  or2  I014_241(w_014_241, w_008_016, w_010_607);
  or2  I014_243(w_014_243, w_009_007, w_006_056);
  or2  I014_245(w_014_245, w_006_259, w_003_126);
  nand2 I014_247(w_014_247, w_012_252, w_004_003);
  or2  I014_248(w_014_248, w_012_268, w_008_079);
  not1 I014_250(w_014_250, w_008_306);
  not1 I014_251(w_014_251, w_004_011);
  nand2 I014_252(w_014_252, w_004_025, w_003_161);
  nand2 I014_253(w_014_253, w_001_471, w_010_601);
  not1 I014_254(w_014_254, w_006_187);
  not1 I014_255(w_014_255, w_010_122);
  nand2 I014_256(w_014_256, w_006_135, w_004_007);
  and2 I014_259(w_014_259, w_006_060, w_011_608);
  or2  I014_260(w_014_260, w_012_523, w_002_136);
  or2  I014_263(w_014_263, w_002_002, w_010_190);
  and2 I014_264(w_014_264, w_007_193, w_012_331);
  nand2 I014_267(w_014_267, w_000_028, w_013_077);
  nand2 I014_268(w_014_268, w_000_736, w_006_322);
  or2  I014_269(w_014_269, w_002_216, w_013_422);
  nand2 I014_270(w_014_270, w_002_424, w_010_110);
  not1 I014_271(w_014_271, w_001_303);
  or2  I014_275(w_014_275, w_010_507, w_006_159);
  not1 I014_276(w_014_276, w_006_248);
  or2  I014_277(w_014_277, w_008_836, w_009_058);
  nand2 I014_279(w_014_279, w_008_373, w_001_219);
  not1 I014_281(w_014_281, w_009_058);
  nand2 I014_282(w_014_282, w_003_156, w_011_001);
  not1 I014_283(w_014_283, w_003_041);
  nand2 I014_285(w_014_285, w_000_570, w_008_043);
  or2  I014_286(w_014_286, w_001_416, w_000_472);
  not1 I014_287(w_014_287, w_000_925);
  not1 I014_289(w_014_289, w_005_365);
  nand2 I014_291(w_014_291, w_007_432, w_002_183);
  nand2 I014_292(w_014_292, w_002_255, w_009_062);
  not1 I014_293(w_014_293, w_010_176);
  nand2 I014_298(w_014_298, w_011_043, w_006_203);
  nand2 I014_300(w_014_300, w_005_270, w_004_014);
  not1 I014_303(w_014_303, w_011_523);
  nand2 I014_305(w_014_305, w_004_021, w_005_247);
  not1 I014_306(w_014_306, w_000_478);
  or2  I014_307(w_014_307, w_003_097, w_001_756);
  nand2 I014_308(w_014_308, w_006_282, w_012_312);
  not1 I014_310(w_014_310, w_000_253);
  not1 I014_311(w_014_311, w_006_237);
  and2 I014_314(w_014_314, w_009_055, w_003_058);
  not1 I014_315(w_014_315, w_010_831);
  not1 I014_320(w_014_320, w_002_314);
  nand2 I014_322(w_014_322, w_002_343, w_011_157);
  nand2 I014_323(w_014_323, w_009_046, w_003_177);
  or2  I014_324(w_014_324, w_006_039, w_007_023);
  or2  I014_325(w_014_325, w_006_158, w_000_308);
  not1 I014_329(w_014_329, w_005_132);
  or2  I014_330(w_014_330, w_012_220, w_004_028);
  nand2 I014_331(w_014_331, w_005_306, w_001_707);
  and2 I014_333(w_014_333, w_003_194, w_012_091);
  or2  I014_337(w_014_337, w_002_266, w_013_305);
  and2 I014_340(w_014_340, w_000_956, w_012_113);
  nand2 I014_341(w_014_341, w_000_383, w_007_413);
  or2  I014_344(w_014_344, w_001_513, w_011_276);
  or2  I014_345(w_014_345, w_006_324, w_005_243);
  and2 I014_346(w_014_346, w_001_838, w_001_835);
  nand2 I014_348(w_014_348, w_006_085, w_002_380);
  or2  I014_349(w_014_349, w_005_289, w_001_639);
  or2  I014_351(w_014_351, w_009_049, w_004_030);
  or2  I014_353(w_014_353, w_002_002, w_011_274);
  nand2 I014_354(w_014_354, w_006_058, w_001_586);
  nand2 I014_356(w_014_356, w_011_337, w_007_081);
  nand2 I014_357(w_014_357, w_000_120, w_007_338);
  or2  I014_359(w_014_359, w_012_076, w_001_147);
  nand2 I014_360(w_014_360, w_006_313, w_006_045);
  nand2 I014_362(w_014_362, w_013_312, w_007_182);
  not1 I014_363(w_014_363, w_002_204);
  not1 I014_365(w_014_365, w_011_514);
  or2  I014_367(w_014_367, w_000_457, w_002_012);
  or2  I014_375(w_014_375, w_001_586, w_006_256);
  not1 I014_380(w_014_380, w_010_165);
  not1 I014_383(w_014_383, w_010_646);
  nand2 I014_389(w_014_389, w_011_631, w_006_195);
  and2 I014_392(w_014_392, w_004_013, w_002_303);
  not1 I014_399(w_014_399, w_013_213);
  nand2 I014_401(w_014_401, w_004_014, w_000_538);
  or2  I014_403(w_014_403, w_004_020, w_011_170);
  nand2 I014_405(w_014_405, w_008_631, w_013_233);
  and2 I014_409(w_014_409, w_013_081, w_003_059);
  nand2 I014_411(w_014_411, w_013_389, w_003_049);
  not1 I014_415(w_014_415, w_007_347);
  nand2 I014_417(w_014_417, w_008_703, w_011_201);
  and2 I014_420(w_014_420, w_012_299, w_006_291);
  not1 I014_424(w_014_424, w_010_693);
  and2 I014_426(w_014_426, w_008_925, w_001_078);
  or2  I014_434(w_014_434, w_009_027, w_000_390);
  nand2 I014_435(w_014_435, w_004_009, w_002_406);
  or2  I014_437(w_014_437, w_010_338, w_004_012);
  and2 I014_442(w_014_442, w_005_226, w_012_179);
  and2 I014_443(w_014_443, w_006_237, w_000_194);
  nand2 I014_444(w_014_444, w_004_011, w_003_117);
  not1 I014_446(w_014_446, w_005_524);
  and2 I014_449(w_014_449, w_012_470, w_007_272);
  not1 I014_451(w_014_451, w_003_022);
  nand2 I014_453(w_014_453, w_001_280, w_000_551);
  nand2 I014_457(w_014_457, w_005_307, w_002_091);
  and2 I014_464(w_014_464, w_002_493, w_005_129);
  not1 I014_465(w_014_465, w_008_234);
  or2  I014_469(w_014_469, w_005_154, w_001_828);
  nand2 I014_470(w_014_470, w_010_834, w_013_074);
  and2 I014_472(w_014_472, w_010_623, w_006_316);
  or2  I014_474(w_014_474, w_012_089, w_000_959);
  and2 I014_479(w_014_479, w_008_396, w_006_132);
  not1 I014_482(w_014_482, w_013_184);
  not1 I014_485(w_014_485, w_008_122);
  and2 I014_487(w_014_487, w_001_794, w_012_006);
  and2 I014_500(w_014_500, w_004_001, w_004_006);
  or2  I014_503(w_014_503, w_013_471, w_009_010);
  or2  I014_504(w_014_504, w_004_001, w_013_488);
  not1 I014_507(w_014_507, w_008_897);
  and2 I014_509(w_014_509, w_008_560, w_003_221);
  not1 I014_515(w_014_515, w_003_050);
  nand2 I014_516(w_014_516, w_011_288, w_004_029);
  not1 I014_518(w_014_518, w_013_057);
  and2 I014_520(w_014_520, w_006_308, w_000_377);
  or2  I014_524(w_014_524, w_002_280, w_010_358);
  and2 I014_527(w_014_527, w_003_133, w_004_012);
  not1 I014_529(w_014_529, w_001_578);
  nand2 I014_533(w_014_533, w_005_216, w_000_062);
  and2 I014_534(w_014_534, w_001_547, w_012_171);
  nand2 I014_538(w_014_538, w_005_244, w_012_337);
  not1 I014_540(w_014_540, w_006_148);
  nand2 I014_542(w_014_542, w_010_579, w_000_124);
  nand2 I014_543(w_014_543, w_002_048, w_004_018);
  nand2 I014_545(w_014_545, w_007_512, w_012_273);
  and2 I014_546(w_014_546, w_010_006, w_005_433);
  or2  I014_549(w_014_549, w_007_260, w_008_943);
  not1 I014_554(w_014_554, w_002_334);
  and2 I014_557(w_014_557, w_007_069, w_005_216);
  and2 I014_559(w_014_559, w_010_392, w_007_018);
  or2  I014_560(w_014_560, w_001_495, w_007_055);
  nand2 I014_564(w_014_564, w_010_445, w_006_162);
  not1 I014_566(w_014_566, w_001_496);
  and2 I014_568(w_014_568, w_000_945, w_000_082);
  and2 I014_571(w_014_571, w_012_424, w_004_038);
  or2  I014_573(w_014_573, w_008_520, w_008_888);
  or2  I014_574(w_014_574, w_007_091, w_004_023);
  nand2 I014_576(w_014_576, w_010_073, w_013_004);
  nand2 I014_577(w_014_577, w_012_472, w_011_312);
  or2  I014_582(w_014_582, w_008_001, w_002_365);
  not1 I014_584(w_014_584, w_000_112);
  not1 I014_586(w_014_586, w_011_277);
  nand2 I014_594(w_014_594, w_006_195, w_002_493);
  or2  I014_595(w_014_595, w_005_201, w_005_184);
  or2  I014_598(w_014_598, w_000_963, w_003_040);
  nand2 I014_602(w_014_602, w_004_008, w_002_379);
  not1 I014_603(w_014_603, w_002_168);
  and2 I014_608(w_014_608, w_013_106, w_007_101);
  nand2 I014_609(w_014_609, w_008_480, w_009_004);
  not1 I014_613(w_014_613, w_003_030);
  and2 I014_626(w_014_626, w_010_499, w_007_392);
  or2  I014_629(w_014_629, w_000_943, w_009_005);
  nand2 I014_632(w_014_632, w_005_190, w_013_444);
  nand2 I014_634(w_014_634, w_012_271, w_001_859);
  and2 I014_635(w_014_635, w_000_844, w_009_028);
  nand2 I014_636(w_014_636, w_002_226, w_006_104);
  not1 I014_637(w_014_637, w_013_116);
  or2  I015_000(w_015_000, w_001_817, w_001_075);
  and2 I015_001(w_015_001, w_002_402, w_005_117);
  or2  I015_002(w_015_002, w_003_030, w_004_028);
  not1 I015_003(w_015_003, w_009_008);
  or2  I015_004(w_015_004, w_002_234, w_000_904);
  or2  I015_008(w_015_008, w_000_648, w_013_102);
  or2  I015_010(w_015_010, w_006_094, w_002_065);
  nand2 I015_011(w_015_011, w_002_321, w_006_041);
  and2 I015_012(w_015_012, w_006_004, w_011_164);
  not1 I015_013(w_015_013, w_008_941);
  not1 I015_015(w_015_015, w_011_265);
  and2 I015_018(w_015_018, w_001_265, w_011_376);
  or2  I015_019(w_015_019, w_002_046, w_007_539);
  or2  I015_021(w_015_021, w_004_018, w_014_417);
  not1 I015_024(w_015_024, w_007_076);
  nand2 I015_025(w_015_025, w_003_138, w_014_507);
  not1 I015_026(w_015_026, w_006_046);
  nand2 I015_027(w_015_027, w_006_212, w_014_307);
  nand2 I015_029(w_015_029, w_013_174, w_011_029);
  or2  I015_031(w_015_031, w_012_089, w_005_102);
  or2  I015_032(w_015_032, w_005_035, w_011_287);
  not1 I015_035(w_015_035, w_008_169);
  or2  I015_036(w_015_036, w_011_198, w_004_003);
  or2  I015_037(w_015_037, w_001_196, w_013_409);
  and2 I015_041(w_015_041, w_012_410, w_013_242);
  nand2 I015_042(w_015_042, w_013_365, w_007_329);
  not1 I015_043(w_015_043, w_003_120);
  not1 I015_044(w_015_044, w_001_881);
  and2 I015_045(w_015_045, w_011_064, w_002_429);
  and2 I015_047(w_015_047, w_003_165, w_013_480);
  nand2 I015_048(w_015_048, w_005_402, w_007_448);
  and2 I015_049(w_015_049, w_011_250, w_000_105);
  not1 I015_051(w_015_051, w_014_435);
  not1 I015_052(w_015_052, w_011_180);
  or2  I015_053(w_015_053, w_008_398, w_009_023);
  and2 I015_057(w_015_057, w_002_111, w_011_419);
  nand2 I015_058(w_015_058, w_000_325, w_004_017);
  nand2 I015_059(w_015_059, w_000_470, w_003_172);
  nand2 I015_061(w_015_061, w_000_566, w_001_014);
  not1 I015_062(w_015_062, w_001_228);
  and2 I015_064(w_015_064, w_002_034, w_003_044);
  not1 I015_067(w_015_067, w_010_234);
  and2 I015_071(w_015_071, w_002_246, w_009_026);
  and2 I015_072(w_015_072, w_008_712, w_005_324);
  not1 I015_078(w_015_078, w_010_385);
  not1 I015_079(w_015_079, w_007_149);
  not1 I015_080(w_015_080, w_008_025);
  not1 I015_081(w_015_081, w_001_020);
  or2  I015_083(w_015_083, w_014_362, w_004_015);
  nand2 I015_084(w_015_084, w_007_278, w_010_780);
  nand2 I015_088(w_015_088, w_010_474, w_009_004);
  or2  I015_089(w_015_089, w_004_034, w_003_035);
  not1 I015_090(w_015_090, w_002_075);
  nand2 I015_092(w_015_092, w_010_540, w_001_890);
  not1 I015_093(w_015_093, w_014_036);
  or2  I015_094(w_015_094, w_008_200, w_003_071);
  and2 I015_095(w_015_095, w_010_082, w_008_396);
  not1 I015_096(w_015_096, w_005_413);
  and2 I015_098(w_015_098, w_012_195, w_011_206);
  nand2 I015_099(w_015_099, w_007_428, w_006_034);
  nand2 I015_101(w_015_101, w_013_106, w_013_470);
  nand2 I015_103(w_015_103, w_000_591, w_010_805);
  or2  I015_106(w_015_106, w_000_084, w_012_307);
  not1 I015_108(w_015_108, w_008_850);
  and2 I015_112(w_015_112, w_014_092, w_005_101);
  and2 I015_114(w_015_114, w_009_058, w_008_882);
  or2  I015_117(w_015_117, w_010_236, w_010_583);
  not1 I015_118(w_015_118, w_007_027);
  and2 I015_122(w_015_122, w_000_170, w_007_219);
  and2 I015_124(w_015_124, w_000_914, w_002_261);
  nand2 I015_126(w_015_126, w_014_285, w_004_001);
  and2 I015_127(w_015_127, w_006_235, w_004_012);
  nand2 I015_128(w_015_128, w_002_439, w_007_082);
  or2  I015_129(w_015_129, w_014_013, w_014_136);
  or2  I015_130(w_015_130, w_008_953, w_011_619);
  and2 I015_131(w_015_131, w_005_305, w_009_035);
  nand2 I015_134(w_015_134, w_003_145, w_009_065);
  nand2 I015_135(w_015_135, w_001_844, w_004_006);
  or2  I015_136(w_015_136, w_004_031, w_014_282);
  not1 I015_138(w_015_138, w_005_226);
  not1 I015_139(w_015_139, w_006_265);
  nand2 I015_140(w_015_140, w_003_087, w_005_291);
  not1 I015_141(w_015_141, w_001_467);
  and2 I015_142(w_015_142, w_006_082, w_010_311);
  not1 I015_143(w_015_143, w_002_160);
  and2 I015_146(w_015_146, w_014_039, w_005_059);
  not1 I015_150(w_015_150, w_011_543);
  or2  I015_151(w_015_151, w_005_129, w_006_113);
  or2  I015_154(w_015_154, w_008_061, w_014_457);
  not1 I015_155(w_015_155, w_006_055);
  not1 I015_156(w_015_156, w_004_027);
  and2 I015_157(w_015_157, w_000_070, w_003_201);
  not1 I015_158(w_015_158, w_006_067);
  nand2 I015_159(w_015_159, w_007_195, w_004_011);
  and2 I015_160(w_015_160, w_011_291, w_010_017);
  and2 I015_164(w_015_164, w_002_377, w_010_013);
  not1 I015_165(w_015_165, w_001_042);
  or2  I015_166(w_015_166, w_006_025, w_000_389);
  not1 I015_168(w_015_168, w_010_079);
  and2 I015_170(w_015_170, w_013_177, w_013_160);
  nand2 I015_171(w_015_171, w_010_178, w_003_095);
  and2 I015_172(w_015_172, w_013_271, w_007_362);
  and2 I015_173(w_015_173, w_006_078, w_005_029);
  and2 I015_175(w_015_175, w_010_813, w_001_622);
  or2  I015_178(w_015_178, w_010_374, w_012_399);
  and2 I015_180(w_015_180, w_006_084, w_009_041);
  not1 I015_187(w_015_187, w_010_475);
  nand2 I015_190(w_015_190, w_012_174, w_010_650);
  not1 I015_191(w_015_191, w_013_309);
  and2 I015_193(w_015_193, w_006_277, w_011_125);
  and2 I015_196(w_015_196, w_000_525, w_008_299);
  nand2 I015_197(w_015_197, w_010_302, w_003_197);
  not1 I015_199(w_015_199, w_000_900);
  or2  I015_201(w_015_201, w_010_645, w_002_013);
  or2  I015_205(w_015_205, w_009_027, w_008_837);
  nand2 I015_206(w_015_206, w_007_076, w_005_153);
  and2 I015_207(w_015_207, w_009_048, w_000_484);
  nand2 I015_209(w_015_209, w_013_237, w_003_048);
  not1 I015_210(w_015_210, w_008_033);
  not1 I015_211(w_015_211, w_009_001);
  and2 I015_214(w_015_214, w_009_068, w_010_003);
  and2 I015_216(w_015_216, w_004_025, w_011_618);
  and2 I015_221(w_015_221, w_014_087, w_004_000);
  nand2 I015_226(w_015_226, w_010_139, w_012_209);
  and2 I015_227(w_015_227, w_012_056, w_011_101);
  or2  I015_233(w_015_233, w_004_001, w_001_542);
  or2  I015_235(w_015_235, w_001_848, w_010_491);
  and2 I015_238(w_015_238, w_012_459, w_009_016);
  nand2 I015_254(w_015_254, w_010_095, w_001_017);
  not1 I015_255(w_015_255, w_003_145);
  or2  I015_258(w_015_258, w_010_136, w_005_089);
  not1 I015_264(w_015_264, w_006_025);
  nand2 I015_265(w_015_265, w_008_331, w_012_524);
  nand2 I015_275(w_015_275, w_010_099, w_007_131);
  or2  I015_277(w_015_277, w_001_656, w_007_128);
  not1 I015_278(w_015_278, w_001_575);
  and2 I015_280(w_015_280, w_006_167, w_003_051);
  or2  I015_282(w_015_282, w_001_892, w_011_168);
  not1 I015_284(w_015_284, w_000_965);
  not1 I015_304(w_015_304, w_002_188);
  nand2 I015_314(w_015_314, w_009_024, w_002_347);
  not1 I015_315(w_015_315, w_013_235);
  and2 I015_316(w_015_316, w_004_000, w_006_109);
  and2 I015_319(w_015_319, w_008_720, w_011_581);
  and2 I015_322(w_015_322, w_004_001, w_008_749);
  or2  I015_323(w_015_323, w_014_236, w_008_184);
  not1 I015_324(w_015_324, w_013_172);
  not1 I015_328(w_015_328, w_010_006);
  and2 I015_330(w_015_330, w_004_000, w_010_480);
  not1 I015_333(w_015_333, w_003_179);
  nand2 I015_339(w_015_339, w_007_130, w_004_019);
  not1 I015_341(w_015_341, w_003_028);
  not1 I015_345(w_015_345, w_002_117);
  not1 I015_346(w_015_346, w_004_017);
  nand2 I015_348(w_015_348, w_004_037, w_000_345);
  nand2 I015_349(w_015_349, w_010_121, w_010_557);
  not1 I015_350(w_015_350, w_001_801);
  or2  I015_359(w_015_359, w_013_034, w_002_031);
  not1 I015_363(w_015_363, w_012_316);
  nand2 I015_365(w_015_365, w_010_595, w_012_066);
  or2  I015_367(w_015_367, w_008_619, w_003_178);
  not1 I015_368(w_015_368, w_007_204);
  or2  I015_369(w_015_369, w_005_310, w_011_281);
  or2  I015_373(w_015_373, w_007_207, w_012_388);
  and2 I015_394(w_015_394, w_012_442, w_008_674);
  nand2 I015_395(w_015_395, w_003_144, w_011_026);
  not1 I015_397(w_015_397, w_014_111);
  or2  I015_404(w_015_404, w_007_317, w_005_408);
  not1 I015_406(w_015_406, w_000_444);
  not1 I015_412(w_015_412, w_004_001);
  not1 I015_418(w_015_418, w_009_035);
  and2 I015_424(w_015_424, w_004_036, w_010_689);
  not1 I015_426(w_015_426, w_006_330);
  and2 I015_427(w_015_427, w_001_438, w_014_603);
  not1 I015_429(w_015_429, w_003_030);
  or2  I015_434(w_015_434, w_001_468, w_013_379);
  nand2 I015_438(w_015_438, w_010_298, w_014_586);
  or2  I015_440(w_015_440, w_008_780, w_011_396);
  and2 I015_442(w_015_442, w_009_001, w_004_010);
  or2  I015_443(w_015_443, w_008_750, w_009_058);
  not1 I015_444(w_015_444, w_008_304);
  and2 I015_445(w_015_445, w_014_250, w_009_051);
  nand2 I015_447(w_015_447, w_009_002, w_013_105);
  or2  I015_450(w_015_450, w_000_770, w_009_022);
  or2  I015_453(w_015_453, w_002_425, w_009_036);
  and2 I015_457(w_015_457, w_012_191, w_001_278);
  and2 I015_458(w_015_458, w_010_570, w_001_173);
  or2  I015_459(w_015_459, w_009_038, w_004_004);
  and2 I015_462(w_015_462, w_007_150, w_011_474);
  and2 I015_465(w_015_465, w_014_359, w_006_040);
  nand2 I015_470(w_015_470, w_004_028, w_008_894);
  not1 I015_474(w_015_474, w_011_369);
  nand2 I015_476(w_015_476, w_003_154, w_002_329);
  nand2 I015_479(w_015_479, w_008_383, w_002_055);
  nand2 I015_482(w_015_482, w_002_140, w_008_021);
  nand2 I015_490(w_015_490, w_010_310, w_013_386);
  or2  I015_492(w_015_492, w_009_004, w_012_272);
  and2 I015_493(w_015_493, w_006_214, w_005_354);
  and2 I015_494(w_015_494, w_009_039, w_002_293);
  or2  I015_496(w_015_496, w_013_150, w_002_145);
  not1 I015_499(w_015_499, w_004_031);
  or2  I015_504(w_015_504, w_002_429, w_008_862);
  nand2 I015_510(w_015_510, w_003_133, w_012_124);
  and2 I015_512(w_015_512, w_009_057, w_009_023);
  nand2 I015_517(w_015_517, w_005_463, w_003_078);
  or2  I015_519(w_015_519, w_004_031, w_005_257);
  nand2 I015_521(w_015_521, w_014_546, w_004_030);
  and2 I015_522(w_015_522, w_001_358, w_009_006);
  or2  I015_525(w_015_525, w_014_566, w_006_320);
  nand2 I015_529(w_015_529, w_008_829, w_004_034);
  or2  I015_532(w_015_532, w_005_496, w_013_288);
  and2 I015_535(w_015_535, w_011_144, w_002_454);
  or2  I015_538(w_015_538, w_012_288, w_001_462);
  or2  I015_541(w_015_541, w_000_310, w_004_035);
  or2  I015_547(w_015_547, w_006_078, w_005_298);
  nand2 I015_554(w_015_554, w_005_272, w_002_307);
  nand2 I015_559(w_015_559, w_014_124, w_002_434);
  nand2 I015_583(w_015_583, w_001_374, w_012_169);
  and2 I015_585(w_015_585, w_008_702, w_013_317);
  not1 I015_592(w_015_592, w_011_513);
  and2 I015_594(w_015_594, w_000_967, w_002_459);
  or2  I015_595(w_015_595, w_004_019, w_014_040);
  and2 I015_597(w_015_597, w_010_499, w_011_096);
  and2 I015_600(w_015_600, w_009_061, w_006_315);
  nand2 I015_603(w_015_603, w_004_008, w_010_370);
  or2  I015_604(w_015_604, w_013_147, w_014_557);
  nand2 I015_605(w_015_605, w_008_597, w_010_744);
  and2 I015_608(w_015_608, w_013_282, w_008_581);
  or2  I015_611(w_015_611, w_007_546, w_004_021);
  or2  I015_618(w_015_618, w_004_025, w_006_255);
  and2 I015_619(w_015_619, w_011_259, w_004_037);
  not1 I015_621(w_015_621, w_014_603);
  or2  I015_624(w_015_624, w_000_173, w_010_403);
  not1 I015_625(w_015_625, w_014_365);
  or2  I015_629(w_015_629, w_004_014, w_006_214);
  and2 I015_631(w_015_631, w_009_024, w_012_312);
  nand2 I015_635(w_015_635, w_003_140, w_002_443);
  or2  I015_636(w_015_636, w_006_030, w_008_007);
  and2 I015_643(w_015_643, w_003_040, w_006_216);
  nand2 I015_644(w_015_644, w_012_149, w_004_036);
  nand2 I015_648(w_015_648, w_012_185, w_011_009);
  or2  I015_652(w_015_652, w_005_048, w_000_177);
  or2  I015_654(w_015_654, w_008_220, w_000_115);
  not1 I015_655(w_015_655, w_011_477);
  nand2 I015_657(w_015_657, w_003_100, w_003_108);
  or2  I015_659(w_015_659, w_012_428, w_009_055);
  and2 I015_661(w_015_661, w_003_152, w_013_243);
  nand2 I015_669(w_015_669, w_013_202, w_005_281);
  and2 I015_676(w_015_676, w_007_303, w_013_207);
  nand2 I015_689(w_015_689, w_013_019, w_004_029);
  or2  I015_691(w_015_691, w_007_446, w_014_092);
  nand2 I015_692(w_015_692, w_002_247, w_011_511);
  and2 I015_693(w_015_693, w_010_082, w_000_751);
  not1 I015_695(w_015_695, w_011_016);
  or2  I015_696(w_015_696, w_009_042, w_009_013);
  or2  I015_699(w_015_699, w_000_446, w_013_197);
  or2  I015_703(w_015_703, w_010_255, w_010_612);
  nand2 I015_704(w_015_704, w_006_035, w_007_504);
  nand2 I015_706(w_015_706, w_000_869, w_002_450);
  nand2 I015_707(w_015_707, w_008_765, w_009_057);
  or2  I015_713(w_015_713, w_004_036, w_010_649);
  not1 I015_714(w_015_714, w_010_766);
  not1 I015_716(w_015_716, w_004_035);
  nand2 I015_718(w_015_718, w_002_235, w_009_016);
  nand2 I015_722(w_015_722, w_004_017, w_011_347);
  not1 I015_730(w_015_730, w_001_457);
  not1 I015_733(w_015_733, w_012_171);
  and2 I015_734(w_015_734, w_010_011, w_008_921);
  nand2 I015_737(w_015_737, w_000_804, w_002_124);
  and2 I015_738(w_015_738, w_009_055, w_002_232);
  and2 I015_742(w_015_742, w_004_033, w_001_038);
  or2  I015_743(w_015_743, w_013_075, w_012_130);
  and2 I015_744(w_015_744, w_006_273, w_003_219);
  nand2 I015_755(w_015_755, w_012_026, w_013_031);
  or2  I015_758(w_015_758, w_004_027, w_010_130);
  and2 I015_759(w_015_759, w_004_004, w_007_142);
  or2  I015_760(w_015_760, w_004_028, w_014_264);
  or2  I015_761(w_015_761, w_003_041, w_012_344);
  and2 I015_763(w_015_763, w_010_388, w_011_568);
  and2 I015_766(w_015_766, w_006_025, w_011_650);
  nand2 I015_773(w_015_773, w_014_293, w_009_035);
  and2 I015_774(w_015_774, w_006_036, w_014_061);
  and2 I015_776(w_015_776, w_013_158, w_003_124);
  and2 I015_778(w_015_778, w_006_286, w_005_544);
  and2 I015_779(w_015_779, w_011_317, w_008_835);
  not1 I015_780(w_015_780, w_010_078);
  or2  I015_782(w_015_782, w_008_276, w_003_067);
  not1 I015_793(w_015_793, w_011_082);
  not1 I016_001(w_016_001, w_009_042);
  nand2 I016_002(w_016_002, w_010_415, w_006_060);
  or2  I016_003(w_016_003, w_015_280, w_012_220);
  not1 I016_004(w_016_004, w_006_322);
  and2 I016_006(w_016_006, w_002_428, w_014_277);
  not1 I016_007(w_016_007, w_005_211);
  nand2 I016_010(w_016_010, w_004_028, w_003_150);
  and2 I016_012(w_016_012, w_011_394, w_012_114);
  not1 I016_013(w_016_013, w_014_542);
  not1 I016_016(w_016_016, w_001_171);
  nand2 I016_021(w_016_021, w_003_024, w_000_770);
  or2  I016_022(w_016_022, w_013_350, w_004_014);
  or2  I016_024(w_016_024, w_007_190, w_004_036);
  and2 I016_025(w_016_025, w_006_295, w_001_771);
  or2  I016_026(w_016_026, w_003_070, w_000_402);
  and2 I016_027(w_016_027, w_007_245, w_011_094);
  nand2 I016_028(w_016_028, w_004_018, w_006_017);
  nand2 I016_029(w_016_029, w_015_027, w_004_011);
  and2 I016_034(w_016_034, w_001_673, w_013_192);
  not1 I016_035(w_016_035, w_000_455);
  or2  I016_036(w_016_036, w_005_013, w_012_238);
  not1 I016_037(w_016_037, w_014_164);
  not1 I016_038(w_016_038, w_011_271);
  not1 I016_039(w_016_039, w_010_034);
  and2 I016_040(w_016_040, w_012_113, w_006_127);
  and2 I016_042(w_016_042, w_009_004, w_004_037);
  not1 I016_043(w_016_043, w_012_389);
  nand2 I016_047(w_016_047, w_015_315, w_002_325);
  not1 I016_048(w_016_048, w_002_149);
  nand2 I016_049(w_016_049, w_011_315, w_007_303);
  not1 I016_050(w_016_050, w_003_019);
  nand2 I016_052(w_016_052, w_005_467, w_010_699);
  nand2 I016_053(w_016_053, w_008_241, w_000_915);
  and2 I016_054(w_016_054, w_000_230, w_002_269);
  or2  I016_057(w_016_057, w_003_052, w_010_688);
  and2 I016_059(w_016_059, w_013_050, w_003_185);
  nand2 I016_060(w_016_060, w_004_006, w_004_009);
  or2  I016_062(w_016_062, w_004_026, w_011_675);
  not1 I016_063(w_016_063, w_000_462);
  nand2 I016_064(w_016_064, w_011_502, w_010_047);
  nand2 I016_065(w_016_065, w_013_235, w_003_092);
  and2 I016_067(w_016_067, w_004_028, w_015_155);
  nand2 I016_070(w_016_070, w_015_173, w_002_056);
  or2  I016_072(w_016_072, w_010_468, w_006_087);
  nand2 I016_074(w_016_074, w_010_097, w_005_109);
  and2 I016_075(w_016_075, w_008_588, w_013_431);
  nand2 I016_076(w_016_076, w_001_422, w_000_643);
  and2 I016_077(w_016_077, w_015_168, w_006_020);
  not1 I016_079(w_016_079, w_006_098);
  or2  I016_081(w_016_081, w_009_027, w_008_927);
  or2  I016_083(w_016_083, w_015_233, w_010_021);
  or2  I016_084(w_016_084, w_014_061, w_008_182);
  and2 I016_085(w_016_085, w_015_049, w_012_072);
  not1 I016_089(w_016_089, w_014_420);
  nand2 I016_090(w_016_090, w_008_793, w_000_030);
  or2  I016_093(w_016_093, w_009_012, w_015_369);
  and2 I016_096(w_016_096, w_013_052, w_007_302);
  nand2 I016_099(w_016_099, w_007_409, w_005_320);
  nand2 I016_100(w_016_100, w_004_003, w_007_218);
  and2 I016_101(w_016_101, w_015_479, w_007_251);
  and2 I016_102(w_016_102, w_007_236, w_000_068);
  nand2 I016_104(w_016_104, w_003_143, w_008_947);
  not1 I016_105(w_016_105, w_008_346);
  nand2 I016_106(w_016_106, w_013_178, w_006_297);
  not1 I016_108(w_016_108, w_009_052);
  nand2 I016_110(w_016_110, w_004_003, w_003_039);
  and2 I016_111(w_016_111, w_003_220, w_007_316);
  not1 I016_112(w_016_112, w_011_662);
  not1 I016_113(w_016_113, w_005_065);
  nand2 I016_114(w_016_114, w_000_767, w_004_037);
  and2 I016_116(w_016_116, w_012_108, w_000_401);
  not1 I016_122(w_016_122, w_000_669);
  nand2 I016_124(w_016_124, w_007_068, w_003_009);
  or2  I016_125(w_016_125, w_002_388, w_011_291);
  not1 I016_127(w_016_127, w_001_629);
  or2  I016_128(w_016_128, w_015_043, w_009_044);
  not1 I016_129(w_016_129, w_009_002);
  or2  I016_135(w_016_135, w_007_472, w_007_288);
  and2 I016_136(w_016_136, w_010_358, w_006_069);
  and2 I016_137(w_016_137, w_003_205, w_006_010);
  and2 I016_138(w_016_138, w_005_368, w_006_309);
  not1 I016_141(w_016_141, w_011_530);
  not1 I016_142(w_016_142, w_002_320);
  not1 I016_143(w_016_143, w_013_039);
  and2 I016_144(w_016_144, w_002_298, w_008_545);
  nand2 I016_146(w_016_146, w_004_007, w_014_124);
  nand2 I016_148(w_016_148, w_015_071, w_011_212);
  or2  I016_155(w_016_155, w_003_026, w_013_167);
  or2  I016_156(w_016_156, w_015_704, w_001_519);
  and2 I016_161(w_016_161, w_015_150, w_013_186);
  and2 I016_162(w_016_162, w_010_683, w_013_121);
  not1 I016_170(w_016_170, w_012_211);
  or2  I016_171(w_016_171, w_015_146, w_006_255);
  and2 I016_172(w_016_172, w_012_223, w_003_120);
  nand2 I016_173(w_016_173, w_007_238, w_004_008);
  nand2 I016_174(w_016_174, w_000_759, w_003_086);
  nand2 I016_175(w_016_175, w_001_026, w_011_161);
  or2  I016_178(w_016_178, w_013_386, w_013_392);
  not1 I016_179(w_016_179, w_000_040);
  or2  I016_181(w_016_181, w_015_209, w_000_344);
  and2 I016_182(w_016_182, w_011_186, w_000_756);
  or2  I016_184(w_016_184, w_002_195, w_007_296);
  nand2 I016_185(w_016_185, w_004_009, w_008_581);
  and2 I016_186(w_016_186, w_008_012, w_013_133);
  and2 I016_188(w_016_188, w_009_024, w_000_316);
  or2  I016_190(w_016_190, w_004_015, w_014_254);
  nand2 I016_191(w_016_191, w_005_103, w_010_642);
  nand2 I016_194(w_016_194, w_007_259, w_015_512);
  nand2 I016_195(w_016_195, w_000_181, w_005_425);
  nand2 I016_197(w_016_197, w_014_282, w_010_043);
  and2 I016_198(w_016_198, w_004_023, w_011_097);
  not1 I016_204(w_016_204, w_003_188);
  not1 I016_206(w_016_206, w_009_039);
  or2  I016_207(w_016_207, w_006_311, w_008_638);
  and2 I016_208(w_016_208, w_006_320, w_015_284);
  and2 I016_209(w_016_209, w_006_262, w_004_004);
  or2  I016_210(w_016_210, w_007_091, w_009_046);
  and2 I016_211(w_016_211, w_007_168, w_007_053);
  or2  I016_213(w_016_213, w_002_011, w_002_136);
  nand2 I016_214(w_016_214, w_011_456, w_005_026);
  or2  I016_215(w_016_215, w_006_012, w_013_057);
  and2 I016_217(w_016_217, w_015_766, w_000_886);
  nand2 I016_218(w_016_218, w_007_004, w_000_312);
  nand2 I016_219(w_016_219, w_001_723, w_008_772);
  or2  I016_220(w_016_220, w_011_327, w_006_143);
  or2  I016_221(w_016_221, w_011_175, w_010_280);
  not1 I016_224(w_016_224, w_006_113);
  not1 I016_225(w_016_225, w_006_091);
  or2  I016_226(w_016_226, w_007_254, w_001_139);
  and2 I016_228(w_016_228, w_013_219, w_014_237);
  or2  I016_232(w_016_232, w_015_214, w_002_292);
  not1 I016_235(w_016_235, w_015_716);
  nand2 I016_239(w_016_239, w_002_075, w_014_201);
  or2  I016_240(w_016_240, w_001_123, w_010_225);
  and2 I016_243(w_016_243, w_010_491, w_015_031);
  and2 I016_247(w_016_247, w_003_120, w_011_463);
  not1 I016_251(w_016_251, w_002_211);
  and2 I016_252(w_016_252, w_010_315, w_008_647);
  and2 I016_253(w_016_253, w_001_894, w_008_908);
  nand2 I016_255(w_016_255, w_015_001, w_011_008);
  nand2 I016_257(w_016_257, w_002_388, w_013_328);
  not1 I016_259(w_016_259, w_005_089);
  not1 I016_260(w_016_260, w_006_003);
  or2  I016_270(w_016_270, w_006_021, w_014_254);
  not1 I016_271(w_016_271, w_015_126);
  nand2 I016_272(w_016_272, w_007_283, w_008_515);
  and2 I016_273(w_016_273, w_012_236, w_015_438);
  not1 I016_274(w_016_274, w_015_482);
  not1 I016_275(w_016_275, w_000_728);
  and2 I016_276(w_016_276, w_015_499, w_007_156);
  and2 I016_278(w_016_278, w_008_941, w_012_262);
  and2 I016_281(w_016_281, w_007_384, w_010_007);
  and2 I016_282(w_016_282, w_006_258, w_003_085);
  not1 I016_285(w_016_285, w_005_445);
  not1 I016_289(w_016_289, w_010_822);
  not1 I016_290(w_016_290, w_001_002);
  or2  I016_295(w_016_295, w_012_025, w_012_109);
  nand2 I016_297(w_016_297, w_013_009, w_015_766);
  or2  I016_298(w_016_298, w_015_474, w_014_333);
  not1 I016_299(w_016_299, w_006_283);
  not1 I016_300(w_016_300, w_007_299);
  not1 I016_301(w_016_301, w_009_025);
  and2 I016_302(w_016_302, w_002_061, w_004_035);
  nand2 I016_303(w_016_303, w_010_491, w_010_198);
  and2 I016_305(w_016_305, w_008_722, w_004_007);
  and2 I016_306(w_016_306, w_009_002, w_007_068);
  not1 I016_307(w_016_307, w_014_287);
  or2  I016_313(w_016_313, w_000_753, w_015_051);
  and2 I016_315(w_016_315, w_001_046, w_006_096);
  not1 I016_316(w_016_316, w_006_075);
  and2 I016_317(w_016_317, w_003_072, w_015_738);
  not1 I016_318(w_016_318, w_006_046);
  nand2 I016_319(w_016_319, w_002_351, w_005_303);
  not1 I016_320(w_016_320, w_005_056);
  or2  I016_322(w_016_322, w_007_179, w_003_204);
  or2  I016_323(w_016_323, w_000_333, w_008_067);
  nand2 I016_326(w_016_326, w_002_469, w_013_470);
  not1 I016_327(w_016_327, w_010_084);
  not1 I016_328(w_016_328, w_008_407);
  and2 I016_329(w_016_329, w_000_586, w_003_078);
  and2 I016_330(w_016_330, w_003_085, w_012_494);
  nand2 I016_333(w_016_333, w_011_402, w_005_035);
  not1 I016_337(w_016_337, w_013_044);
  not1 I016_338(w_016_338, w_003_030);
  not1 I016_345(w_016_345, w_005_010);
  not1 I016_347(w_016_347, w_009_053);
  and2 I016_348(w_016_348, w_011_646, w_008_939);
  and2 I016_349(w_016_349, w_011_064, w_003_016);
  and2 I016_351(w_016_351, w_007_239, w_005_145);
  nand2 I016_353(w_016_353, w_010_092, w_001_036);
  nand2 I016_354(w_016_354, w_010_607, w_000_310);
  not1 I016_356(w_016_356, w_012_500);
  or2  I016_358(w_016_358, w_002_099, w_001_085);
  nand2 I016_359(w_016_359, w_014_251, w_011_209);
  not1 I016_362(w_016_362, w_012_276);
  and2 I016_363(w_016_363, w_009_059, w_001_022);
  nand2 I016_364(w_016_364, w_014_444, w_012_400);
  not1 I016_367(w_016_367, w_005_292);
  not1 I016_368(w_016_368, w_012_321);
  not1 I016_370(w_016_370, w_015_328);
  nand2 I016_371(w_016_371, w_008_889, w_003_171);
  and2 I016_372(w_016_372, w_006_277, w_013_419);
  or2  I016_374(w_016_374, w_006_045, w_003_104);
  not1 I016_376(w_016_376, w_015_064);
  not1 I016_378(w_016_378, w_014_053);
  nand2 I016_380(w_016_380, w_007_317, w_002_326);
  not1 I016_381(w_016_381, w_006_283);
  and2 I016_387(w_016_387, w_002_451, w_006_312);
  or2  I016_390(w_016_390, w_005_037, w_004_037);
  or2  I016_393(w_016_393, w_007_209, w_012_429);
  nand2 I016_394(w_016_394, w_001_882, w_003_178);
  nand2 I016_397(w_016_397, w_000_499, w_012_262);
  and2 I016_398(w_016_398, w_005_378, w_003_014);
  nand2 I016_400(w_016_400, w_000_740, w_007_042);
  not1 I016_404(w_016_404, w_012_221);
  nand2 I016_405(w_016_405, w_015_170, w_001_407);
  nand2 I016_406(w_016_406, w_003_215, w_007_229);
  nand2 I016_407(w_016_407, w_006_225, w_000_235);
  not1 I016_411(w_016_411, w_005_168);
  and2 I016_416(w_016_416, w_006_085, w_008_474);
  not1 I016_418(w_016_418, w_004_024);
  not1 I016_420(w_016_420, w_002_294);
  and2 I016_422(w_016_422, w_000_969, w_002_066);
  not1 I016_423(w_016_423, w_012_374);
  nand2 I016_424(w_016_424, w_008_893, w_005_105);
  nand2 I016_425(w_016_425, w_015_058, w_001_566);
  not1 I016_428(w_016_428, w_008_310);
  not1 I016_429(w_016_429, w_008_288);
  or2  I016_435(w_016_435, w_014_367, w_011_558);
  nand2 I016_436(w_016_436, w_008_024, w_009_049);
  not1 I016_437(w_016_437, w_007_252);
  and2 I016_438(w_016_438, w_010_049, w_013_107);
  nand2 I016_439(w_016_439, w_004_037, w_005_073);
  nand2 I016_440(w_016_440, w_015_036, w_011_261);
  or2  I016_442(w_016_442, w_000_661, w_012_280);
  or2  I016_445(w_016_445, w_006_317, w_000_882);
  and2 I016_448(w_016_448, w_000_209, w_005_097);
  nand2 I016_450(w_016_450, w_014_131, w_001_622);
  not1 I016_452(w_016_452, w_011_068);
  not1 I016_453(w_016_453, w_009_012);
  or2  I016_455(w_016_455, w_013_011, w_013_430);
  or2  I016_459(w_016_459, w_004_003, w_008_899);
  nand2 I016_461(w_016_461, w_008_609, w_004_019);
  nand2 I016_465(w_016_465, w_010_073, w_015_134);
  not1 I016_466(w_016_466, w_004_021);
  not1 I016_467(w_016_467, w_015_490);
  or2  I016_471(w_016_471, w_012_279, w_006_157);
  not1 I016_472(w_016_472, w_005_034);
  and2 I016_473(w_016_473, w_014_137, w_015_368);
  or2  I016_474(w_016_474, w_014_034, w_012_424);
  and2 I016_475(w_016_475, w_000_776, w_013_123);
  nand2 I016_476(w_016_476, w_003_192, w_012_182);
  and2 I016_477(w_016_477, w_006_262, w_013_481);
  nand2 I016_481(w_016_481, w_010_160, w_015_094);
  not1 I016_484(w_016_484, w_007_201);
  and2 I016_485(w_016_485, w_005_542, w_014_091);
  or2  I016_487(w_016_487, w_000_254, w_001_623);
  or2  I016_492(w_016_492, w_012_039, w_003_051);
  and2 I016_494(w_016_494, w_003_110, w_005_026);
  not1 I016_495(w_016_495, w_000_162);
  and2 I016_496(w_016_496, w_014_322, w_009_044);
  nand2 I016_500(w_016_500, w_015_458, w_002_181);
  not1 I016_501(w_016_501, w_005_394);
  and2 I017_000(w_017_000, w_007_404, w_001_608);
  not1 I017_001(w_017_001, w_016_171);
  and2 I017_002(w_017_002, w_006_117, w_003_174);
  not1 I017_003(w_017_003, w_002_421);
  or2  I017_004(w_017_004, w_001_088, w_008_599);
  not1 I017_005(w_017_005, w_008_598);
  and2 I017_006(w_017_006, w_000_131, w_012_429);
  or2  I017_007(w_017_007, w_014_269, w_014_123);
  nand2 I017_008(w_017_008, w_005_262, w_012_478);
  not1 I017_009(w_017_009, w_001_050);
  nand2 I017_010(w_017_010, w_005_023, w_005_253);
  nand2 I017_011(w_017_011, w_014_268, w_012_054);
  nand2 I017_012(w_017_012, w_011_004, w_000_340);
  and2 I017_013(w_017_013, w_012_321, w_002_139);
  nand2 I017_014(w_017_014, w_016_259, w_007_383);
  nand2 I017_015(w_017_015, w_002_421, w_003_084);
  and2 I017_016(w_017_016, w_006_062, w_004_005);
  and2 I017_017(w_017_017, w_016_349, w_008_275);
  or2  I017_018(w_017_018, w_000_535, w_012_375);
  nand2 I017_019(w_017_019, w_015_057, w_016_338);
  nand2 I017_020(w_017_020, w_011_476, w_015_418);
  nand2 I017_021(w_017_021, w_010_525, w_001_192);
  or2  I017_022(w_017_022, w_007_357, w_015_583);
  or2  I017_023(w_017_023, w_014_533, w_013_329);
  and2 I017_024(w_017_024, w_014_052, w_001_683);
  nand2 I017_025(w_017_025, w_008_432, w_002_120);
  nand2 I017_026(w_017_026, w_015_604, w_007_224);
  nand2 I017_027(w_017_027, w_010_467, w_006_211);
  or2  I018_000(w_018_000, w_002_430, w_001_060);
  not1 I018_002(w_018_002, w_013_105);
  and2 I018_003(w_018_003, w_009_042, w_013_375);
  or2  I018_006(w_018_006, w_003_047, w_008_154);
  nand2 I018_008(w_018_008, w_007_117, w_007_138);
  or2  I018_010(w_018_010, w_004_031, w_004_033);
  nand2 I018_013(w_018_013, w_008_727, w_010_468);
  or2  I018_014(w_018_014, w_001_006, w_017_006);
  and2 I018_015(w_018_015, w_006_091, w_008_327);
  nand2 I018_016(w_018_016, w_015_139, w_004_017);
  not1 I018_017(w_018_017, w_008_884);
  nand2 I018_019(w_018_019, w_009_045, w_002_355);
  or2  I018_020(w_018_020, w_012_321, w_001_811);
  or2  I018_021(w_018_021, w_000_097, w_003_008);
  and2 I018_023(w_018_023, w_009_060, w_014_608);
  nand2 I018_024(w_018_024, w_003_196, w_001_731);
  or2  I018_025(w_018_025, w_002_270, w_005_033);
  nand2 I018_026(w_018_026, w_003_073, w_009_009);
  nand2 I018_027(w_018_027, w_008_340, w_004_025);
  or2  I018_030(w_018_030, w_003_004, w_006_024);
  not1 I018_031(w_018_031, w_007_422);
  and2 I018_032(w_018_032, w_008_692, w_017_015);
  and2 I018_033(w_018_033, w_000_734, w_007_100);
  or2  I018_034(w_018_034, w_013_303, w_014_574);
  nand2 I018_035(w_018_035, w_010_335, w_015_031);
  or2  I018_036(w_018_036, w_003_075, w_002_186);
  nand2 I018_038(w_018_038, w_008_400, w_005_374);
  nand2 I018_039(w_018_039, w_003_032, w_017_012);
  nand2 I018_040(w_018_040, w_009_043, w_015_429);
  not1 I018_041(w_018_041, w_012_329);
  nand2 I018_043(w_018_043, w_001_531, w_003_190);
  or2  I018_046(w_018_046, w_012_245, w_016_353);
  and2 I018_047(w_018_047, w_005_078, w_007_162);
  and2 I018_048(w_018_048, w_002_051, w_010_519);
  nand2 I018_049(w_018_049, w_009_036, w_007_038);
  and2 I018_051(w_018_051, w_004_020, w_004_006);
  nand2 I018_052(w_018_052, w_003_109, w_010_226);
  and2 I018_053(w_018_053, w_002_167, w_013_136);
  not1 I018_054(w_018_054, w_005_170);
  not1 I018_056(w_018_056, w_010_181);
  not1 I018_057(w_018_057, w_000_970);
  not1 I018_058(w_018_058, w_009_019);
  not1 I018_059(w_018_059, w_004_008);
  or2  I018_060(w_018_060, w_013_114, w_009_020);
  and2 I018_062(w_018_062, w_009_032, w_002_249);
  and2 I018_064(w_018_064, w_009_018, w_016_370);
  or2  I018_066(w_018_066, w_009_038, w_008_557);
  nand2 I018_067(w_018_067, w_017_001, w_015_453);
  or2  I018_068(w_018_068, w_010_551, w_002_268);
  or2  I018_069(w_018_069, w_004_015, w_017_016);
  nand2 I018_070(w_018_070, w_013_285, w_009_021);
  or2  I018_072(w_018_072, w_009_023, w_016_298);
  and2 I018_073(w_018_073, w_006_043, w_015_462);
  not1 I018_074(w_018_074, w_010_078);
  and2 I018_075(w_018_075, w_000_818, w_014_472);
  and2 I018_076(w_018_076, w_000_839, w_009_039);
  not1 I018_077(w_018_077, w_004_018);
  or2  I018_079(w_018_079, w_014_253, w_007_010);
  not1 I018_081(w_018_081, w_000_848);
  not1 I018_082(w_018_082, w_001_667);
  and2 I018_084(w_018_084, w_004_028, w_006_009);
  and2 I018_086(w_018_086, w_000_898, w_009_065);
  or2  I018_088(w_018_088, w_002_353, w_007_097);
  and2 I018_089(w_018_089, w_010_665, w_007_299);
  and2 I018_090(w_018_090, w_009_008, w_015_275);
  and2 I018_091(w_018_091, w_014_409, w_006_038);
  or2  I018_092(w_018_092, w_008_078, w_017_000);
  or2  I018_093(w_018_093, w_009_047, w_009_022);
  nand2 I018_096(w_018_096, w_014_098, w_014_529);
  or2  I018_097(w_018_097, w_006_280, w_014_636);
  and2 I018_098(w_018_098, w_016_063, w_003_203);
  and2 I018_101(w_018_101, w_004_012, w_002_470);
  and2 I018_102(w_018_102, w_017_006, w_006_075);
  nand2 I018_103(w_018_103, w_016_475, w_011_201);
  and2 I018_104(w_018_104, w_016_272, w_009_040);
  and2 I018_106(w_018_106, w_006_044, w_002_371);
  and2 I018_107(w_018_107, w_009_056, w_004_025);
  not1 I018_108(w_018_108, w_004_027);
  not1 I018_109(w_018_109, w_003_013);
  and2 I018_110(w_018_110, w_014_026, w_004_009);
  and2 I018_111(w_018_111, w_015_706, w_010_121);
  nand2 I018_112(w_018_112, w_007_451, w_003_008);
  and2 I018_113(w_018_113, w_009_032, w_014_160);
  or2  I018_114(w_018_114, w_005_478, w_009_000);
  and2 I018_115(w_018_115, w_012_203, w_000_025);
  not1 I018_116(w_018_116, w_006_163);
  and2 I018_117(w_018_117, w_009_021, w_000_971);
  and2 I018_118(w_018_118, w_010_103, w_007_073);
  nand2 I018_119(w_018_119, w_010_060, w_009_020);
  not1 I018_120(w_018_120, w_005_379);
  nand2 I018_121(w_018_121, w_008_209, w_004_022);
  or2  I018_122(w_018_122, w_016_191, w_003_028);
  nand2 I018_123(w_018_123, w_008_015, w_015_621);
  not1 I018_124(w_018_124, w_016_101);
  not1 I018_125(w_018_125, w_008_706);
  or2  I018_126(w_018_126, w_006_280, w_015_053);
  nand2 I018_129(w_018_129, w_013_129, w_005_237);
  not1 I018_130(w_018_130, w_017_007);
  and2 I018_131(w_018_131, w_001_723, w_011_503);
  nand2 I018_132(w_018_132, w_012_069, w_013_054);
  not1 I018_133(w_018_133, w_001_020);
  nand2 I018_134(w_018_134, w_001_856, w_007_058);
  not1 I018_135(w_018_135, w_009_025);
  nand2 I018_136(w_018_136, w_010_011, w_009_036);
  or2  I018_139(w_018_139, w_001_597, w_014_240);
  and2 I018_141(w_018_141, w_003_013, w_000_314);
  not1 I018_143(w_018_143, w_003_044);
  and2 I018_144(w_018_144, w_014_357, w_015_079);
  or2  I018_145(w_018_145, w_003_125, w_005_380);
  not1 I018_146(w_018_146, w_004_008);
  not1 I018_150(w_018_150, w_006_098);
  not1 I018_151(w_018_151, w_001_121);
  or2  I018_153(w_018_153, w_008_050, w_010_633);
  nand2 I018_155(w_018_155, w_010_304, w_016_472);
  nand2 I018_156(w_018_156, w_006_317, w_011_159);
  and2 I018_157(w_018_157, w_015_127, w_009_030);
  and2 I018_158(w_018_158, w_000_073, w_011_669);
  or2  I018_159(w_018_159, w_016_398, w_013_258);
  and2 I018_163(w_018_163, w_016_155, w_012_192);
  not1 I018_164(w_018_164, w_003_050);
  nand2 I018_165(w_018_165, w_002_379, w_006_133);
  and2 I018_166(w_018_166, w_002_033, w_012_173);
  nand2 I018_167(w_018_167, w_003_130, w_009_016);
  not1 I018_168(w_018_168, w_012_218);
  or2  I018_170(w_018_170, w_001_055, w_006_235);
  or2  I018_171(w_018_171, w_016_144, w_006_286);
  or2  I018_172(w_018_172, w_008_332, w_009_036);
  and2 I018_174(w_018_174, w_005_302, w_005_403);
  nand2 I018_175(w_018_175, w_017_020, w_003_135);
  or2  I018_176(w_018_176, w_010_226, w_015_008);
  not1 I018_177(w_018_177, w_000_006);
  nand2 I018_180(w_018_180, w_000_886, w_001_539);
  nand2 I018_181(w_018_181, w_007_309, w_008_892);
  not1 I018_182(w_018_182, w_011_057);
  nand2 I018_183(w_018_183, w_002_137, w_016_038);
  or2  I018_184(w_018_184, w_015_045, w_014_626);
  nand2 I018_186(w_018_186, w_014_097, w_016_136);
  nand2 I018_188(w_018_188, w_011_318, w_003_021);
  or2  I018_190(w_018_190, w_017_016, w_010_751);
  not1 I018_191(w_018_191, w_002_445);
  nand2 I018_192(w_018_192, w_017_001, w_004_020);
  not1 I018_193(w_018_193, w_002_160);
  or2  I018_194(w_018_194, w_000_188, w_016_182);
  and2 I018_196(w_018_196, w_000_722, w_016_197);
  nand2 I018_197(w_018_197, w_013_026, w_006_065);
  or2  I018_198(w_018_198, w_006_027, w_002_062);
  or2  I019_002(w_019_002, w_016_327, w_012_098);
  and2 I019_004(w_019_004, w_016_206, w_017_000);
  nand2 I019_005(w_019_005, w_016_500, w_013_291);
  and2 I019_008(w_019_008, w_006_253, w_005_363);
  not1 I019_010(w_019_010, w_014_143);
  not1 I019_011(w_019_011, w_011_309);
  and2 I019_012(w_019_012, w_008_505, w_005_239);
  or2  I019_014(w_019_014, w_016_315, w_010_127);
  or2  I019_015(w_019_015, w_013_224, w_016_295);
  or2  I019_019(w_019_019, w_008_761, w_017_010);
  nand2 I019_020(w_019_020, w_003_157, w_004_030);
  and2 I019_021(w_019_021, w_015_742, w_017_007);
  nand2 I019_024(w_019_024, w_012_117, w_006_131);
  and2 I019_025(w_019_025, w_004_008, w_016_329);
  and2 I019_026(w_019_026, w_014_503, w_013_415);
  or2  I019_027(w_019_027, w_017_011, w_009_066);
  and2 I019_032(w_019_032, w_016_093, w_014_392);
  or2  I019_037(w_019_037, w_014_042, w_006_186);
  or2  I019_039(w_019_039, w_016_235, w_010_278);
  not1 I019_040(w_019_040, w_004_017);
  and2 I019_042(w_019_042, w_013_313, w_017_002);
  not1 I019_043(w_019_043, w_006_084);
  and2 I019_044(w_019_044, w_001_127, w_000_581);
  and2 I019_046(w_019_046, w_018_090, w_003_027);
  nand2 I019_048(w_019_048, w_017_019, w_003_050);
  and2 I019_049(w_019_049, w_001_768, w_001_516);
  or2  I019_050(w_019_050, w_014_245, w_015_165);
  nand2 I019_051(w_019_051, w_017_019, w_003_078);
  or2  I019_055(w_019_055, w_013_424, w_004_000);
  and2 I019_056(w_019_056, w_002_236, w_016_016);
  or2  I019_057(w_019_057, w_009_062, w_008_874);
  or2  I019_060(w_019_060, w_008_107, w_016_074);
  or2  I019_064(w_019_064, w_010_486, w_017_018);
  nand2 I019_065(w_019_065, w_000_153, w_003_012);
  or2  I019_067(w_019_067, w_014_063, w_003_075);
  not1 I019_068(w_019_068, w_014_017);
  and2 I019_069(w_019_069, w_003_162, w_008_794);
  and2 I019_070(w_019_070, w_010_406, w_017_010);
  not1 I019_072(w_019_072, w_016_362);
  not1 I019_073(w_019_073, w_001_188);
  nand2 I019_074(w_019_074, w_010_474, w_003_093);
  not1 I019_077(w_019_077, w_004_014);
  nand2 I019_078(w_019_078, w_005_453, w_018_130);
  not1 I019_082(w_019_082, w_016_144);
  nand2 I019_084(w_019_084, w_018_086, w_007_423);
  nand2 I019_085(w_019_085, w_009_023, w_010_514);
  nand2 I019_088(w_019_088, w_002_246, w_009_049);
  and2 I019_089(w_019_089, w_000_163, w_017_025);
  or2  I019_092(w_019_092, w_015_084, w_002_087);
  and2 I019_093(w_019_093, w_017_013, w_018_183);
  or2  I019_094(w_019_094, w_000_891, w_011_259);
  or2  I019_096(w_019_096, w_015_427, w_016_282);
  nand2 I019_097(w_019_097, w_011_011, w_013_303);
  nand2 I019_099(w_019_099, w_004_011, w_001_244);
  nand2 I019_100(w_019_100, w_000_506, w_018_136);
  nand2 I019_101(w_019_101, w_018_027, w_003_033);
  nand2 I019_102(w_019_102, w_001_119, w_014_534);
  not1 I019_103(w_019_103, w_008_318);
  or2  I019_111(w_019_111, w_011_673, w_016_329);
  not1 I019_116(w_019_116, w_014_150);
  nand2 I019_118(w_019_118, w_005_232, w_013_112);
  nand2 I019_121(w_019_121, w_001_820, w_017_002);
  not1 I019_124(w_019_124, w_016_072);
  or2  I019_125(w_019_125, w_003_158, w_003_057);
  nand2 I019_126(w_019_126, w_004_036, w_012_043);
  or2  I019_128(w_019_128, w_011_258, w_014_303);
  not1 I019_129(w_019_129, w_015_214);
  not1 I019_130(w_019_130, w_000_191);
  nand2 I019_133(w_019_133, w_009_032, w_008_900);
  or2  I019_135(w_019_135, w_009_064, w_009_039);
  or2  I019_138(w_019_138, w_017_000, w_008_232);
  or2  I019_144(w_019_144, w_009_050, w_007_417);
  nand2 I019_145(w_019_145, w_010_450, w_012_321);
  nand2 I019_146(w_019_146, w_015_780, w_005_317);
  not1 I019_147(w_019_147, w_011_583);
  and2 I019_148(w_019_148, w_011_560, w_018_131);
  nand2 I019_149(w_019_149, w_002_439, w_014_219);
  or2  I019_152(w_019_152, w_015_761, w_015_737);
  or2  I019_153(w_019_153, w_017_026, w_012_077);
  or2  I019_154(w_019_154, w_016_259, w_011_467);
  nand2 I019_155(w_019_155, w_000_266, w_014_337);
  or2  I019_157(w_019_157, w_009_022, w_005_173);
  and2 I019_160(w_019_160, w_005_134, w_004_008);
  not1 I019_163(w_019_163, w_005_059);
  not1 I019_165(w_019_165, w_001_011);
  nand2 I019_168(w_019_168, w_007_035, w_004_009);
  or2  I019_169(w_019_169, w_000_602, w_001_800);
  or2  I019_170(w_019_170, w_003_108, w_014_298);
  nand2 I019_171(w_019_171, w_008_717, w_013_405);
  and2 I019_173(w_019_173, w_011_131, w_017_004);
  not1 I019_174(w_019_174, w_000_362);
  or2  I019_179(w_019_179, w_011_250, w_017_015);
  and2 I019_182(w_019_182, w_005_089, w_018_054);
  nand2 I019_184(w_019_184, w_012_427, w_005_366);
  not1 I019_185(w_019_185, w_007_021);
  or2  I019_186(w_019_186, w_002_126, w_011_495);
  and2 I019_187(w_019_187, w_005_099, w_008_722);
  not1 I019_191(w_019_191, w_012_154);
  and2 I019_192(w_019_192, w_011_253, w_002_293);
  or2  I019_197(w_019_197, w_009_046, w_012_411);
  and2 I019_200(w_019_200, w_005_005, w_009_064);
  nand2 I019_205(w_019_205, w_014_006, w_008_442);
  not1 I019_207(w_019_207, w_002_441);
  nand2 I019_209(w_019_209, w_015_450, w_000_647);
  or2  I019_213(w_019_213, w_011_163, w_017_006);
  not1 I019_214(w_019_214, w_016_053);
  or2  I019_215(w_019_215, w_018_046, w_012_069);
  nand2 I019_219(w_019_219, w_000_236, w_013_278);
  nand2 I019_228(w_019_228, w_010_295, w_005_142);
  and2 I019_229(w_019_229, w_002_080, w_004_004);
  nand2 I019_230(w_019_230, w_015_755, w_018_013);
  and2 I019_233(w_019_233, w_011_631, w_015_081);
  not1 I019_234(w_019_234, w_004_009);
  or2  I019_235(w_019_235, w_007_142, w_017_025);
  nand2 I019_241(w_019_241, w_014_069, w_018_165);
  and2 I019_242(w_019_242, w_014_221, w_010_453);
  not1 I019_243(w_019_243, w_015_035);
  and2 I019_245(w_019_245, w_010_261, w_001_322);
  and2 I019_246(w_019_246, w_000_795, w_012_188);
  or2  I019_248(w_019_248, w_012_197, w_007_045);
  or2  I019_249(w_019_249, w_018_067, w_013_320);
  nand2 I019_255(w_019_255, w_002_243, w_015_015);
  or2  I019_258(w_019_258, w_001_247, w_017_021);
  nand2 I019_259(w_019_259, w_011_233, w_007_524);
  and2 I019_260(w_019_260, w_018_097, w_013_470);
  not1 I019_261(w_019_261, w_003_209);
  nand2 I019_265(w_019_265, w_005_088, w_004_007);
  and2 I019_269(w_019_269, w_000_777, w_011_158);
  and2 I019_274(w_019_274, w_008_609, w_015_519);
  and2 I019_275(w_019_275, w_010_542, w_010_409);
  not1 I019_277(w_019_277, w_003_145);
  or2  I019_279(w_019_279, w_016_319, w_017_012);
  nand2 I019_286(w_019_286, w_012_374, w_017_015);
  or2  I019_288(w_019_288, w_004_001, w_006_068);
  not1 I019_291(w_019_291, w_009_019);
  not1 I019_294(w_019_294, w_009_028);
  and2 I019_295(w_019_295, w_010_392, w_013_285);
  and2 I019_296(w_019_296, w_001_263, w_017_010);
  and2 I019_297(w_019_297, w_011_171, w_018_003);
  not1 I019_299(w_019_299, w_011_679);
  not1 I019_300(w_019_300, w_010_020);
  and2 I019_303(w_019_303, w_007_147, w_015_071);
  or2  I019_305(w_019_305, w_016_393, w_002_253);
  and2 I019_306(w_019_306, w_014_142, w_008_861);
  not1 I019_307(w_019_307, w_014_300);
  and2 I019_308(w_019_308, w_011_297, w_002_257);
  not1 I019_310(w_019_310, w_003_038);
  nand2 I019_314(w_019_314, w_002_289, w_016_029);
  and2 I019_317(w_019_317, w_011_309, w_005_417);
  or2  I019_318(w_019_318, w_018_034, w_007_134);
  or2  I019_319(w_019_319, w_012_040, w_006_025);
  and2 I019_320(w_019_320, w_013_177, w_007_186);
  and2 I019_321(w_019_321, w_002_131, w_015_763);
  and2 I019_322(w_019_322, w_013_188, w_001_082);
  nand2 I019_327(w_019_327, w_007_020, w_012_447);
  not1 I019_329(w_019_329, w_002_253);
  not1 I019_332(w_019_332, w_017_010);
  and2 I019_335(w_019_335, w_011_097, w_008_158);
  and2 I019_339(w_019_339, w_002_235, w_000_671);
  nand2 I019_340(w_019_340, w_000_427, w_009_032);
  and2 I019_342(w_019_342, w_008_374, w_003_083);
  and2 I019_344(w_019_344, w_010_146, w_016_089);
  and2 I019_345(w_019_345, w_016_278, w_014_574);
  nand2 I019_347(w_019_347, w_007_161, w_008_176);
  or2  I019_352(w_019_352, w_005_330, w_008_213);
  nand2 I019_353(w_019_353, w_017_023, w_004_033);
  not1 I019_357(w_019_357, w_009_036);
  nand2 I019_359(w_019_359, w_016_381, w_017_025);
  and2 I019_360(w_019_360, w_002_139, w_011_274);
  or2  I019_362(w_019_362, w_005_026, w_015_197);
  nand2 I019_363(w_019_363, w_005_240, w_018_066);
  nand2 I019_364(w_019_364, w_004_025, w_012_306);
  nand2 I019_371(w_019_371, w_018_125, w_017_014);
  not1 I019_374(w_019_374, w_006_064);
  not1 I019_377(w_019_377, w_017_011);
  or2  I019_378(w_019_378, w_017_010, w_012_337);
  not1 I019_384(w_019_384, w_000_508);
  and2 I019_386(w_019_386, w_006_147, w_012_018);
  not1 I019_389(w_019_389, w_000_022);
  or2  I019_396(w_019_396, w_012_184, w_018_197);
  or2  I019_402(w_019_402, w_011_068, w_009_022);
  and2 I019_403(w_019_403, w_008_046, w_005_210);
  not1 I019_404(w_019_404, w_015_755);
  not1 I019_406(w_019_406, w_006_109);
  and2 I019_407(w_019_407, w_003_031, w_017_014);
  and2 I019_413(w_019_413, w_001_892, w_013_148);
  not1 I019_416(w_019_416, w_004_016);
  nand2 I019_417(w_019_417, w_002_435, w_012_023);
  and2 I019_421(w_019_421, w_009_026, w_014_632);
  or2  I020_000(w_020_000, w_008_604, w_009_068);
  or2  I020_001(w_020_001, w_003_190, w_006_165);
  and2 I020_002(w_020_002, w_019_384, w_011_374);
  not1 I020_003(w_020_003, w_000_923);
  nand2 I020_004(w_020_004, w_004_034, w_002_480);
  and2 I020_005(w_020_005, w_012_190, w_014_598);
  nand2 I020_006(w_020_006, w_006_067, w_000_794);
  and2 I020_007(w_020_007, w_009_007, w_006_104);
  nand2 I020_008(w_020_008, w_012_050, w_004_025);
  or2  I020_009(w_020_009, w_007_010, w_019_307);
  or2  I020_010(w_020_010, w_002_323, w_019_152);
  or2  I020_011(w_020_011, w_019_389, w_015_733);
  nand2 I020_012(w_020_012, w_003_033, w_012_151);
  or2  I020_013(w_020_013, w_008_425, w_016_026);
  or2  I020_014(w_020_014, w_003_045, w_004_003);
  nand2 I020_015(w_020_015, w_017_027, w_017_016);
  not1 I020_016(w_020_016, w_010_590);
  not1 I020_017(w_020_017, w_001_042);
  nand2 I020_019(w_020_019, w_014_256, w_011_269);
  or2  I020_020(w_020_020, w_012_142, w_001_041);
  and2 I020_021(w_020_021, w_016_059, w_012_236);
  and2 I020_022(w_020_022, w_001_175, w_005_294);
  or2  I020_023(w_020_023, w_007_459, w_003_020);
  not1 I020_024(w_020_024, w_007_272);
  not1 I020_025(w_020_025, w_010_377);
  not1 I020_026(w_020_026, w_004_010);
  or2  I020_027(w_020_027, w_013_450, w_013_420);
  nand2 I020_028(w_020_028, w_004_036, w_008_677);
  and2 I020_029(w_020_029, w_016_204, w_013_171);
  nand2 I020_030(w_020_030, w_002_446, w_011_153);
  not1 I020_032(w_020_032, w_017_005);
  and2 I020_033(w_020_033, w_013_013, w_006_260);
  or2  I020_034(w_020_034, w_011_017, w_005_360);
  not1 I020_035(w_020_035, w_005_038);
  not1 I020_036(w_020_036, w_001_671);
  nand2 I020_037(w_020_037, w_004_014, w_017_000);
  or2  I020_038(w_020_038, w_011_340, w_001_087);
  nand2 I020_039(w_020_039, w_009_007, w_008_294);
  not1 I020_040(w_020_040, w_001_285);
  and2 I020_041(w_020_041, w_000_079, w_007_318);
  and2 I020_042(w_020_042, w_003_051, w_001_328);
  nand2 I020_043(w_020_043, w_014_359, w_011_430);
  or2  I020_044(w_020_044, w_008_130, w_015_631);
  nand2 I020_045(w_020_045, w_016_070, w_002_167);
  and2 I020_046(w_020_046, w_011_278, w_002_324);
  or2  I020_047(w_020_047, w_018_106, w_016_085);
  nand2 I020_048(w_020_048, w_012_248, w_004_010);
  and2 I020_049(w_020_049, w_011_347, w_019_274);
  or2  I020_050(w_020_050, w_005_075, w_019_340);
  or2  I020_052(w_020_052, w_017_001, w_001_228);
  and2 I020_053(w_020_053, w_003_000, w_013_033);
  or2  I020_054(w_020_054, w_009_049, w_016_253);
  or2  I020_057(w_020_057, w_014_260, w_019_096);
  and2 I020_058(w_020_058, w_008_253, w_005_169);
  or2  I020_060(w_020_060, w_019_168, w_008_347);
  not1 I020_061(w_020_061, w_019_207);
  and2 I020_062(w_020_062, w_010_570, w_014_013);
  and2 I020_063(w_020_063, w_008_861, w_001_742);
  or2  I020_064(w_020_064, w_013_191, w_013_241);
  nand2 I020_066(w_020_066, w_012_139, w_017_011);
  nand2 I020_067(w_020_067, w_017_022, w_001_308);
  or2  I020_068(w_020_068, w_010_730, w_007_196);
  and2 I020_069(w_020_069, w_008_484, w_017_025);
  nand2 I020_070(w_020_070, w_011_222, w_010_144);
  and2 I020_071(w_020_071, w_018_136, w_019_056);
  nand2 I020_072(w_020_072, w_018_176, w_010_827);
  nand2 I020_073(w_020_073, w_009_050, w_005_336);
  and2 I020_074(w_020_074, w_002_341, w_015_042);
  or2  I020_075(w_020_075, w_019_228, w_005_261);
  and2 I020_077(w_020_077, w_010_257, w_019_149);
  or2  I020_078(w_020_078, w_018_188, w_002_228);
  and2 I020_080(w_020_080, w_016_035, w_001_011);
  nand2 I020_081(w_020_081, w_002_104, w_001_748);
  not1 I020_082(w_020_082, w_013_475);
  not1 I020_083(w_020_083, w_019_303);
  not1 I020_084(w_020_084, w_009_008);
  or2  I020_085(w_020_085, w_010_717, w_011_029);
  nand2 I020_086(w_020_086, w_011_596, w_001_160);
  and2 I020_087(w_020_087, w_016_481, w_016_065);
  not1 I020_088(w_020_088, w_019_153);
  or2  I020_089(w_020_089, w_001_033, w_005_316);
  nand2 I020_090(w_020_090, w_001_229, w_014_324);
  nand2 I020_091(w_020_091, w_015_088, w_004_006);
  not1 I020_092(w_020_092, w_007_427);
  or2  I020_093(w_020_093, w_018_023, w_018_113);
  not1 I020_095(w_020_095, w_002_231);
  nand2 I020_096(w_020_096, w_015_659, w_000_687);
  and2 I020_098(w_020_098, w_017_015, w_016_174);
  or2  I020_099(w_020_099, w_016_099, w_018_110);
  or2  I020_100(w_020_100, w_017_025, w_012_403);
  and2 I020_102(w_020_102, w_011_314, w_004_036);
  or2  I020_103(w_020_103, w_011_066, w_009_028);
  and2 I020_104(w_020_104, w_001_081, w_011_129);
  and2 I020_105(w_020_105, w_004_015, w_001_743);
  and2 I020_106(w_020_106, w_018_036, w_002_373);
  nand2 I020_107(w_020_107, w_011_047, w_003_021);
  or2  I020_108(w_020_108, w_007_183, w_011_111);
  or2  I020_111(w_020_111, w_000_869, w_007_094);
  and2 I020_112(w_020_112, w_000_192, w_008_254);
  or2  I020_114(w_020_114, w_000_046, w_012_411);
  not1 I020_115(w_020_115, w_019_126);
  and2 I020_116(w_020_116, w_004_028, w_015_517);
  or2  I020_117(w_020_117, w_000_242, w_007_532);
  and2 I020_118(w_020_118, w_014_186, w_008_186);
  nand2 I020_119(w_020_119, w_009_026, w_006_332);
  not1 I020_120(w_020_120, w_009_062);
  nand2 I020_121(w_020_121, w_001_874, w_019_234);
  and2 I020_122(w_020_122, w_010_204, w_013_146);
  not1 I020_123(w_020_123, w_000_015);
  and2 I020_124(w_020_124, w_000_258, w_007_065);
  not1 I020_126(w_020_126, w_008_542);
  nand2 I020_127(w_020_127, w_000_689, w_000_370);
  not1 I020_128(w_020_128, w_016_475);
  nand2 I020_129(w_020_129, w_003_110, w_007_239);
  not1 I020_130(w_020_130, w_004_038);
  and2 I020_131(w_020_131, w_018_089, w_004_008);
  or2  I020_132(w_020_132, w_002_467, w_002_288);
  nand2 I020_133(w_020_133, w_006_142, w_007_308);
  not1 I020_134(w_020_134, w_019_153);
  not1 I020_135(w_020_135, w_010_162);
  nand2 I020_136(w_020_136, w_019_342, w_010_111);
  not1 I020_137(w_020_137, w_001_390);
  not1 I021_000(w_021_000, w_006_116);
  nand2 I021_001(w_021_001, w_014_515, w_006_131);
  nand2 I021_003(w_021_003, w_001_333, w_001_090);
  not1 I021_006(w_021_006, w_015_265);
  and2 I021_007(w_021_007, w_000_381, w_008_684);
  and2 I021_008(w_021_008, w_013_481, w_005_004);
  not1 I021_009(w_021_009, w_013_252);
  or2  I021_010(w_021_010, w_015_141, w_005_493);
  and2 I021_012(w_021_012, w_004_006, w_004_008);
  or2  I021_013(w_021_013, w_019_242, w_011_118);
  or2  I021_014(w_021_014, w_019_413, w_014_225);
  and2 I021_016(w_021_016, w_016_048, w_005_030);
  nand2 I021_018(w_021_018, w_013_164, w_014_637);
  and2 I021_019(w_021_019, w_001_687, w_013_477);
  not1 I021_020(w_021_020, w_001_871);
  not1 I021_024(w_021_024, w_006_060);
  not1 I021_025(w_021_025, w_019_065);
  and2 I021_026(w_021_026, w_015_470, w_020_084);
  not1 I021_027(w_021_027, w_009_060);
  and2 I021_028(w_021_028, w_016_285, w_015_559);
  not1 I021_029(w_021_029, w_005_516);
  or2  I021_030(w_021_030, w_001_234, w_003_085);
  not1 I021_033(w_021_033, w_014_389);
  and2 I021_035(w_021_035, w_018_079, w_008_896);
  and2 I021_036(w_021_036, w_017_018, w_000_142);
  nand2 I021_037(w_021_037, w_001_376, w_006_254);
  and2 I021_039(w_021_039, w_019_069, w_018_035);
  or2  I021_040(w_021_040, w_017_012, w_002_104);
  nand2 I021_041(w_021_041, w_015_363, w_015_214);
  and2 I021_042(w_021_042, w_012_287, w_009_034);
  and2 I021_044(w_021_044, w_011_203, w_000_557);
  nand2 I021_045(w_021_045, w_010_822, w_018_163);
  or2  I021_046(w_021_046, w_012_068, w_002_154);
  and2 I021_047(w_021_047, w_015_654, w_016_429);
  and2 I021_048(w_021_048, w_012_281, w_005_186);
  nand2 I021_049(w_021_049, w_000_692, w_002_309);
  or2  I021_050(w_021_050, w_018_049, w_000_563);
  or2  I021_051(w_021_051, w_010_143, w_018_166);
  nand2 I021_052(w_021_052, w_009_049, w_013_017);
  or2  I021_053(w_021_053, w_012_470, w_017_010);
  and2 I021_055(w_021_055, w_018_115, w_009_021);
  nand2 I021_058(w_021_058, w_003_011, w_014_270);
  not1 I021_059(w_021_059, w_001_035);
  or2  I021_060(w_021_060, w_011_109, w_004_026);
  and2 I021_061(w_021_061, w_009_031, w_014_264);
  and2 I021_063(w_021_063, w_002_196, w_003_144);
  not1 I021_064(w_021_064, w_017_020);
  not1 I021_065(w_021_065, w_020_003);
  and2 I021_066(w_021_066, w_010_757, w_020_069);
  or2  I021_070(w_021_070, w_002_049, w_017_002);
  nand2 I021_071(w_021_071, w_005_119, w_002_327);
  and2 I021_075(w_021_075, w_001_050, w_003_020);
  not1 I021_076(w_021_076, w_003_201);
  and2 I021_079(w_021_079, w_014_072, w_003_129);
  not1 I021_082(w_021_082, w_003_028);
  or2  I021_083(w_021_083, w_004_009, w_017_022);
  or2  I021_084(w_021_084, w_005_344, w_004_005);
  or2  I021_086(w_021_086, w_006_262, w_003_082);
  not1 I021_088(w_021_088, w_011_376);
  or2  I021_089(w_021_089, w_012_083, w_008_922);
  and2 I021_091(w_021_091, w_001_624, w_008_143);
  and2 I021_093(w_021_093, w_011_355, w_018_025);
  or2  I021_095(w_021_095, w_017_017, w_004_008);
  not1 I021_099(w_021_099, w_008_748);
  and2 I021_101(w_021_101, w_008_896, w_012_028);
  nand2 I021_105(w_021_105, w_000_544, w_017_002);
  or2  I021_106(w_021_106, w_017_016, w_008_210);
  not1 I021_107(w_021_107, w_020_080);
  nand2 I021_108(w_021_108, w_008_880, w_006_237);
  nand2 I021_111(w_021_111, w_002_374, w_005_121);
  nand2 I021_119(w_021_119, w_014_564, w_008_263);
  and2 I021_120(w_021_120, w_010_315, w_015_474);
  nand2 I021_122(w_021_122, w_009_028, w_010_772);
  and2 I021_123(w_021_123, w_004_028, w_005_045);
  or2  I021_126(w_021_126, w_003_222, w_019_163);
  not1 I021_127(w_021_127, w_009_004);
  nand2 I021_128(w_021_128, w_005_463, w_007_196);
  not1 I021_129(w_021_129, w_016_224);
  not1 I021_130(w_021_130, w_015_044);
  not1 I021_131(w_021_131, w_001_590);
  not1 I021_133(w_021_133, w_009_005);
  and2 I021_136(w_021_136, w_012_058, w_002_451);
  or2  I021_137(w_021_137, w_007_497, w_003_006);
  not1 I021_138(w_021_138, w_019_130);
  not1 I021_139(w_021_139, w_020_004);
  not1 I021_141(w_021_141, w_014_165);
  and2 I021_142(w_021_142, w_005_031, w_000_530);
  not1 I021_143(w_021_143, w_013_375);
  not1 I021_145(w_021_145, w_003_043);
  nand2 I021_149(w_021_149, w_008_490, w_003_018);
  and2 I021_151(w_021_151, w_010_565, w_016_001);
  and2 I021_152(w_021_152, w_009_038, w_013_189);
  nand2 I021_154(w_021_154, w_002_131, w_001_522);
  not1 I021_155(w_021_155, w_002_461);
  and2 I021_156(w_021_156, w_004_034, w_017_019);
  and2 I021_157(w_021_157, w_018_048, w_003_163);
  or2  I021_158(w_021_158, w_019_345, w_015_165);
  or2  I021_159(w_021_159, w_006_021, w_007_390);
  and2 I021_161(w_021_161, w_000_859, w_001_084);
  and2 I021_162(w_021_162, w_011_053, w_017_022);
  and2 I021_163(w_021_163, w_016_405, w_010_381);
  and2 I021_164(w_021_164, w_005_471, w_004_018);
  and2 I021_166(w_021_166, w_004_004, w_003_181);
  nand2 I021_169(w_021_169, w_020_063, w_009_006);
  not1 I021_170(w_021_170, w_019_317);
  not1 I021_171(w_021_171, w_001_210);
  and2 I021_172(w_021_172, w_020_061, w_015_090);
  or2  I021_178(w_021_178, w_016_106, w_018_024);
  or2  I021_179(w_021_179, w_018_006, w_012_158);
  or2  I021_181(w_021_181, w_015_151, w_008_595);
  and2 I021_183(w_021_183, w_020_063, w_015_349);
  nand2 I021_184(w_021_184, w_015_026, w_010_340);
  not1 I021_185(w_021_185, w_018_079);
  and2 I021_186(w_021_186, w_009_022, w_019_032);
  and2 I021_187(w_021_187, w_008_884, w_005_197);
  nand2 I021_190(w_021_190, w_020_082, w_001_446);
  nand2 I021_191(w_021_191, w_014_472, w_003_104);
  nand2 I021_192(w_021_192, w_019_186, w_007_200);
  and2 I021_194(w_021_194, w_004_014, w_015_304);
  or2  I021_195(w_021_195, w_015_029, w_013_045);
  or2  I021_198(w_021_198, w_005_247, w_007_068);
  not1 I021_199(w_021_199, w_003_023);
  not1 I021_201(w_021_201, w_004_008);
  nand2 I021_204(w_021_204, w_013_462, w_009_002);
  and2 I021_209(w_021_209, w_002_398, w_006_297);
  nand2 I021_210(w_021_210, w_006_263, w_006_222);
  and2 I021_211(w_021_211, w_013_449, w_010_768);
  not1 I021_215(w_021_215, w_015_730);
  and2 I021_218(w_021_218, w_008_806, w_006_055);
  or2  I021_219(w_021_219, w_019_146, w_007_394);
  not1 I021_220(w_021_220, w_006_087);
  or2  I021_221(w_021_221, w_018_158, w_011_142);
  or2  I021_222(w_021_222, w_004_014, w_011_372);
  not1 I021_224(w_021_224, w_011_659);
  nand2 I021_228(w_021_228, w_004_004, w_020_129);
  and2 I021_229(w_021_229, w_003_090, w_004_029);
  nand2 I021_230(w_021_230, w_007_033, w_019_069);
  or2  I021_234(w_021_234, w_008_379, w_004_005);
  not1 I021_236(w_021_236, w_015_193);
  nand2 I021_237(w_021_237, w_014_192, w_012_061);
  not1 I021_239(w_021_239, w_005_363);
  not1 I021_240(w_021_240, w_004_011);
  nand2 I021_243(w_021_243, w_020_010, w_002_085);
  and2 I021_244(w_021_244, w_014_270, w_013_213);
  or2  I021_245(w_021_245, w_013_006, w_008_636);
  not1 I021_247(w_021_247, w_018_046);
  nand2 I021_248(w_021_248, w_019_025, w_020_095);
  not1 I021_252(w_021_252, w_003_001);
  nand2 I021_256(w_021_256, w_013_396, w_013_449);
  not1 I021_257(w_021_257, w_010_597);
  not1 I021_259(w_021_259, w_005_029);
  or2  I021_261(w_021_261, w_003_100, w_001_115);
  nand2 I021_264(w_021_264, w_010_378, w_010_141);
  not1 I021_266(w_021_266, w_001_042);
  nand2 I021_270(w_021_270, w_005_165, w_004_037);
  nand2 I021_272(w_021_272, w_014_568, w_007_228);
  and2 I021_273(w_021_273, w_011_604, w_018_017);
  and2 I021_275(w_021_275, w_009_015, w_016_039);
  not1 I021_277(w_021_277, w_003_170);
  not1 I021_281(w_021_281, w_020_087);
  and2 I021_283(w_021_283, w_004_028, w_013_450);
  or2  I021_284(w_021_284, w_014_424, w_009_022);
  nand2 I021_289(w_021_289, w_009_055, w_007_099);
  nand2 I021_290(w_021_290, w_011_084, w_017_025);
  not1 I021_294(w_021_294, w_020_060);
  not1 I021_298(w_021_298, w_020_123);
  nand2 I021_303(w_021_303, w_006_256, w_014_230);
  nand2 I021_305(w_021_305, w_014_437, w_017_012);
  and2 I021_306(w_021_306, w_002_015, w_011_198);
  nand2 I021_307(w_021_307, w_002_074, w_004_000);
  or2  I021_310(w_021_310, w_015_597, w_014_070);
  not1 I021_313(w_021_313, w_005_486);
  or2  I021_314(w_021_314, w_005_560, w_010_714);
  not1 I021_317(w_021_317, w_008_010);
  or2  I021_319(w_021_319, w_005_574, w_006_013);
  not1 I021_320(w_021_320, w_003_178);
  and2 I021_322(w_021_322, w_018_014, w_018_123);
  nand2 I021_324(w_021_324, w_011_565, w_013_022);
  nand2 I021_326(w_021_326, w_016_037, w_005_024);
  not1 I021_328(w_021_328, w_006_074);
  and2 I021_329(w_021_329, w_001_813, w_010_749);
  not1 I021_330(w_021_330, w_007_304);
  or2  I021_335(w_021_335, w_002_305, w_012_504);
  nand2 I021_337(w_021_337, w_016_220, w_019_163);
  not1 I021_340(w_021_340, w_016_110);
  not1 I021_341(w_021_341, w_003_121);
  nand2 I021_342(w_021_342, w_000_452, w_013_005);
  nand2 I021_343(w_021_343, w_012_349, w_020_124);
  or2  I021_348(w_021_348, w_006_279, w_018_113);
  or2  I021_352(w_021_352, w_000_064, w_004_026);
  not1 I021_353(w_021_353, w_019_377);
  nand2 I021_360(w_021_360, w_015_559, w_004_016);
  or2  I022_002(w_022_002, w_017_014, w_012_378);
  or2  I022_003(w_022_003, w_013_273, w_013_194);
  and2 I022_006(w_022_006, w_009_037, w_008_194);
  nand2 I022_008(w_022_008, w_008_086, w_021_010);
  nand2 I022_010(w_022_010, w_004_028, w_000_765);
  or2  I022_020(w_022_020, w_018_016, w_003_106);
  or2  I022_021(w_022_021, w_002_497, w_006_058);
  or2  I022_025(w_022_025, w_015_078, w_008_737);
  nand2 I022_026(w_022_026, w_002_171, w_011_504);
  nand2 I022_031(w_022_031, w_003_150, w_018_051);
  or2  I022_032(w_022_032, w_007_551, w_012_098);
  nand2 I022_033(w_022_033, w_000_895, w_016_190);
  and2 I022_034(w_022_034, w_020_128, w_006_004);
  not1 I022_039(w_022_039, w_014_311);
  or2  I022_043(w_022_043, w_004_034, w_019_255);
  not1 I022_046(w_022_046, w_019_039);
  or2  I022_049(w_022_049, w_006_144, w_012_040);
  not1 I022_052(w_022_052, w_001_764);
  or2  I022_054(w_022_054, w_007_137, w_006_076);
  or2  I022_055(w_022_055, w_020_131, w_017_014);
  not1 I022_057(w_022_057, w_002_389);
  nand2 I022_061(w_022_061, w_010_014, w_004_017);
  or2  I022_065(w_022_065, w_017_021, w_017_015);
  and2 I022_066(w_022_066, w_005_116, w_000_730);
  and2 I022_067(w_022_067, w_021_061, w_020_005);
  not1 I022_068(w_022_068, w_008_346);
  or2  I022_072(w_022_072, w_005_333, w_018_089);
  or2  I022_073(w_022_073, w_018_023, w_014_307);
  or2  I022_076(w_022_076, w_000_482, w_006_115);
  and2 I022_081(w_022_081, w_015_603, w_011_645);
  nand2 I022_084(w_022_084, w_009_035, w_014_405);
  nand2 I022_087(w_022_087, w_021_224, w_003_142);
  nand2 I022_088(w_022_088, w_017_009, w_009_057);
  or2  I022_090(w_022_090, w_017_018, w_020_021);
  and2 I022_097(w_022_097, w_014_080, w_000_169);
  not1 I022_099(w_022_099, w_008_442);
  not1 I022_100(w_022_100, w_021_247);
  or2  I022_101(w_022_101, w_009_027, w_016_281);
  nand2 I022_103(w_022_103, w_008_034, w_016_076);
  and2 I022_105(w_022_105, w_008_213, w_013_405);
  and2 I022_109(w_022_109, w_001_514, w_015_604);
  not1 I022_110(w_022_110, w_001_093);
  and2 I022_113(w_022_113, w_018_090, w_021_047);
  and2 I022_117(w_022_117, w_005_031, w_017_008);
  not1 I022_118(w_022_118, w_010_074);
  nand2 I022_119(w_022_119, w_009_039, w_005_070);
  not1 I022_124(w_022_124, w_003_208);
  not1 I022_126(w_022_126, w_015_525);
  not1 I022_128(w_022_128, w_021_224);
  not1 I022_129(w_022_129, w_018_139);
  nand2 I022_139(w_022_139, w_017_022, w_005_353);
  not1 I022_143(w_022_143, w_014_582);
  not1 I022_144(w_022_144, w_008_545);
  or2  I022_146(w_022_146, w_002_181, w_014_420);
  and2 I022_149(w_022_149, w_017_008, w_015_625);
  not1 I022_151(w_022_151, w_009_040);
  not1 I022_152(w_022_152, w_010_484);
  or2  I022_155(w_022_155, w_012_096, w_014_417);
  nand2 I022_159(w_022_159, w_021_009, w_016_239);
  nand2 I022_160(w_022_160, w_005_094, w_013_357);
  nand2 I022_161(w_022_161, w_021_042, w_012_151);
  or2  I022_162(w_022_162, w_005_569, w_021_234);
  nand2 I022_163(w_022_163, w_007_347, w_007_234);
  not1 I022_165(w_022_165, w_017_023);
  not1 I022_168(w_022_168, w_016_347);
  not1 I022_169(w_022_169, w_006_227);
  and2 I022_174(w_022_174, w_001_481, w_014_191);
  or2  I022_175(w_022_175, w_021_122, w_000_535);
  nand2 I022_177(w_022_177, w_018_135, w_009_059);
  or2  I022_181(w_022_181, w_015_348, w_012_040);
  or2  I022_183(w_022_183, w_009_052, w_018_088);
  and2 I022_185(w_022_185, w_018_150, w_009_012);
  or2  I022_187(w_022_187, w_020_123, w_000_671);
  not1 I022_193(w_022_193, w_001_707);
  not1 I022_197(w_022_197, w_016_211);
  and2 I022_198(w_022_198, w_009_006, w_008_179);
  or2  I022_202(w_022_202, w_006_239, w_002_494);
  nand2 I022_205(w_022_205, w_018_116, w_009_032);
  not1 I022_206(w_022_206, w_019_032);
  or2  I022_209(w_022_209, w_003_112, w_015_394);
  not1 I022_210(w_022_210, w_003_094);
  or2  I022_213(w_022_213, w_015_655, w_003_113);
  and2 I022_222(w_022_222, w_000_305, w_000_057);
  nand2 I022_225(w_022_225, w_005_189, w_003_167);
  and2 I022_226(w_022_226, w_014_055, w_012_159);
  nand2 I022_229(w_022_229, w_010_193, w_009_038);
  and2 I022_234(w_022_234, w_012_422, w_003_188);
  nand2 I022_236(w_022_236, w_021_204, w_015_090);
  not1 I022_239(w_022_239, w_005_173);
  nand2 I022_242(w_022_242, w_006_058, w_005_069);
  or2  I022_243(w_022_243, w_020_116, w_018_036);
  not1 I022_244(w_022_244, w_007_254);
  and2 I022_246(w_022_246, w_013_187, w_013_045);
  not1 I022_256(w_022_256, w_010_099);
  not1 I022_258(w_022_258, w_005_167);
  nand2 I022_259(w_022_259, w_010_141, w_000_247);
  or2  I022_260(w_022_260, w_020_117, w_017_004);
  not1 I022_262(w_022_262, w_006_305);
  or2  I022_267(w_022_267, w_012_321, w_019_327);
  nand2 I022_268(w_022_268, w_018_164, w_021_126);
  or2  I022_269(w_022_269, w_017_005, w_009_016);
  nand2 I022_270(w_022_270, w_008_609, w_009_002);
  nand2 I022_271(w_022_271, w_000_169, w_015_779);
  nand2 I022_274(w_022_274, w_021_065, w_015_529);
  nand2 I022_275(w_022_275, w_009_011, w_015_114);
  and2 I022_276(w_022_276, w_012_113, w_004_003);
  and2 I022_277(w_022_277, w_019_364, w_016_358);
  or2  I022_278(w_022_278, w_012_409, w_021_178);
  and2 I022_280(w_022_280, w_009_039, w_001_321);
  nand2 I022_281(w_022_281, w_017_012, w_003_060);
  not1 I022_282(w_022_282, w_013_417);
  and2 I022_286(w_022_286, w_012_523, w_020_032);
  nand2 I022_290(w_022_290, w_014_594, w_019_148);
  nand2 I022_291(w_022_291, w_016_438, w_015_010);
  and2 I022_293(w_022_293, w_020_073, w_021_049);
  or2  I022_294(w_022_294, w_002_318, w_006_239);
  not1 I022_297(w_022_297, w_005_328);
  or2  I022_301(w_022_301, w_012_002, w_017_011);
  not1 I022_304(w_022_304, w_006_084);
  and2 I022_305(w_022_305, w_018_145, w_001_281);
  not1 I022_307(w_022_307, w_019_318);
  and2 I022_310(w_022_310, w_005_381, w_006_088);
  and2 I022_311(w_022_311, w_016_274, w_015_611);
  or2  I022_314(w_022_314, w_009_032, w_020_083);
  not1 I022_315(w_022_315, w_014_056);
  nand2 I022_316(w_022_316, w_012_453, w_000_022);
  nand2 I022_318(w_022_318, w_003_023, w_011_546);
  or2  I022_319(w_022_319, w_006_020, w_003_178);
  not1 I022_320(w_022_320, w_018_155);
  and2 I022_321(w_022_321, w_006_091, w_006_211);
  not1 I022_322(w_022_322, w_017_027);
  not1 I022_323(w_022_323, w_018_091);
  or2  I022_325(w_022_325, w_019_192, w_011_101);
  or2  I022_326(w_022_326, w_016_102, w_021_036);
  nand2 I022_328(w_022_328, w_010_407, w_007_463);
  and2 I022_335(w_022_335, w_016_027, w_009_004);
  and2 I022_336(w_022_336, w_013_254, w_002_060);
  nand2 I022_337(w_022_337, w_010_591, w_000_051);
  not1 I022_339(w_022_339, w_010_294);
  or2  I022_341(w_022_341, w_020_085, w_018_000);
  or2  I022_343(w_022_343, w_012_042, w_019_042);
  not1 I022_344(w_022_344, w_005_410);
  not1 I022_345(w_022_345, w_014_000);
  or2  I022_349(w_022_349, w_020_085, w_016_367);
  or2  I022_352(w_022_352, w_016_372, w_018_192);
  not1 I022_353(w_022_353, w_003_200);
  not1 I022_358(w_022_358, w_021_101);
  nand2 I022_360(w_022_360, w_018_114, w_012_216);
  nand2 I022_361(w_022_361, w_005_175, w_020_098);
  or2  I022_364(w_022_364, w_015_059, w_007_098);
  or2  I022_370(w_022_370, w_007_346, w_009_051);
  or2  I022_372(w_022_372, w_017_017, w_011_272);
  nand2 I022_375(w_022_375, w_006_196, w_018_074);
  not1 I022_376(w_022_376, w_015_061);
  not1 I022_383(w_022_383, w_018_024);
  and2 I022_385(w_022_385, w_008_675, w_020_061);
  or2  I022_388(w_022_388, w_007_484, w_002_396);
  or2  I022_391(w_022_391, w_006_257, w_008_282);
  or2  I022_392(w_022_392, w_004_013, w_010_323);
  nand2 I022_395(w_022_395, w_021_071, w_009_009);
  not1 I022_398(w_022_398, w_014_228);
  not1 I022_400(w_022_400, w_015_793);
  not1 I022_401(w_022_401, w_007_244);
  not1 I022_402(w_022_402, w_021_091);
  not1 I022_405(w_022_405, w_014_571);
  nand2 I022_406(w_022_406, w_002_081, w_007_000);
  nand2 I022_412(w_022_412, w_010_543, w_007_393);
  not1 I022_414(w_022_414, w_014_201);
  or2  I022_415(w_022_415, w_007_343, w_016_411);
  or2  I022_416(w_022_416, w_020_046, w_008_881);
  not1 I022_418(w_022_418, w_000_531);
  or2  I022_421(w_022_421, w_014_543, w_008_304);
  and2 I022_426(w_022_426, w_008_267, w_002_015);
  not1 I022_427(w_022_427, w_002_356);
  nand2 I022_428(w_022_428, w_016_247, w_007_342);
  nand2 I022_429(w_022_429, w_010_058, w_005_062);
  and2 I022_430(w_022_430, w_018_180, w_021_154);
  and2 I022_431(w_022_431, w_001_402, w_007_459);
  and2 I022_432(w_022_432, w_012_290, w_008_167);
  or2  I022_433(w_022_433, w_008_680, w_016_270);
  or2  I022_436(w_022_436, w_010_043, w_017_013);
  not1 I022_439(w_022_439, w_017_027);
  or2  I022_446(w_022_446, w_013_281, w_012_451);
  or2  I022_453(w_022_453, w_015_166, w_002_218);
  nand2 I022_455(w_022_455, w_001_391, w_016_099);
  not1 I022_457(w_022_457, w_003_223);
  and2 I022_464(w_022_464, w_009_061, w_007_346);
  nand2 I022_469(w_022_469, w_009_056, w_005_070);
  and2 I022_472(w_022_472, w_004_038, w_003_181);
  not1 I022_479(w_022_479, w_004_019);
  or2  I022_482(w_022_482, w_007_373, w_001_173);
  and2 I022_486(w_022_486, w_018_031, w_007_198);
  nand2 I022_489(w_022_489, w_008_827, w_016_065);
  nand2 I022_495(w_022_495, w_014_487, w_001_750);
  nand2 I022_498(w_022_498, w_005_169, w_005_181);
  nand2 I022_503(w_022_503, w_014_087, w_009_050);
  nand2 I022_506(w_022_506, w_013_463, w_015_157);
  nand2 I022_508(w_022_508, w_000_895, w_006_053);
  and2 I022_511(w_022_511, w_000_701, w_016_465);
  or2  I022_512(w_022_512, w_018_170, w_006_126);
  or2  I022_516(w_022_516, w_014_241, w_003_062);
  and2 I022_517(w_022_517, w_019_184, w_020_008);
  not1 I022_519(w_022_519, w_015_459);
  not1 I022_524(w_022_524, w_012_183);
  and2 I022_527(w_022_527, w_016_059, w_010_396);
  not1 I022_537(w_022_537, w_008_780);
  nand2 I022_540(w_022_540, w_011_044, w_021_061);
  or2  I022_543(w_022_543, w_010_005, w_018_129);
  or2  I023_002(w_023_002, w_002_325, w_006_154);
  or2  I023_012(w_023_012, w_002_490, w_003_152);
  and2 I023_013(w_023_013, w_006_168, w_003_173);
  not1 I023_015(w_023_015, w_006_324);
  nand2 I023_020(w_023_020, w_000_939, w_007_538);
  and2 I023_024(w_023_024, w_011_656, w_005_327);
  and2 I023_037(w_023_037, w_012_224, w_015_080);
  and2 I023_038(w_023_038, w_011_167, w_002_354);
  not1 I023_040(w_023_040, w_009_019);
  nand2 I023_041(w_023_041, w_013_373, w_008_216);
  nand2 I023_047(w_023_047, w_009_063, w_003_135);
  not1 I023_049(w_023_049, w_009_013);
  nand2 I023_051(w_023_051, w_022_002, w_017_021);
  nand2 I023_053(w_023_053, w_000_110, w_012_105);
  or2  I023_054(w_023_054, w_021_040, w_005_374);
  or2  I023_058(w_023_058, w_004_012, w_003_131);
  nand2 I023_059(w_023_059, w_016_281, w_008_383);
  and2 I023_064(w_023_064, w_018_060, w_019_092);
  nand2 I023_065(w_023_065, w_019_407, w_001_091);
  or2  I023_068(w_023_068, w_008_108, w_017_014);
  nand2 I023_071(w_023_071, w_000_190, w_007_105);
  not1 I023_073(w_023_073, w_017_015);
  not1 I023_078(w_023_078, w_005_369);
  or2  I023_079(w_023_079, w_018_008, w_005_311);
  and2 I023_086(w_023_086, w_005_042, w_007_164);
  or2  I023_088(w_023_088, w_022_129, w_007_121);
  nand2 I023_089(w_023_089, w_008_392, w_020_037);
  not1 I023_092(w_023_092, w_020_015);
  and2 I023_093(w_023_093, w_005_429, w_015_470);
  not1 I023_099(w_023_099, w_010_326);
  nand2 I023_100(w_023_100, w_021_329, w_012_218);
  nand2 I023_104(w_023_104, w_000_198, w_022_436);
  nand2 I023_106(w_023_106, w_017_012, w_015_150);
  not1 I023_108(w_023_108, w_009_014);
  not1 I023_109(w_023_109, w_019_103);
  not1 I023_110(w_023_110, w_006_085);
  not1 I023_111(w_023_111, w_019_089);
  nand2 I023_112(w_023_112, w_019_182, w_014_141);
  nand2 I023_118(w_023_118, w_001_599, w_018_167);
  nand2 I023_120(w_023_120, w_017_007, w_014_184);
  not1 I023_127(w_023_127, w_011_093);
  or2  I023_132(w_023_132, w_012_007, w_019_121);
  or2  I023_134(w_023_134, w_016_359, w_002_147);
  not1 I023_136(w_023_136, w_008_877);
  or2  I023_137(w_023_137, w_019_386, w_016_439);
  not1 I023_138(w_023_138, w_010_265);
  and2 I023_139(w_023_139, w_015_211, w_019_187);
  or2  I023_140(w_023_140, w_006_090, w_012_458);
  and2 I023_143(w_023_143, w_003_138, w_010_037);
  nand2 I023_148(w_023_148, w_012_519, w_007_194);
  not1 I023_153(w_023_153, w_006_073);
  or2  I023_154(w_023_154, w_013_107, w_001_689);
  and2 I023_157(w_023_157, w_018_174, w_001_820);
  not1 I023_158(w_023_158, w_006_318);
  not1 I023_161(w_023_161, w_000_378);
  or2  I023_166(w_023_166, w_005_184, w_014_403);
  and2 I023_170(w_023_170, w_016_440, w_012_128);
  and2 I023_172(w_023_172, w_002_002, w_003_164);
  and2 I023_174(w_023_174, w_005_023, w_008_044);
  or2  I023_175(w_023_175, w_015_155, w_004_036);
  or2  I023_177(w_023_177, w_002_041, w_016_476);
  and2 I023_178(w_023_178, w_009_003, w_011_078);
  or2  I023_181(w_023_181, w_013_330, w_019_295);
  or2  I023_184(w_023_184, w_012_432, w_008_604);
  or2  I023_186(w_023_186, w_002_129, w_004_020);
  nand2 I023_188(w_023_188, w_021_019, w_021_199);
  and2 I023_190(w_023_190, w_014_169, w_011_201);
  not1 I023_193(w_023_193, w_001_587);
  not1 I023_196(w_023_196, w_020_119);
  nand2 I023_197(w_023_197, w_007_136, w_007_101);
  or2  I023_200(w_023_200, w_022_152, w_011_351);
  nand2 I023_206(w_023_206, w_006_273, w_001_346);
  and2 I023_211(w_023_211, w_008_459, w_015_696);
  or2  I023_212(w_023_212, w_008_218, w_005_364);
  not1 I023_215(w_023_215, w_018_084);
  or2  I023_216(w_023_216, w_015_159, w_017_009);
  not1 I023_226(w_023_226, w_018_133);
  and2 I023_228(w_023_228, w_008_632, w_015_043);
  not1 I023_230(w_023_230, w_017_006);
  nand2 I023_231(w_023_231, w_005_356, w_018_126);
  nand2 I023_232(w_023_232, w_012_062, w_013_060);
  and2 I023_234(w_023_234, w_000_593, w_002_296);
  nand2 I023_239(w_023_239, w_003_037, w_022_103);
  not1 I023_240(w_023_240, w_022_181);
  not1 I023_241(w_023_241, w_022_126);
  not1 I023_242(w_023_242, w_019_055);
  nand2 I023_248(w_023_248, w_013_274, w_002_495);
  not1 I023_249(w_023_249, w_022_401);
  or2  I023_250(w_023_250, w_019_040, w_014_158);
  and2 I023_251(w_023_251, w_009_010, w_012_077);
  not1 I023_252(w_023_252, w_001_080);
  and2 I023_253(w_023_253, w_005_260, w_016_351);
  not1 I023_255(w_023_255, w_022_305);
  and2 I023_267(w_023_267, w_002_403, w_016_217);
  not1 I023_269(w_023_269, w_007_213);
  nand2 I023_271(w_023_271, w_010_004, w_022_155);
  not1 I023_274(w_023_274, w_017_009);
  nand2 I023_277(w_023_277, w_011_107, w_015_151);
  nand2 I023_278(w_023_278, w_003_048, w_011_106);
  or2  I023_291(w_023_291, w_006_314, w_016_471);
  nand2 I023_293(w_023_293, w_002_043, w_009_026);
  not1 I023_295(w_023_295, w_016_143);
  not1 I023_297(w_023_297, w_020_026);
  nand2 I023_302(w_023_302, w_012_179, w_018_047);
  or2  I023_305(w_023_305, w_000_053, w_021_161);
  and2 I023_306(w_023_306, w_015_554, w_001_387);
  not1 I023_307(w_023_307, w_014_140);
  not1 I023_309(w_023_309, w_020_034);
  and2 I023_311(w_023_311, w_019_078, w_020_086);
  and2 I023_316(w_023_316, w_020_019, w_001_046);
  and2 I023_321(w_023_321, w_007_158, w_012_149);
  nand2 I023_325(w_023_325, w_018_070, w_017_020);
  not1 I023_326(w_023_326, w_011_422);
  and2 I023_333(w_023_333, w_011_292, w_011_191);
  and2 I023_334(w_023_334, w_021_221, w_022_315);
  and2 I023_348(w_023_348, w_007_220, w_008_930);
  and2 I023_351(w_023_351, w_015_492, w_022_282);
  not1 I023_352(w_023_352, w_004_019);
  not1 I023_358(w_023_358, w_004_022);
  and2 I023_359(w_023_359, w_005_542, w_011_000);
  nand2 I023_369(w_023_369, w_012_456, w_013_119);
  not1 I023_383(w_023_383, w_002_127);
  and2 I023_387(w_023_387, w_007_192, w_020_035);
  nand2 I023_400(w_023_400, w_013_003, w_006_243);
  and2 I023_403(w_023_403, w_000_890, w_014_192);
  or2  I023_405(w_023_405, w_013_423, w_006_216);
  not1 I023_413(w_023_413, w_010_708);
  and2 I023_416(w_023_416, w_013_065, w_019_306);
  and2 I023_423(w_023_423, w_019_125, w_013_157);
  or2  I023_427(w_023_427, w_000_194, w_005_004);
  or2  I023_429(w_023_429, w_011_039, w_021_209);
  or2  I023_432(w_023_432, w_022_262, w_021_128);
  and2 I023_435(w_023_435, w_004_021, w_015_510);
  not1 I023_444(w_023_444, w_017_025);
  and2 I023_445(w_023_445, w_002_345, w_001_381);
  nand2 I023_448(w_023_448, w_005_059, w_019_026);
  not1 I023_451(w_023_451, w_022_020);
  nand2 I023_455(w_023_455, w_006_132, w_005_299);
  not1 I023_457(w_023_457, w_010_793);
  nand2 I023_459(w_023_459, w_006_322, w_017_024);
  nand2 I023_462(w_023_462, w_002_314, w_000_463);
  or2  I023_468(w_023_468, w_007_399, w_019_179);
  and2 I023_470(w_023_470, w_015_618, w_008_236);
  or2  I023_472(w_023_472, w_022_256, w_016_138);
  not1 I023_477(w_023_477, w_003_112);
  or2  I023_489(w_023_489, w_011_272, w_015_367);
  or2  I023_493(w_023_493, w_022_345, w_016_075);
  nand2 I023_499(w_023_499, w_022_400, w_012_154);
  or2  I023_500(w_023_500, w_005_284, w_005_384);
  or2  I023_502(w_023_502, w_016_173, w_007_188);
  or2  I023_503(w_023_503, w_015_333, w_019_286);
  and2 I023_507(w_023_507, w_006_163, w_012_415);
  and2 I023_513(w_023_513, w_007_322, w_006_015);
  or2  I023_518(w_023_518, w_001_486, w_009_062);
  not1 I023_520(w_023_520, w_013_431);
  or2  I023_522(w_023_522, w_011_227, w_020_070);
  nand2 I023_528(w_023_528, w_016_090, w_003_078);
  not1 I023_529(w_023_529, w_017_010);
  nand2 I023_530(w_023_530, w_007_413, w_012_185);
  or2  I023_531(w_023_531, w_016_495, w_013_406);
  nand2 I023_547(w_023_547, w_009_020, w_020_123);
  not1 I023_548(w_023_548, w_007_487);
  or2  I023_551(w_023_551, w_000_501, w_015_493);
  not1 I023_553(w_023_553, w_016_081);
  not1 I023_558(w_023_558, w_002_289);
  or2  I023_559(w_023_559, w_009_012, w_021_326);
  or2  I023_569(w_023_569, w_021_142, w_001_355);
  and2 I023_572(w_023_572, w_004_003, w_016_459);
  and2 I023_576(w_023_576, w_004_007, w_020_118);
  not1 I023_578(w_023_578, w_001_409);
  and2 I023_584(w_023_584, w_020_026, w_006_306);
  and2 I023_588(w_023_588, w_014_283, w_010_834);
  not1 I023_594(w_023_594, w_018_106);
  and2 I023_601(w_023_601, w_003_180, w_007_057);
  nand2 I023_603(w_023_603, w_019_173, w_017_005);
  nand2 I023_604(w_023_604, w_003_131, w_004_013);
  nand2 I023_611(w_023_611, w_009_000, w_019_082);
  not1 I023_614(w_023_614, w_012_022);
  and2 I023_621(w_023_621, w_004_016, w_009_024);
  or2  I023_622(w_023_622, w_006_319, w_000_687);
  nand2 I023_624(w_023_624, w_000_553, w_013_362);
  and2 I023_628(w_023_628, w_004_025, w_004_000);
  nand2 I023_633(w_023_633, w_006_112, w_014_064);
  and2 I023_656(w_023_656, w_006_009, w_011_125);
  nand2 I023_659(w_023_659, w_013_301, w_003_177);
  not1 I023_660(w_023_660, w_005_380);
  not1 I023_664(w_023_664, w_002_304);
  or2  I023_666(w_023_666, w_002_203, w_020_052);
  or2  I023_668(w_023_668, w_016_148, w_006_125);
  or2  I023_670(w_023_670, w_010_034, w_008_678);
  or2  I023_679(w_023_679, w_014_035, w_003_138);
  and2 I024_000(w_024_000, w_013_014, w_001_727);
  not1 I024_008(w_024_008, w_022_372);
  nand2 I024_012(w_024_012, w_014_310, w_012_107);
  or2  I024_014(w_024_014, w_000_395, w_020_060);
  or2  I024_019(w_024_019, w_001_027, w_010_103);
  not1 I024_020(w_024_020, w_003_150);
  nand2 I024_024(w_024_024, w_018_112, w_016_065);
  nand2 I024_029(w_024_029, w_015_238, w_008_172);
  not1 I024_034(w_024_034, w_008_406);
  and2 I024_037(w_024_037, w_009_032, w_003_088);
  not1 I024_040(w_024_040, w_017_019);
  or2  I024_041(w_024_041, w_022_021, w_023_228);
  not1 I024_042(w_024_042, w_021_058);
  and2 I024_050(w_024_050, w_018_043, w_020_068);
  nand2 I024_051(w_024_051, w_001_190, w_008_679);
  or2  I024_052(w_024_052, w_018_097, w_007_343);
  not1 I024_053(w_024_053, w_011_283);
  nand2 I024_056(w_024_056, w_014_609, w_019_012);
  not1 I024_057(w_024_057, w_015_171);
  nand2 I024_068(w_024_068, w_006_099, w_017_027);
  or2  I024_069(w_024_069, w_003_165, w_004_037);
  nand2 I024_070(w_024_070, w_008_862, w_012_317);
  and2 I024_072(w_024_072, w_007_262, w_013_170);
  and2 I024_076(w_024_076, w_001_127, w_007_089);
  not1 I024_079(w_024_079, w_011_231);
  nand2 I024_080(w_024_080, w_022_345, w_004_008);
  nand2 I024_082(w_024_082, w_004_015, w_012_301);
  nand2 I024_083(w_024_083, w_013_428, w_002_036);
  not1 I024_084(w_024_084, w_014_116);
  not1 I024_089(w_024_089, w_013_048);
  not1 I024_090(w_024_090, w_010_003);
  and2 I024_093(w_024_093, w_018_031, w_009_035);
  not1 I024_094(w_024_094, w_008_853);
  nand2 I024_096(w_024_096, w_011_150, w_012_426);
  not1 I024_103(w_024_103, w_021_156);
  or2  I024_104(w_024_104, w_004_019, w_019_362);
  nand2 I024_105(w_024_105, w_008_646, w_023_572);
  or2  I024_108(w_024_108, w_001_716, w_007_113);
  nand2 I024_112(w_024_112, w_022_301, w_002_082);
  nand2 I024_122(w_024_122, w_002_330, w_013_034);
  nand2 I024_128(w_024_128, w_001_024, w_013_310);
  and2 I024_129(w_024_129, w_015_644, w_023_068);
  or2  I024_130(w_024_130, w_009_033, w_002_112);
  not1 I024_131(w_024_131, w_018_092);
  nand2 I024_133(w_024_133, w_005_526, w_016_146);
  nand2 I024_136(w_024_136, w_019_165, w_001_492);
  nand2 I024_138(w_024_138, w_006_113, w_007_350);
  nand2 I024_141(w_024_141, w_007_041, w_011_569);
  and2 I024_142(w_024_142, w_007_315, w_020_067);
  or2  I024_145(w_024_145, w_019_342, w_003_207);
  not1 I024_146(w_024_146, w_019_048);
  nand2 I024_158(w_024_158, w_009_036, w_020_105);
  or2  I024_159(w_024_159, w_014_349, w_012_050);
  not1 I024_161(w_024_161, w_016_174);
  not1 I024_162(w_024_162, w_018_059);
  and2 I024_164(w_024_164, w_018_120, w_019_214);
  nand2 I024_166(w_024_166, w_015_062, w_014_268);
  nand2 I024_170(w_024_170, w_014_285, w_003_028);
  and2 I024_171(w_024_171, w_022_469, w_004_018);
  and2 I024_174(w_024_174, w_012_190, w_007_341);
  nand2 I024_176(w_024_176, w_017_017, w_009_039);
  nand2 I024_180(w_024_180, w_016_295, w_023_040);
  nand2 I024_182(w_024_182, w_016_285, w_006_110);
  or2  I024_183(w_024_183, w_015_773, w_002_244);
  not1 I024_189(w_024_189, w_002_219);
  and2 I024_191(w_024_191, w_020_014, w_011_260);
  not1 I024_192(w_024_192, w_021_106);
  or2  I024_194(w_024_194, w_016_240, w_014_635);
  nand2 I024_196(w_024_196, w_018_076, w_006_172);
  or2  I024_200(w_024_200, w_022_269, w_017_020);
  not1 I024_207(w_024_207, w_014_255);
  nand2 I024_209(w_024_209, w_017_021, w_021_289);
  and2 I024_217(w_024_217, w_015_442, w_006_243);
  or2  I024_218(w_024_218, w_010_157, w_007_460);
  and2 I024_220(w_024_220, w_004_030, w_022_151);
  and2 I024_225(w_024_225, w_015_635, w_022_343);
  or2  I024_228(w_024_228, w_009_009, w_010_158);
  not1 I024_229(w_024_229, w_010_632);
  not1 I024_231(w_024_231, w_013_032);
  or2  I024_236(w_024_236, w_020_008, w_013_013);
  and2 I024_238(w_024_238, w_006_260, w_010_023);
  not1 I024_244(w_024_244, w_008_434);
  not1 I024_247(w_024_247, w_022_540);
  and2 I024_249(w_024_249, w_022_202, w_001_369);
  or2  I024_251(w_024_251, w_019_148, w_009_052);
  not1 I024_255(w_024_255, w_020_092);
  nand2 I024_257(w_024_257, w_008_143, w_010_520);
  and2 I024_259(w_024_259, w_010_088, w_016_007);
  or2  I024_263(w_024_263, w_013_404, w_009_036);
  or2  I024_264(w_024_264, w_010_249, w_007_234);
  not1 I024_265(w_024_265, w_021_237);
  and2 I024_266(w_024_266, w_023_249, w_022_464);
  or2  I024_267(w_024_267, w_003_106, w_019_103);
  or2  I024_268(w_024_268, w_006_208, w_004_027);
  nand2 I024_270(w_024_270, w_021_240, w_009_038);
  and2 I024_276(w_024_276, w_010_234, w_000_515);
  nand2 I024_283(w_024_283, w_015_124, w_012_221);
  not1 I024_284(w_024_284, w_005_129);
  not1 I024_285(w_024_285, w_019_191);
  and2 I024_287(w_024_287, w_020_087, w_016_025);
  and2 I024_289(w_024_289, w_016_194, w_023_158);
  or2  I024_291(w_024_291, w_023_120, w_015_346);
  not1 I024_292(w_024_292, w_007_420);
  not1 I024_293(w_024_293, w_011_229);
  not1 I024_297(w_024_297, w_018_033);
  and2 I024_298(w_024_298, w_000_517, w_015_002);
  or2  I024_302(w_024_302, w_003_069, w_001_771);
  or2  I024_307(w_024_307, w_017_005, w_006_087);
  or2  I024_309(w_024_309, w_019_046, w_014_509);
  nand2 I024_316(w_024_316, w_011_003, w_017_012);
  or2  I024_319(w_024_319, w_012_463, w_003_049);
  nand2 I024_321(w_024_321, w_017_001, w_016_485);
  nand2 I024_322(w_024_322, w_008_279, w_006_279);
  and2 I024_323(w_024_323, w_000_676, w_013_208);
  and2 I024_326(w_024_326, w_017_025, w_004_027);
  and2 I024_331(w_024_331, w_011_180, w_005_026);
  nand2 I024_333(w_024_333, w_001_194, w_017_012);
  or2  I024_334(w_024_334, w_017_015, w_005_397);
  nand2 I024_335(w_024_335, w_017_001, w_011_112);
  nand2 I024_336(w_024_336, w_012_133, w_016_306);
  or2  I024_339(w_024_339, w_023_132, w_012_456);
  and2 I024_341(w_024_341, w_007_351, w_013_154);
  nand2 I024_342(w_024_342, w_006_232, w_010_463);
  nand2 I024_343(w_024_343, w_022_395, w_008_897);
  or2  I024_344(w_024_344, w_009_032, w_003_205);
  or2  I024_345(w_024_345, w_005_015, w_014_340);
  and2 I024_347(w_024_347, w_016_428, w_008_335);
  nand2 I024_351(w_024_351, w_012_226, w_016_035);
  not1 I024_353(w_024_353, w_003_111);
  and2 I024_357(w_024_357, w_001_022, w_016_135);
  and2 I024_361(w_024_361, w_014_263, w_010_212);
  and2 I024_364(w_024_364, w_001_167, w_019_171);
  not1 I024_366(w_024_366, w_015_143);
  and2 I024_367(w_024_367, w_006_162, w_018_107);
  not1 I024_377(w_024_377, w_003_045);
  not1 I024_380(w_024_380, w_011_232);
  not1 I024_381(w_024_381, w_010_536);
  not1 I024_382(w_024_382, w_009_001);
  and2 I024_388(w_024_388, w_005_033, w_019_010);
  or2  I024_391(w_024_391, w_005_403, w_014_221);
  and2 I024_393(w_024_393, w_014_538, w_001_093);
  and2 I024_394(w_024_394, w_020_027, w_005_314);
  not1 I024_397(w_024_397, w_000_491);
  and2 I024_398(w_024_398, w_006_046, w_003_044);
  nand2 I024_399(w_024_399, w_011_192, w_019_085);
  nand2 I024_400(w_024_400, w_020_022, w_019_069);
  nand2 I024_401(w_024_401, w_000_579, w_009_033);
  nand2 I024_402(w_024_402, w_013_260, w_021_209);
  and2 I024_404(w_024_404, w_006_264, w_004_015);
  or2  I024_407(w_024_407, w_015_096, w_016_065);
  nand2 I024_416(w_024_416, w_008_879, w_017_021);
  not1 I024_426(w_024_426, w_018_072);
  nand2 I024_429(w_024_429, w_004_003, w_015_154);
  not1 I024_435(w_024_435, w_018_097);
  not1 I024_437(w_024_437, w_010_116);
  nand2 I024_446(w_024_446, w_000_405, w_018_034);
  not1 I024_452(w_024_452, w_010_514);
  or2  I024_455(w_024_455, w_018_141, w_000_389);
  and2 I024_473(w_024_473, w_000_591, w_004_026);
  and2 I024_476(w_024_476, w_007_353, w_008_018);
  and2 I024_486(w_024_486, w_015_158, w_015_611);
  or2  I024_491(w_024_491, w_019_339, w_014_595);
  nand2 I024_495(w_024_495, w_000_788, w_006_031);
  and2 I024_496(w_024_496, w_005_408, w_001_510);
  nand2 I024_497(w_024_497, w_016_358, w_008_676);
  not1 I024_501(w_024_501, w_003_003);
  nand2 I024_507(w_024_507, w_010_297, w_004_023);
  and2 I024_511(w_024_511, w_019_032, w_021_000);
  or2  I024_515(w_024_515, w_006_067, w_014_311);
  and2 I024_522(w_024_522, w_010_606, w_011_121);
  and2 I024_523(w_024_523, w_002_007, w_005_163);
  or2  I024_529(w_024_529, w_003_048, w_017_026);
  not1 I024_537(w_024_537, w_015_049);
  not1 I024_539(w_024_539, w_022_160);
  nand2 I024_540(w_024_540, w_014_275, w_020_093);
  and2 I024_546(w_024_546, w_020_122, w_023_226);
  not1 I024_549(w_024_549, w_013_175);
  and2 I024_555(w_024_555, w_014_104, w_003_011);
  not1 I024_556(w_024_556, w_009_036);
  or2  I024_557(w_024_557, w_011_305, w_020_093);
  or2  I024_560(w_024_560, w_023_351, w_016_111);
  or2  I024_570(w_024_570, w_023_559, w_021_275);
  or2  I024_574(w_024_574, w_002_031, w_000_856);
  or2  I024_577(w_024_577, w_002_367, w_017_018);
  not1 I024_588(w_024_588, w_022_486);
  or2  I024_590(w_024_590, w_003_097, w_001_400);
  and2 I024_592(w_024_592, w_016_022, w_000_173);
  not1 I025_003(w_025_003, w_010_163);
  nand2 I025_005(w_025_005, w_024_264, w_012_091);
  or2  I025_008(w_025_008, w_008_002, w_012_367);
  and2 I025_009(w_025_009, w_001_850, w_008_036);
  not1 I025_011(w_025_011, w_000_964);
  not1 I025_012(w_025_012, w_013_407);
  nand2 I025_014(w_025_014, w_003_084, w_018_166);
  and2 I025_015(w_025_015, w_015_258, w_004_010);
  not1 I025_018(w_025_018, w_010_016);
  or2  I025_020(w_025_020, w_014_487, w_017_015);
  not1 I025_022(w_025_022, w_004_022);
  and2 I025_025(w_025_025, w_004_037, w_017_018);
  or2  I025_026(w_025_026, w_018_190, w_004_036);
  and2 I025_032(w_025_032, w_014_093, w_015_657);
  nand2 I025_033(w_025_033, w_022_239, w_015_175);
  nand2 I025_036(w_025_036, w_001_483, w_023_423);
  nand2 I025_039(w_025_039, w_005_517, w_005_250);
  not1 I025_041(w_025_041, w_007_297);
  or2  I025_042(w_025_042, w_016_108, w_011_109);
  and2 I025_047(w_025_047, w_001_124, w_009_061);
  or2  I025_050(w_025_050, w_004_032, w_002_125);
  not1 I025_056(w_025_056, w_018_059);
  nand2 I025_057(w_025_057, w_018_180, w_023_316);
  or2  I025_060(w_025_060, w_019_296, w_005_225);
  and2 I025_061(w_025_061, w_015_032, w_018_183);
  or2  I025_066(w_025_066, w_018_084, w_017_007);
  not1 I025_067(w_025_067, w_022_339);
  nand2 I025_068(w_025_068, w_014_520, w_019_169);
  and2 I025_071(w_025_071, w_012_070, w_004_012);
  or2  I025_075(w_025_075, w_014_267, w_007_350);
  and2 I025_077(w_025_077, w_005_346, w_020_010);
  not1 I025_079(w_025_079, w_003_156);
  or2  I025_083(w_025_083, w_023_584, w_021_322);
  or2  I025_087(w_025_087, w_010_628, w_016_042);
  nand2 I025_090(w_025_090, w_000_311, w_021_261);
  or2  I025_093(w_025_093, w_002_024, w_014_225);
  nand2 I025_094(w_025_094, w_007_347, w_016_416);
  or2  I025_100(w_025_100, w_022_391, w_002_430);
  and2 I025_103(w_025_103, w_010_680, w_014_269);
  or2  I025_105(w_025_105, w_022_055, w_010_461);
  and2 I025_107(w_025_107, w_005_147, w_020_048);
  not1 I025_108(w_025_108, w_002_201);
  and2 I025_115(w_025_115, w_016_003, w_011_186);
  and2 I025_125(w_025_125, w_017_002, w_011_280);
  or2  I025_126(w_025_126, w_007_250, w_001_213);
  or2  I025_131(w_025_131, w_023_297, w_011_534);
  nand2 I025_132(w_025_132, w_001_118, w_003_023);
  not1 I025_136(w_025_136, w_014_291);
  and2 I025_144(w_025_144, w_022_418, w_022_025);
  not1 I025_145(w_025_145, w_011_192);
  or2  I025_146(w_025_146, w_009_042, w_012_154);
  not1 I025_147(w_025_147, w_010_281);
  not1 I025_153(w_025_153, w_003_039);
  nand2 I025_154(w_025_154, w_007_177, w_008_866);
  or2  I025_155(w_025_155, w_014_399, w_023_321);
  nand2 I025_156(w_025_156, w_018_170, w_006_205);
  nand2 I025_157(w_025_157, w_001_679, w_001_328);
  or2  I025_158(w_025_158, w_014_198, w_017_012);
  nand2 I025_159(w_025_159, w_011_652, w_005_139);
  nand2 I025_160(w_025_160, w_003_145, w_023_489);
  nand2 I025_163(w_025_163, w_009_007, w_000_313);
  nand2 I025_169(w_025_169, w_005_143, w_008_389);
  not1 I025_171(w_025_171, w_022_003);
  not1 I025_177(w_025_177, w_000_309);
  not1 I025_180(w_025_180, w_023_216);
  nand2 I025_181(w_025_181, w_006_294, w_012_217);
  or2  I025_183(w_025_183, w_014_348, w_004_019);
  not1 I025_187(w_025_187, w_003_148);
  nand2 I025_188(w_025_188, w_015_122, w_013_451);
  or2  I025_189(w_025_189, w_013_096, w_020_127);
  not1 I025_195(w_025_195, w_005_336);
  and2 I025_199(w_025_199, w_003_163, w_024_336);
  and2 I025_202(w_025_202, w_004_002, w_005_388);
  or2  I025_203(w_025_203, w_011_044, w_006_031);
  not1 I025_206(w_025_206, w_023_369);
  and2 I025_208(w_025_208, w_018_193, w_008_004);
  not1 I025_215(w_025_215, w_013_280);
  nand2 I025_221(w_025_221, w_000_959, w_016_307);
  or2  I025_223(w_025_223, w_013_391, w_002_078);
  nand2 I025_225(w_025_225, w_018_196, w_015_350);
  or2  I025_226(w_025_226, w_000_831, w_001_474);
  or2  I025_228(w_025_228, w_015_691, w_015_053);
  or2  I025_232(w_025_232, w_020_089, w_024_220);
  and2 I025_233(w_025_233, w_002_196, w_001_020);
  and2 I025_238(w_025_238, w_008_474, w_021_136);
  nand2 I025_239(w_025_239, w_016_436, w_019_044);
  nand2 I025_246(w_025_246, w_013_448, w_009_001);
  and2 I025_247(w_025_247, w_023_212, w_008_182);
  or2  I025_250(w_025_250, w_018_102, w_009_011);
  and2 I025_251(w_025_251, w_003_075, w_000_271);
  or2  I025_262(w_025_262, w_006_059, w_013_272);
  or2  I025_269(w_025_269, w_013_264, w_015_499);
  not1 I025_272(w_025_272, w_015_156);
  and2 I025_274(w_025_274, w_014_130, w_022_226);
  nand2 I025_275(w_025_275, w_021_028, w_003_032);
  or2  I025_280(w_025_280, w_022_415, w_006_086);
  nand2 I025_281(w_025_281, w_005_217, w_007_551);
  not1 I025_282(w_025_282, w_012_162);
  not1 I025_286(w_025_286, w_019_173);
  not1 I025_290(w_025_290, w_010_404);
  nand2 I025_292(w_025_292, w_002_059, w_019_214);
  nand2 I025_294(w_025_294, w_020_131, w_004_029);
  nand2 I025_295(w_025_295, w_010_278, w_004_032);
  and2 I025_297(w_025_297, w_000_419, w_003_099);
  or2  I025_306(w_025_306, w_021_218, w_020_069);
  or2  I025_307(w_025_307, w_018_049, w_005_347);
  not1 I025_308(w_025_308, w_009_011);
  or2  I025_314(w_025_314, w_013_080, w_018_076);
  not1 I025_317(w_025_317, w_017_005);
  or2  I025_339(w_025_339, w_023_047, w_001_532);
  not1 I025_342(w_025_342, w_017_006);
  nand2 I025_346(w_025_346, w_010_061, w_019_057);
  nand2 I025_347(w_025_347, w_004_019, w_013_004);
  and2 I025_348(w_025_348, w_003_057, w_007_027);
  or2  I025_358(w_025_358, w_016_135, w_010_821);
  or2  I025_362(w_025_362, w_009_006, w_013_441);
  not1 I025_373(w_025_373, w_016_487);
  or2  I025_378(w_025_378, w_000_505, w_018_171);
  or2  I025_382(w_025_382, w_017_002, w_007_456);
  or2  I025_396(w_025_396, w_021_006, w_003_030);
  nand2 I025_405(w_025_405, w_016_065, w_006_210);
  not1 I025_406(w_025_406, w_022_405);
  and2 I025_412(w_025_412, w_003_073, w_010_523);
  nand2 I025_419(w_025_419, w_000_303, w_020_048);
  or2  I025_428(w_025_428, w_014_311, w_013_384);
  or2  I025_429(w_025_429, w_002_202, w_011_031);
  nand2 I025_437(w_025_437, w_006_276, w_024_333);
  or2  I025_454(w_025_454, w_002_154, w_018_066);
  nand2 I025_465(w_025_465, w_016_301, w_014_010);
  not1 I025_468(w_025_468, w_003_225);
  not1 I025_473(w_025_473, w_022_229);
  not1 I025_477(w_025_477, w_006_320);
  not1 I025_478(w_025_478, w_011_167);
  not1 I025_480(w_025_480, w_023_444);
  nand2 I025_488(w_025_488, w_006_242, w_013_486);
  and2 I025_497(w_025_497, w_017_022, w_013_064);
  not1 I025_498(w_025_498, w_021_187);
  not1 I025_506(w_025_506, w_008_450);
  and2 I025_510(w_025_510, w_005_478, w_010_218);
  or2  I025_514(w_025_514, w_017_003, w_014_443);
  not1 I025_516(w_025_516, w_021_245);
  and2 I025_519(w_025_519, w_019_260, w_017_022);
  nand2 I025_530(w_025_530, w_011_082, w_018_116);
  or2  I025_531(w_025_531, w_018_019, w_000_143);
  not1 I025_532(w_025_532, w_018_079);
  or2  I025_535(w_025_535, w_022_512, w_005_002);
  not1 I025_539(w_025_539, w_004_023);
  and2 I025_542(w_025_542, w_013_292, w_003_041);
  nand2 I025_552(w_025_552, w_002_173, w_017_006);
  and2 I025_553(w_025_553, w_019_010, w_000_649);
  not1 I025_554(w_025_554, w_006_214);
  not1 I025_555(w_025_555, w_022_316);
  or2  I025_556(w_025_556, w_015_080, w_019_160);
  nand2 I025_557(w_025_557, w_009_056, w_016_228);
  or2  I025_571(w_025_571, w_006_056, w_004_024);
  nand2 I025_572(w_025_572, w_000_723, w_020_060);
  nand2 I025_576(w_025_576, w_022_206, w_009_043);
  and2 I025_585(w_025_585, w_015_199, w_018_058);
  and2 I025_591(w_025_591, w_002_358, w_016_116);
  nand2 I025_595(w_025_595, w_014_043, w_019_040);
  not1 I025_606(w_025_606, w_006_166);
  nand2 I025_613(w_025_613, w_011_004, w_009_065);
  and2 I025_614(w_025_614, w_016_298, w_014_340);
  not1 I025_625(w_025_625, w_013_175);
  not1 I025_626(w_025_626, w_008_038);
  nand2 I025_630(w_025_630, w_021_036, w_017_001);
  or2  I025_635(w_025_635, w_022_168, w_018_086);
  or2  I025_640(w_025_640, w_011_464, w_019_032);
  and2 I025_648(w_025_648, w_011_395, w_011_224);
  or2  I025_654(w_025_654, w_008_319, w_000_487);
  and2 I025_656(w_025_656, w_016_012, w_010_819);
  nand2 I025_657(w_025_657, w_021_141, w_001_678);
  or2  I025_658(w_025_658, w_013_237, w_020_002);
  and2 I025_660(w_025_660, w_016_077, w_001_005);
  or2  I025_663(w_025_663, w_019_299, w_022_162);
  and2 I025_665(w_025_665, w_020_107, w_023_522);
  and2 I025_668(w_025_668, w_007_094, w_006_002);
  and2 I025_678(w_025_678, w_019_318, w_010_479);
  or2  I026_001(w_026_001, w_021_036, w_022_242);
  and2 I026_003(w_026_003, w_000_877, w_011_349);
  nand2 I026_007(w_026_007, w_001_082, w_023_099);
  not1 I026_008(w_026_008, w_011_176);
  nand2 I026_009(w_026_009, w_005_560, w_007_333);
  and2 I026_011(w_026_011, w_019_396, w_002_138);
  or2  I026_012(w_026_012, w_002_071, w_007_233);
  or2  I026_014(w_026_014, w_010_479, w_012_057);
  or2  I026_017(w_026_017, w_001_111, w_010_446);
  and2 I026_023(w_026_023, w_024_540, w_000_900);
  nand2 I026_024(w_026_024, w_010_698, w_001_752);
  or2  I026_025(w_026_025, w_024_342, w_002_344);
  or2  I026_026(w_026_026, w_023_049, w_017_017);
  or2  I026_028(w_026_028, w_014_247, w_012_308);
  or2  I026_029(w_026_029, w_018_139, w_008_582);
  and2 I026_030(w_026_030, w_010_834, w_006_179);
  or2  I026_031(w_026_031, w_009_057, w_024_400);
  not1 I026_032(w_026_032, w_002_242);
  not1 I026_034(w_026_034, w_007_109);
  nand2 I026_035(w_026_035, w_021_187, w_005_315);
  and2 I026_037(w_026_037, w_020_032, w_022_143);
  and2 I026_038(w_026_038, w_018_030, w_022_076);
  and2 I026_039(w_026_039, w_004_006, w_016_300);
  or2  I026_040(w_026_040, w_018_048, w_008_261);
  or2  I026_045(w_026_045, w_015_180, w_003_059);
  not1 I026_046(w_026_046, w_022_213);
  and2 I026_047(w_026_047, w_016_062, w_010_657);
  or2  I026_048(w_026_048, w_003_035, w_004_037);
  nand2 I026_049(w_026_049, w_018_174, w_023_601);
  or2  I026_051(w_026_051, w_024_170, w_008_145);
  nand2 I026_054(w_026_054, w_002_005, w_003_044);
  not1 I026_055(w_026_055, w_007_418);
  or2  I026_056(w_026_056, w_001_703, w_022_087);
  not1 I026_058(w_026_058, w_011_426);
  and2 I026_061(w_026_061, w_008_260, w_025_071);
  not1 I026_062(w_026_062, w_006_080);
  and2 I026_063(w_026_063, w_007_224, w_004_023);
  nand2 I026_064(w_026_064, w_012_373, w_012_345);
  and2 I026_065(w_026_065, w_024_079, w_019_219);
  not1 I026_068(w_026_068, w_024_130);
  not1 I026_073(w_026_073, w_005_175);
  nand2 I026_075(w_026_075, w_018_041, w_007_266);
  nand2 I026_078(w_026_078, w_015_779, w_002_369);
  nand2 I026_079(w_026_079, w_011_075, w_007_189);
  or2  I026_080(w_026_080, w_012_365, w_024_176);
  not1 I026_088(w_026_088, w_004_019);
  nand2 I026_089(w_026_089, w_002_132, w_024_259);
  not1 I026_091(w_026_091, w_006_239);
  nand2 I026_092(w_026_092, w_023_186, w_020_060);
  or2  I026_094(w_026_094, w_018_153, w_022_163);
  or2  I026_095(w_026_095, w_000_119, w_004_004);
  nand2 I026_096(w_026_096, w_002_429, w_001_846);
  not1 I026_097(w_026_097, w_012_460);
  and2 I026_098(w_026_098, w_020_033, w_012_375);
  nand2 I026_100(w_026_100, w_011_112, w_003_079);
  or2  I026_103(w_026_103, w_003_016, w_005_314);
  not1 I026_106(w_026_106, w_007_423);
  not1 I026_108(w_026_108, w_012_345);
  not1 I026_110(w_026_110, w_017_003);
  or2  I026_116(w_026_116, w_009_009, w_002_466);
  or2  I026_124(w_026_124, w_016_318, w_023_193);
  nand2 I026_125(w_026_125, w_004_034, w_015_319);
  and2 I026_131(w_026_131, w_025_262, w_012_269);
  and2 I026_139(w_026_139, w_005_311, w_005_039);
  and2 I026_142(w_026_142, w_020_134, w_020_063);
  not1 I026_149(w_026_149, w_003_166);
  and2 I026_155(w_026_155, w_004_015, w_014_256);
  or2  I026_156(w_026_156, w_009_061, w_015_535);
  not1 I026_158(w_026_158, w_021_277);
  nand2 I026_161(w_026_161, w_022_328, w_004_021);
  and2 I026_170(w_026_170, w_006_038, w_005_200);
  and2 I026_172(w_026_172, w_004_025, w_005_248);
  nand2 I026_174(w_026_174, w_013_446, w_021_089);
  nand2 I026_175(w_026_175, w_005_011, w_005_063);
  and2 I026_176(w_026_176, w_000_434, w_000_382);
  or2  I026_180(w_026_180, w_011_112, w_023_174);
  or2  I026_181(w_026_181, w_020_127, w_000_795);
  nand2 I026_183(w_026_183, w_017_019, w_025_556);
  nand2 I026_189(w_026_189, w_018_139, w_001_095);
  nand2 I026_194(w_026_194, w_010_074, w_013_363);
  and2 I026_195(w_026_195, w_016_105, w_013_291);
  not1 I026_200(w_026_200, w_009_030);
  nand2 I026_206(w_026_206, w_020_105, w_013_078);
  nand2 I026_209(w_026_209, w_016_420, w_004_020);
  and2 I026_210(w_026_210, w_013_458, w_001_251);
  nand2 I026_215(w_026_215, w_021_101, w_022_383);
  not1 I026_216(w_026_216, w_012_306);
  not1 I026_217(w_026_217, w_016_040);
  or2  I026_218(w_026_218, w_004_012, w_025_079);
  not1 I026_219(w_026_219, w_011_261);
  or2  I026_224(w_026_224, w_009_032, w_020_001);
  not1 I026_226(w_026_226, w_022_175);
  and2 I026_228(w_026_228, w_003_016, w_015_692);
  and2 I026_231(w_026_231, w_010_070, w_016_394);
  nand2 I026_232(w_026_232, w_022_197, w_020_137);
  not1 I026_235(w_026_235, w_016_024);
  not1 I026_236(w_026_236, w_002_325);
  and2 I026_239(w_026_239, w_006_270, w_016_142);
  or2  I026_243(w_026_243, w_018_089, w_005_016);
  and2 I026_246(w_026_246, w_013_277, w_023_111);
  nand2 I026_247(w_026_247, w_010_571, w_013_017);
  or2  I026_249(w_026_249, w_008_054, w_020_116);
  not1 I026_252(w_026_252, w_003_180);
  nand2 I026_253(w_026_253, w_017_025, w_008_926);
  or2  I026_257(w_026_257, w_019_261, w_011_094);
  nand2 I026_264(w_026_264, w_005_057, w_000_303);
  and2 I026_265(w_026_265, w_021_343, w_012_211);
  and2 I026_266(w_026_266, w_012_469, w_011_295);
  not1 I026_269(w_026_269, w_000_935);
  nand2 I026_272(w_026_272, w_002_294, w_015_058);
  and2 I026_273(w_026_273, w_003_075, w_001_771);
  and2 I026_274(w_026_274, w_023_271, w_021_211);
  or2  I026_275(w_026_275, w_002_490, w_003_174);
  and2 I026_277(w_026_277, w_011_434, w_009_019);
  and2 I026_279(w_026_279, w_013_488, w_020_122);
  nand2 I026_280(w_026_280, w_024_399, w_002_171);
  nand2 I026_282(w_026_282, w_005_436, w_025_221);
  or2  I026_283(w_026_283, w_005_168, w_020_004);
  and2 I026_294(w_026_294, w_011_022, w_024_322);
  and2 I026_295(w_026_295, w_015_776, w_001_127);
  and2 I026_296(w_026_296, w_004_003, w_022_315);
  or2  I026_297(w_026_297, w_006_057, w_010_376);
  or2  I026_298(w_026_298, w_013_279, w_006_018);
  or2  I026_301(w_026_301, w_012_058, w_021_230);
  not1 I026_303(w_026_303, w_015_462);
  or2  I026_305(w_026_305, w_003_124, w_016_374);
  and2 I026_307(w_026_307, w_023_211, w_009_007);
  or2  I026_308(w_026_308, w_004_037, w_014_061);
  and2 I026_309(w_026_309, w_007_200, w_010_746);
  not1 I026_310(w_026_310, w_014_442);
  not1 I026_311(w_026_311, w_004_006);
  not1 I026_317(w_026_317, w_025_317);
  nand2 I026_321(w_026_321, w_015_519, w_000_867);
  or2  I026_323(w_026_323, w_019_128, w_000_233);
  and2 I026_325(w_026_325, w_011_268, w_000_151);
  nand2 I026_326(w_026_326, w_000_352, w_025_075);
  not1 I026_328(w_026_328, w_006_036);
  or2  I026_331(w_026_331, w_004_026, w_003_013);
  and2 I026_332(w_026_332, w_005_069, w_015_278);
  or2  I026_333(w_026_333, w_014_032, w_013_375);
  and2 I026_338(w_026_338, w_023_321, w_020_093);
  nand2 I026_340(w_026_340, w_024_231, w_013_174);
  not1 I026_341(w_026_341, w_006_226);
  not1 I026_349(w_026_349, w_009_013);
  not1 I026_351(w_026_351, w_017_009);
  or2  I026_353(w_026_353, w_004_016, w_002_351);
  and2 I026_355(w_026_355, w_006_119, w_010_740);
  nand2 I026_356(w_026_356, w_019_174, w_000_183);
  and2 I026_358(w_026_358, w_018_040, w_018_033);
  nand2 I026_361(w_026_361, w_023_250, w_023_413);
  or2  I026_364(w_026_364, w_021_030, w_011_601);
  not1 I026_365(w_026_365, w_006_051);
  and2 I026_368(w_026_368, w_016_127, w_012_006);
  or2  I026_370(w_026_370, w_020_107, w_012_112);
  nand2 I026_374(w_026_374, w_012_048, w_008_555);
  or2  I026_375(w_026_375, w_020_009, w_024_207);
  nand2 I026_376(w_026_376, w_006_030, w_002_082);
  nand2 I026_377(w_026_377, w_015_692, w_010_171);
  and2 I026_379(w_026_379, w_015_330, w_021_324);
  nand2 I026_381(w_026_381, w_013_054, w_022_543);
  and2 I026_382(w_026_382, w_023_058, w_003_119);
  or2  I026_383(w_026_383, w_006_063, w_022_335);
  not1 I026_387(w_026_387, w_006_252);
  or2  I026_388(w_026_388, w_021_306, w_020_038);
  not1 I026_390(w_026_390, w_022_052);
  or2  I026_392(w_026_392, w_001_054, w_005_180);
  and2 I026_393(w_026_393, w_022_495, w_007_371);
  and2 I026_395(w_026_395, w_023_507, w_003_124);
  or2  I026_396(w_026_396, w_007_190, w_020_033);
  and2 I026_399(w_026_399, w_012_324, w_022_175);
  and2 I026_400(w_026_400, w_019_046, w_012_206);
  and2 I026_401(w_026_401, w_023_024, w_023_184);
  not1 I026_407(w_026_407, w_024_069);
  not1 I026_408(w_026_408, w_023_158);
  or2  I026_410(w_026_410, w_021_219, w_024_161);
  or2  I026_419(w_026_419, w_025_281, w_013_271);
  nand2 I026_421(w_026_421, w_011_423, w_025_429);
  not1 I026_424(w_026_424, w_000_734);
  and2 I026_430(w_026_430, w_014_210, w_025_136);
  or2  I026_431(w_026_431, w_017_026, w_013_104);
  and2 I026_435(w_026_435, w_008_665, w_005_104);
  and2 I026_436(w_026_436, w_009_007, w_000_475);
  or2  I026_438(w_026_438, w_018_020, w_025_066);
  not1 I027_006(w_027_006, w_016_322);
  nand2 I027_007(w_027_007, w_001_769, w_006_211);
  nand2 I027_011(w_027_011, w_019_144, w_010_200);
  nand2 I027_014(w_027_014, w_021_264, w_005_143);
  or2  I027_016(w_027_016, w_002_271, w_016_303);
  or2  I027_027(w_027_027, w_021_145, w_000_274);
  and2 I027_035(w_027_035, w_018_132, w_018_168);
  or2  I027_040(w_027_040, w_008_503, w_015_108);
  or2  I027_041(w_027_041, w_022_109, w_016_243);
  not1 I027_042(w_027_042, w_002_077);
  not1 I027_050(w_027_050, w_003_056);
  nand2 I027_054(w_027_054, w_005_100, w_018_064);
  and2 I027_055(w_027_055, w_004_003, w_018_159);
  nand2 I027_063(w_027_063, w_020_116, w_001_192);
  nand2 I027_067(w_027_067, w_026_277, w_018_025);
  or2  I027_069(w_027_069, w_010_741, w_020_107);
  or2  I027_075(w_027_075, w_019_133, w_008_692);
  not1 I027_077(w_027_077, w_019_297);
  or2  I027_080(w_027_080, w_008_610, w_016_418);
  or2  I027_083(w_027_083, w_021_079, w_021_158);
  and2 I027_085(w_027_085, w_000_158, w_012_357);
  and2 I027_087(w_027_087, w_023_502, w_020_133);
  and2 I027_091(w_027_091, w_020_070, w_026_170);
  nand2 I027_095(w_027_095, w_015_373, w_014_060);
  not1 I027_101(w_027_101, w_004_005);
  or2  I027_108(w_027_108, w_005_148, w_016_184);
  nand2 I027_111(w_027_111, w_011_520, w_000_405);
  and2 I027_114(w_027_114, w_020_133, w_000_301);
  not1 I027_115(w_027_115, w_021_088);
  and2 I027_118(w_027_118, w_001_170, w_007_007);
  nand2 I027_124(w_027_124, w_002_492, w_022_431);
  and2 I027_127(w_027_127, w_001_046, w_025_083);
  and2 I027_128(w_027_128, w_012_436, w_019_295);
  nand2 I027_130(w_027_130, w_003_145, w_019_245);
  not1 I027_134(w_027_134, w_017_004);
  or2  I027_141(w_027_141, w_006_124, w_005_011);
  nand2 I027_143(w_027_143, w_024_108, w_022_021);
  and2 I027_144(w_027_144, w_015_140, w_019_403);
  not1 I027_145(w_027_145, w_016_116);
  nand2 I027_154(w_027_154, w_021_184, w_016_435);
  and2 I027_162(w_027_162, w_023_518, w_005_380);
  not1 I027_164(w_027_164, w_023_251);
  nand2 I027_165(w_027_165, w_013_159, w_000_468);
  or2  I027_168(w_027_168, w_000_891, w_026_235);
  not1 I027_171(w_027_171, w_004_022);
  or2  I027_172(w_027_172, w_018_177, w_017_009);
  not1 I027_173(w_027_173, w_020_095);
  nand2 I027_177(w_027_177, w_020_036, w_016_257);
  and2 I027_189(w_027_189, w_014_329, w_017_012);
  and2 I027_195(w_027_195, w_009_028, w_006_144);
  and2 I027_198(w_027_198, w_018_066, w_010_111);
  and2 I027_207(w_027_207, w_013_013, w_012_012);
  and2 I027_208(w_027_208, w_024_367, w_004_025);
  nand2 I027_222(w_027_222, w_008_163, w_001_198);
  not1 I027_225(w_027_225, w_020_067);
  not1 I027_227(w_027_227, w_025_226);
  not1 I027_234(w_027_234, w_007_414);
  and2 I027_236(w_027_236, w_021_070, w_021_247);
  or2  I027_250(w_027_250, w_010_615, w_019_342);
  or2  I027_257(w_027_257, w_017_000, w_019_135);
  or2  I027_259(w_027_259, w_005_136, w_022_099);
  not1 I027_267(w_027_267, w_023_500);
  or2  I027_272(w_027_272, w_020_120, w_013_203);
  not1 I027_280(w_027_280, w_022_293);
  or2  I027_285(w_027_285, w_019_327, w_022_427);
  not1 I027_294(w_027_294, w_007_248);
  and2 I027_299(w_027_299, w_000_452, w_008_135);
  not1 I027_300(w_027_300, w_021_239);
  nand2 I027_307(w_027_307, w_010_392, w_013_487);
  nand2 I027_311(w_027_311, w_006_020, w_005_172);
  and2 I027_320(w_027_320, w_010_152, w_022_341);
  and2 I027_324(w_027_324, w_005_284, w_008_487);
  not1 I027_336(w_027_336, w_026_156);
  or2  I027_339(w_027_339, w_001_853, w_000_749);
  nand2 I027_343(w_027_343, w_002_000, w_009_045);
  and2 I027_344(w_027_344, w_004_009, w_006_028);
  nand2 I027_348(w_027_348, w_000_753, w_011_308);
  and2 I027_353(w_027_353, w_008_297, w_006_201);
  not1 I027_373(w_027_373, w_018_072);
  nand2 I027_383(w_027_383, w_006_300, w_018_122);
  not1 I027_400(w_027_400, w_003_168);
  or2  I027_401(w_027_401, w_015_322, w_004_031);
  or2  I027_412(w_027_412, w_009_000, w_024_336);
  or2  I027_413(w_027_413, w_019_012, w_020_084);
  nand2 I027_414(w_027_414, w_003_161, w_003_037);
  nand2 I027_419(w_027_419, w_015_758, w_012_045);
  nand2 I027_426(w_027_426, w_021_186, w_020_086);
  or2  I027_429(w_027_429, w_019_073, w_014_243);
  nand2 I027_431(w_027_431, w_001_020, w_000_636);
  or2  I027_433(w_027_433, w_020_046, w_026_195);
  not1 I027_434(w_027_434, w_005_462);
  and2 I027_437(w_027_437, w_001_829, w_007_054);
  and2 I027_440(w_027_440, w_026_008, w_024_050);
  or2  I027_445(w_027_445, w_018_188, w_012_314);
  not1 I027_459(w_027_459, w_019_342);
  and2 I027_460(w_027_460, w_026_333, w_002_422);
  nand2 I027_466(w_027_466, w_003_108, w_018_062);
  nand2 I027_470(w_027_470, w_012_383, w_019_130);
  and2 I027_478(w_027_478, w_023_184, w_017_017);
  nand2 I027_486(w_027_486, w_023_078, w_017_022);
  and2 I027_497(w_027_497, w_020_090, w_010_562);
  and2 I027_522(w_027_522, w_024_577, w_001_000);
  not1 I027_525(w_027_525, w_025_180);
  or2  I027_526(w_027_526, w_013_329, w_021_229);
  and2 I027_535(w_027_535, w_009_006, w_026_189);
  nand2 I027_537(w_027_537, w_014_573, w_003_147);
  or2  I027_543(w_027_543, w_008_527, w_003_062);
  nand2 I027_546(w_027_546, w_003_218, w_010_082);
  and2 I027_548(w_027_548, w_006_282, w_019_205);
  not1 I027_564(w_027_564, w_012_266);
  not1 I027_565(w_027_565, w_007_173);
  nand2 I027_568(w_027_568, w_006_169, w_003_174);
  not1 I027_573(w_027_573, w_016_013);
  or2  I027_576(w_027_576, w_022_270, w_003_106);
  and2 I027_584(w_027_584, w_014_602, w_006_056);
  and2 I027_600(w_027_600, w_008_237, w_007_276);
  and2 I027_602(w_027_602, w_012_284, w_003_202);
  not1 I027_606(w_027_606, w_005_155);
  not1 I027_614(w_027_614, w_006_326);
  and2 I027_619(w_027_619, w_022_361, w_013_307);
  nand2 I027_622(w_027_622, w_012_439, w_009_037);
  or2  I027_624(w_027_624, w_020_077, w_017_013);
  and2 I027_625(w_027_625, w_005_053, w_001_860);
  or2  I027_628(w_027_628, w_011_136, w_010_747);
  nand2 I027_629(w_027_629, w_008_474, w_011_221);
  and2 I027_635(w_027_635, w_001_146, w_007_513);
  or2  I027_647(w_027_647, w_026_161, w_019_246);
  and2 I027_656(w_027_656, w_022_068, w_023_079);
  nand2 I027_658(w_027_658, w_006_303, w_004_035);
  nand2 I027_659(w_027_659, w_025_208, w_005_214);
  or2  I027_663(w_027_663, w_025_157, w_007_436);
  not1 I027_668(w_027_668, w_016_333);
  or2  I027_671(w_027_671, w_020_108, w_020_041);
  or2  I027_672(w_027_672, w_017_023, w_018_060);
  nand2 I027_676(w_027_676, w_015_349, w_001_041);
  not1 I027_678(w_027_678, w_008_037);
  not1 I027_681(w_027_681, w_007_485);
  not1 I027_683(w_027_683, w_025_189);
  nand2 I027_690(w_027_690, w_020_048, w_018_155);
  or2  I027_696(w_027_696, w_016_037, w_003_159);
  or2  I027_699(w_027_699, w_001_771, w_020_006);
  or2  I027_707(w_027_707, w_013_143, w_017_001);
  not1 I027_712(w_027_712, w_018_077);
  nand2 I027_717(w_027_717, w_012_069, w_006_125);
  not1 I027_725(w_027_725, w_024_076);
  nand2 I027_736(w_027_736, w_023_138, w_025_626);
  and2 I027_742(w_027_742, w_016_368, w_021_228);
  not1 I027_757(w_027_757, w_014_331);
  or2  I027_762(w_027_762, w_011_126, w_017_001);
  not1 I027_768(w_027_768, w_022_061);
  or2  I027_776(w_027_776, w_021_266, w_003_138);
  not1 I027_779(w_027_779, w_017_024);
  and2 I027_791(w_027_791, w_007_311, w_020_098);
  and2 I027_794(w_027_794, w_011_033, w_023_086);
  and2 I027_796(w_027_796, w_024_497, w_009_027);
  or2  I027_797(w_027_797, w_012_289, w_020_038);
  and2 I027_811(w_027_811, w_002_021, w_003_095);
  and2 I027_813(w_027_813, w_004_023, w_008_830);
  and2 I027_816(w_027_816, w_005_472, w_007_169);
  nand2 I027_819(w_027_819, w_025_635, w_015_776);
  or2  I027_826(w_027_826, w_020_091, w_022_118);
  nand2 I028_004(w_028_004, w_011_213, w_010_344);
  not1 I028_012(w_028_012, w_001_311);
  nand2 I028_013(w_028_013, w_021_215, w_016_081);
  or2  I028_015(w_028_015, w_003_067, w_019_145);
  nand2 I028_017(w_028_017, w_011_056, w_012_287);
  not1 I028_020(w_028_020, w_027_696);
  nand2 I028_024(w_028_024, w_009_009, w_022_349);
  and2 I028_025(w_028_025, w_009_019, w_018_040);
  not1 I028_027(w_028_027, w_011_164);
  or2  I028_028(w_028_028, w_027_207, w_021_095);
  or2  I028_029(w_028_029, w_024_209, w_006_306);
  not1 I028_030(w_028_030, w_024_164);
  and2 I028_033(w_028_033, w_019_049, w_018_082);
  not1 I028_036(w_028_036, w_019_307);
  or2  I028_042(w_028_042, w_014_420, w_016_330);
  or2  I028_043(w_028_043, w_000_977, w_025_663);
  not1 I028_049(w_028_049, w_015_595);
  or2  I028_052(w_028_052, w_020_014, w_002_257);
  and2 I028_062(w_028_062, w_011_125, w_017_022);
  nand2 I028_065(w_028_065, w_027_294, w_006_214);
  not1 I028_066(w_028_066, w_006_240);
  or2  I028_067(w_028_067, w_004_005, w_001_399);
  and2 I028_070(w_028_070, w_009_044, w_020_037);
  not1 I028_073(w_028_073, w_019_099);
  or2  I028_076(w_028_076, w_025_342, w_020_123);
  or2  I028_078(w_028_078, w_003_056, w_010_012);
  or2  I028_079(w_028_079, w_026_421, w_018_144);
  not1 I028_081(w_028_081, w_002_123);
  and2 I028_087(w_028_087, w_027_725, w_005_547);
  nand2 I028_088(w_028_088, w_017_013, w_013_372);
  and2 I028_092(w_028_092, w_027_811, w_020_058);
  not1 I028_102(w_028_102, w_010_184);
  or2  I028_107(w_028_107, w_001_286, w_019_037);
  and2 I028_108(w_028_108, w_026_092, w_006_100);
  or2  I028_109(w_028_109, w_015_605, w_008_496);
  and2 I028_112(w_028_112, w_011_478, w_001_779);
  not1 I028_119(w_028_119, w_026_224);
  not1 I028_125(w_028_125, w_019_235);
  or2  I028_128(w_028_128, w_015_482, w_006_177);
  and2 I028_131(w_028_131, w_005_190, w_026_216);
  or2  I028_132(w_028_132, w_001_451, w_011_648);
  and2 I028_135(w_028_135, w_017_007, w_027_035);
  not1 I028_143(w_028_143, w_005_497);
  not1 I028_144(w_028_144, w_006_096);
  or2  I028_146(w_028_146, w_027_622, w_011_622);
  not1 I028_156(w_028_156, w_009_023);
  nand2 I028_161(w_028_161, w_013_300, w_011_407);
  and2 I028_162(w_028_162, w_017_022, w_024_053);
  nand2 I028_167(w_028_167, w_001_529, w_018_046);
  and2 I028_171(w_028_171, w_004_031, w_020_136);
  not1 I028_180(w_028_180, w_003_110);
  not1 I028_186(w_028_186, w_010_139);
  not1 I028_201(w_028_201, w_018_129);
  and2 I028_202(w_028_202, w_016_096, w_005_404);
  nand2 I028_206(w_028_206, w_011_650, w_021_317);
  nand2 I028_210(w_028_210, w_002_388, w_021_192);
  nand2 I028_211(w_028_211, w_017_011, w_024_189);
  and2 I028_216(w_028_216, w_000_726, w_004_021);
  nand2 I028_218(w_028_218, w_024_159, w_003_150);
  and2 I028_219(w_028_219, w_012_268, w_011_087);
  or2  I028_220(w_028_220, w_015_282, w_022_430);
  nand2 I028_222(w_028_222, w_005_413, w_018_000);
  nand2 I028_234(w_028_234, w_022_274, w_016_209);
  nand2 I028_235(w_028_235, w_016_299, w_020_064);
  or2  I028_237(w_028_237, w_010_833, w_002_364);
  or2  I028_241(w_028_241, w_003_180, w_017_003);
  and2 I028_246(w_028_246, w_002_182, w_019_269);
  or2  I028_258(w_028_258, w_013_311, w_025_272);
  not1 I028_276(w_028_276, w_011_172);
  not1 I028_277(w_028_277, w_023_232);
  or2  I028_281(w_028_281, w_020_069, w_010_061);
  nand2 I028_289(w_028_289, w_003_147, w_005_221);
  not1 I028_294(w_028_294, w_017_022);
  nand2 I028_296(w_028_296, w_026_045, w_017_019);
  not1 I028_302(w_028_302, w_000_290);
  and2 I028_311(w_028_311, w_011_278, w_008_918);
  nand2 I028_313(w_028_313, w_027_127, w_006_313);
  not1 I028_318(w_028_318, w_018_144);
  or2  I028_323(w_028_323, w_018_130, w_014_111);
  not1 I028_326(w_028_326, w_007_282);
  and2 I028_328(w_028_328, w_010_065, w_024_361);
  not1 I028_345(w_028_345, w_007_155);
  or2  I028_349(w_028_349, w_006_278, w_000_848);
  not1 I028_358(w_028_358, w_000_856);
  not1 I028_359(w_028_359, w_019_352);
  or2  I028_360(w_028_360, w_022_006, w_008_548);
  or2  I028_366(w_028_366, w_027_629, w_012_203);
  not1 I028_368(w_028_368, w_016_214);
  not1 I028_369(w_028_369, w_010_059);
  or2  I028_371(w_028_371, w_014_064, w_011_496);
  nand2 I028_376(w_028_376, w_015_397, w_017_001);
  not1 I028_397(w_028_397, w_024_336);
  nand2 I028_403(w_028_403, w_010_196, w_019_396);
  not1 I028_404(w_028_404, w_027_154);
  not1 I028_406(w_028_406, w_001_658);
  and2 I028_411(w_028_411, w_019_421, w_006_268);
  or2  I028_424(w_028_424, w_009_044, w_004_005);
  and2 I028_427(w_028_427, w_026_375, w_005_311);
  or2  I028_429(w_028_429, w_000_003, w_001_188);
  not1 I028_432(w_028_432, w_001_163);
  and2 I028_436(w_028_436, w_011_042, w_014_220);
  nand2 I028_439(w_028_439, w_008_642, w_016_260);
  not1 I028_440(w_028_440, w_024_229);
  nand2 I028_442(w_028_442, w_016_209, w_003_177);
  not1 I028_456(w_028_456, w_014_145);
  or2  I028_462(w_028_462, w_001_071, w_011_135);
  or2  I028_468(w_028_468, w_011_376, w_000_783);
  nand2 I028_470(w_028_470, w_025_012, w_013_009);
  nand2 I028_472(w_028_472, w_027_250, w_004_030);
  not1 I028_475(w_028_475, w_025_437);
  or2  I028_482(w_028_482, w_003_173, w_011_031);
  not1 I028_487(w_028_487, w_017_001);
  and2 I028_492(w_028_492, w_010_057, w_003_165);
  not1 I028_494(w_028_494, w_024_093);
  nand2 I028_496(w_028_496, w_019_074, w_004_036);
  and2 I028_506(w_028_506, w_010_117, w_022_149);
  nand2 I028_509(w_028_509, w_018_048, w_008_671);
  nand2 I028_511(w_028_511, w_027_486, w_017_018);
  and2 I028_527(w_028_527, w_003_210, w_022_008);
  and2 I028_535(w_028_535, w_027_115, w_021_169);
  not1 I028_544(w_028_544, w_021_305);
  nand2 I028_546(w_028_546, w_023_231, w_020_091);
  and2 I028_566(w_028_566, w_022_321, w_020_062);
  or2  I028_567(w_028_567, w_025_497, w_003_070);
  or2  I028_573(w_028_573, w_000_369, w_010_618);
  not1 I028_574(w_028_574, w_007_116);
  nand2 I028_577(w_028_577, w_009_012, w_007_418);
  and2 I028_581(w_028_581, w_001_297, w_004_010);
  not1 I028_590(w_028_590, w_015_559);
  nand2 I028_595(w_028_595, w_006_320, w_018_006);
  not1 I028_599(w_028_599, w_010_148);
  and2 I028_613(w_028_613, w_021_172, w_010_459);
  nand2 I028_615(w_028_615, w_016_162, w_026_295);
  nand2 I028_625(w_028_625, w_019_305, w_024_020);
  and2 I028_626(w_028_626, w_005_039, w_001_032);
  or2  I028_629(w_028_629, w_006_111, w_023_293);
  not1 I028_630(w_028_630, w_027_171);
  or2  I028_631(w_028_631, w_011_067, w_004_035);
  nand2 I028_638(w_028_638, w_012_405, w_026_283);
  not1 I028_647(w_028_647, w_017_023);
  nand2 I028_648(w_028_648, w_001_136, w_014_449);
  or2  I028_652(w_028_652, w_016_170, w_021_303);
  and2 I028_664(w_028_664, w_003_019, w_012_300);
  not1 I028_682(w_028_682, w_011_584);
  nand2 I028_693(w_028_693, w_008_658, w_024_452);
  nand2 I028_709(w_028_709, w_003_202, w_013_100);
  not1 I028_715(w_028_715, w_006_041);
  not1 I028_728(w_028_728, w_023_551);
  and2 I028_729(w_028_729, w_010_118, w_020_023);
  not1 I028_735(w_028_735, w_008_808);
  or2  I028_739(w_028_739, w_004_016, w_024_267);
  nand2 I028_745(w_028_745, w_010_088, w_020_134);
  or2  I028_762(w_028_762, w_021_003, w_015_024);
  not1 I028_764(w_028_764, w_014_341);
  and2 I028_767(w_028_767, w_016_313, w_010_719);
  nand2 I028_768(w_028_768, w_001_637, w_011_034);
  not1 I028_777(w_028_777, w_014_360);
  and2 I028_783(w_028_783, w_007_067, w_011_088);
  and2 I028_785(w_028_785, w_024_429, w_023_267);
  or2  I028_793(w_028_793, w_006_132, w_011_068);
  and2 I028_799(w_028_799, w_009_025, w_009_058);
  nand2 I028_811(w_028_811, w_007_356, w_002_139);
  nand2 I028_817(w_028_817, w_012_172, w_026_161);
  and2 I028_827(w_028_827, w_012_231, w_016_501);
  or2  I028_848(w_028_848, w_026_026, w_016_445);
  and2 I028_854(w_028_854, w_008_122, w_017_002);
  not1 I028_855(w_028_855, w_017_024);
  not1 I028_862(w_028_862, w_016_471);
  or2  I028_875(w_028_875, w_023_548, w_027_584);
  or2  I028_876(w_028_876, w_011_240, w_019_155);
  or2  I028_877(w_028_877, w_015_494, w_009_063);
  and2 I028_882(w_028_882, w_026_200, w_016_367);
  nand2 I028_885(w_028_885, w_027_663, w_026_096);
  or2  I028_886(w_028_886, w_010_449, w_004_013);
  not1 I028_890(w_028_890, w_024_257);
  nand2 I028_895(w_028_895, w_021_008, w_007_212);
  and2 I028_899(w_028_899, w_003_029, w_013_157);
  and2 I028_900(w_028_900, w_027_014, w_026_266);
  nand2 I029_004(w_029_004, w_015_201, w_012_406);
  nand2 I029_007(w_029_007, w_022_139, w_020_066);
  or2  I029_008(w_029_008, w_007_021, w_017_000);
  and2 I029_009(w_029_009, w_027_690, w_013_220);
  or2  I029_010(w_029_010, w_013_267, w_005_551);
  or2  I029_011(w_029_011, w_017_006, w_005_195);
  nand2 I029_016(w_029_016, w_001_446, w_028_799);
  or2  I029_020(w_029_020, w_003_167, w_018_117);
  or2  I029_021(w_029_021, w_009_009, w_011_667);
  nand2 I029_024(w_029_024, w_024_041, w_022_210);
  not1 I029_026(w_029_026, w_024_476);
  and2 I029_027(w_029_027, w_013_104, w_021_138);
  or2  I029_029(w_029_029, w_009_034, w_003_096);
  and2 I029_030(w_029_030, w_001_719, w_020_121);
  and2 I029_031(w_029_031, w_005_137, w_020_117);
  nand2 I029_034(w_029_034, w_028_566, w_023_181);
  and2 I029_035(w_029_035, w_015_178, w_019_100);
  or2  I029_036(w_029_036, w_015_648, w_021_008);
  and2 I029_038(w_029_038, w_007_095, w_001_601);
  or2  I029_039(w_029_039, w_027_165, w_018_155);
  or2  I029_040(w_029_040, w_007_190, w_022_032);
  nand2 I029_041(w_029_041, w_019_389, w_008_169);
  and2 I029_042(w_029_042, w_020_063, w_013_416);
  nand2 I029_044(w_029_044, w_021_191, w_019_322);
  nand2 I029_046(w_029_046, w_012_044, w_007_224);
  or2  I029_047(w_029_047, w_010_020, w_014_603);
  nand2 I029_050(w_029_050, w_009_059, w_020_119);
  and2 I029_051(w_029_051, w_002_081, w_015_155);
  or2  I029_054(w_029_054, w_005_009, w_022_006);
  or2  I029_056(w_029_056, w_004_020, w_003_197);
  and2 I029_061(w_029_061, w_026_236, w_014_181);
  not1 I029_062(w_029_062, w_017_023);
  nand2 I029_063(w_029_063, w_014_135, w_002_388);
  and2 I029_064(w_029_064, w_002_442, w_021_283);
  and2 I029_067(w_029_067, w_007_430, w_002_016);
  or2  I029_070(w_029_070, w_015_151, w_015_404);
  nand2 I029_071(w_029_071, w_009_018, w_008_411);
  and2 I029_072(w_029_072, w_017_006, w_017_020);
  or2  I029_073(w_029_073, w_002_453, w_021_162);
  not1 I029_075(w_029_075, w_012_301);
  or2  I029_077(w_029_077, w_001_700, w_028_432);
  not1 I029_080(w_029_080, w_000_033);
  not1 I029_082(w_029_082, w_007_336);
  nand2 I029_084(w_029_084, w_028_885, w_008_712);
  nand2 I029_086(w_029_086, w_013_441, w_025_406);
  nand2 I029_087(w_029_087, w_012_389, w_002_270);
  or2  I029_089(w_029_089, w_005_366, w_004_001);
  and2 I029_092(w_029_092, w_028_036, w_016_453);
  not1 I029_093(w_029_093, w_018_021);
  nand2 I029_094(w_029_094, w_020_092, w_028_328);
  nand2 I029_096(w_029_096, w_004_016, w_002_172);
  or2  I029_099(w_029_099, w_020_006, w_018_003);
  not1 I029_101(w_029_101, w_026_374);
  and2 I029_103(w_029_103, w_004_001, w_014_577);
  and2 I029_106(w_029_106, w_005_276, w_012_299);
  nand2 I029_110(w_029_110, w_007_509, w_007_123);
  or2  I029_111(w_029_111, w_003_215, w_020_024);
  nand2 I029_113(w_029_113, w_014_276, w_021_273);
  nand2 I029_114(w_029_114, w_026_056, w_007_390);
  and2 I029_115(w_029_115, w_001_700, w_015_594);
  and2 I029_116(w_029_116, w_022_344, w_011_449);
  nand2 I029_117(w_029_117, w_001_411, w_021_272);
  or2  I029_118(w_029_118, w_016_450, w_020_127);
  or2  I029_119(w_029_119, w_002_245, w_027_658);
  nand2 I029_120(w_029_120, w_018_103, w_026_252);
  not1 I029_123(w_029_123, w_020_012);
  not1 I029_124(w_029_124, w_021_328);
  and2 I029_125(w_029_125, w_006_139, w_014_213);
  nand2 I029_126(w_029_126, w_004_017, w_017_020);
  or2  I029_129(w_029_129, w_012_357, w_027_280);
  not1 I029_130(w_029_130, w_025_382);
  or2  I029_131(w_029_131, w_008_304, w_024_259);
  and2 I029_133(w_029_133, w_007_200, w_012_470);
  and2 I029_134(w_029_134, w_008_666, w_021_220);
  and2 I029_135(w_029_135, w_024_537, w_021_041);
  not1 I029_136(w_029_136, w_011_001);
  or2  I029_138(w_029_138, w_007_029, w_017_025);
  not1 I029_139(w_029_139, w_020_105);
  not1 I029_140(w_029_140, w_019_209);
  and2 I029_148(w_029_148, w_025_068, w_023_065);
  not1 I029_149(w_029_149, w_018_112);
  and2 I029_151(w_029_151, w_025_306, w_012_336);
  nand2 I029_154(w_029_154, w_011_023, w_010_086);
  and2 I029_157(w_029_157, w_010_583, w_004_016);
  nand2 I029_158(w_029_158, w_022_385, w_009_051);
  and2 I029_160(w_029_160, w_017_008, w_009_056);
  not1 I029_162(w_029_162, w_014_040);
  and2 I029_163(w_029_163, w_025_477, w_010_042);
  not1 I029_166(w_029_166, w_015_036);
  not1 I029_171(w_029_171, w_014_250);
  nand2 I029_173(w_029_173, w_007_390, w_015_611);
  nand2 I029_174(w_029_174, w_028_029, w_001_306);
  not1 I029_178(w_029_178, w_009_014);
  and2 I029_183(w_029_183, w_027_434, w_025_057);
  nand2 I029_186(w_029_186, w_001_095, w_002_142);
  not1 I029_187(w_029_187, w_021_016);
  nand2 I029_188(w_029_188, w_003_195, w_016_455);
  or2  I029_189(w_029_189, w_001_455, w_022_222);
  nand2 I029_190(w_029_190, w_012_008, w_024_309);
  not1 I029_191(w_029_191, w_016_400);
  not1 I029_192(w_029_192, w_000_769);
  and2 I029_193(w_029_193, w_012_416, w_003_147);
  and2 I029_196(w_029_196, w_024_326, w_016_397);
  and2 I029_199(w_029_199, w_000_613, w_007_299);
  nand2 I029_202(w_029_202, w_000_536, w_024_251);
  and2 I029_207(w_029_207, w_009_039, w_018_081);
  and2 I029_209(w_029_209, w_012_539, w_022_072);
  and2 I029_211(w_029_211, w_016_477, w_022_311);
  and2 I029_214(w_029_214, w_015_412, w_028_156);
  and2 I029_215(w_029_215, w_005_293, w_000_732);
  or2  I029_216(w_029_216, w_011_380, w_026_331);
  and2 I029_217(w_029_217, w_010_396, w_000_178);
  and2 I029_218(w_029_218, w_009_015, w_028_277);
  nand2 I030_001(w_030_001, w_006_026, w_001_551);
  and2 I030_002(w_030_002, w_007_387, w_015_277);
  and2 I030_003(w_030_003, w_015_196, w_005_103);
  or2  I030_004(w_030_004, w_020_104, w_025_042);
  not1 I030_005(w_030_005, w_006_324);
  not1 I030_010(w_030_010, w_001_665);
  nand2 I030_011(w_030_011, w_026_149, w_012_106);
  and2 I030_012(w_030_012, w_024_069, w_014_251);
  or2  I030_016(w_030_016, w_007_448, w_007_256);
  not1 I030_019(w_030_019, w_021_111);
  or2  I030_028(w_030_028, w_016_039, w_014_534);
  or2  I030_030(w_030_030, w_014_226, w_004_008);
  nand2 I030_031(w_030_031, w_029_160, w_002_063);
  and2 I030_033(w_030_033, w_000_657, w_021_183);
  nand2 I030_035(w_030_035, w_026_064, w_009_023);
  not1 I030_038(w_030_038, w_005_256);
  nand2 I030_041(w_030_041, w_008_100, w_027_267);
  not1 I030_044(w_030_044, w_004_022);
  and2 I030_045(w_030_045, w_022_406, w_019_042);
  nand2 I030_046(w_030_046, w_018_051, w_006_087);
  or2  I030_049(w_030_049, w_021_264, w_009_053);
  nand2 I030_050(w_030_050, w_018_119, w_011_353);
  nand2 I030_052(w_030_052, w_022_209, w_019_088);
  or2  I030_053(w_030_053, w_029_158, w_009_020);
  not1 I030_064(w_030_064, w_028_728);
  or2  I030_071(w_030_071, w_019_258, w_005_517);
  not1 I030_072(w_030_072, w_014_635);
  not1 I030_073(w_030_073, w_010_010);
  or2  I030_075(w_030_075, w_007_116, w_011_239);
  nand2 I030_076(w_030_076, w_008_231, w_028_202);
  and2 I030_080(w_030_080, w_026_080, w_029_116);
  or2  I030_082(w_030_082, w_025_159, w_008_685);
  nand2 I030_089(w_030_089, w_021_259, w_002_259);
  nand2 I030_105(w_030_105, w_022_421, w_023_239);
  and2 I030_109(w_030_109, w_014_228, w_016_054);
  nand2 I030_123(w_030_123, w_024_162, w_019_296);
  nand2 I030_133(w_030_133, w_023_053, w_029_029);
  or2  I030_145(w_030_145, w_013_010, w_023_569);
  not1 I030_149(w_030_149, w_029_134);
  not1 I030_151(w_030_151, w_029_075);
  and2 I030_152(w_030_152, w_008_347, w_016_442);
  not1 I030_158(w_030_158, w_023_038);
  not1 I030_160(w_030_160, w_018_134);
  nand2 I030_163(w_030_163, w_014_465, w_022_110);
  or2  I030_166(w_030_166, w_026_038, w_027_816);
  or2  I030_174(w_030_174, w_024_094, w_005_252);
  or2  I030_176(w_030_176, w_002_491, w_005_274);
  and2 I030_177(w_030_177, w_024_366, w_012_462);
  nand2 I030_178(w_030_178, w_008_652, w_027_168);
  or2  I030_182(w_030_182, w_028_131, w_001_133);
  or2  I030_184(w_030_184, w_008_268, w_023_305);
  nand2 I030_186(w_030_186, w_023_624, w_000_156);
  and2 I030_189(w_030_189, w_005_204, w_023_230);
  not1 I030_193(w_030_193, w_004_006);
  not1 I030_194(w_030_194, w_020_063);
  nand2 I030_196(w_030_196, w_003_165, w_014_073);
  nand2 I030_198(w_030_198, w_018_198, w_028_900);
  and2 I030_201(w_030_201, w_002_479, w_004_020);
  nand2 I030_202(w_030_202, w_002_298, w_002_207);
  or2  I030_203(w_030_203, w_009_011, w_000_366);
  or2  I030_205(w_030_205, w_003_093, w_027_663);
  and2 I030_206(w_030_206, w_001_218, w_014_127);
  not1 I030_210(w_030_210, w_021_341);
  nand2 I030_216(w_030_216, w_011_154, w_013_123);
  not1 I030_217(w_030_217, w_021_257);
  not1 I030_230(w_030_230, w_014_046);
  or2  I030_231(w_030_231, w_017_020, w_002_146);
  not1 I030_234(w_030_234, w_019_010);
  not1 I030_239(w_030_239, w_021_001);
  or2  I030_240(w_030_240, w_009_040, w_000_635);
  or2  I030_242(w_030_242, w_016_001, w_005_117);
  and2 I030_244(w_030_244, w_011_195, w_014_314);
  or2  I030_246(w_030_246, w_015_094, w_010_768);
  nand2 I030_247(w_030_247, w_011_222, w_011_337);
  and2 I030_248(w_030_248, w_014_259, w_027_130);
  nand2 I030_252(w_030_252, w_000_937, w_015_150);
  not1 I030_253(w_030_253, w_026_410);
  and2 I030_255(w_030_255, w_016_484, w_006_271);
  not1 I030_258(w_030_258, w_003_183);
  and2 I030_265(w_030_265, w_001_772, w_007_052);
  not1 I030_269(w_030_269, w_002_009);
  or2  I030_271(w_030_271, w_006_110, w_021_284);
  and2 I030_274(w_030_274, w_002_232, w_029_009);
  and2 I030_275(w_030_275, w_004_023, w_016_436);
  or2  I030_281(w_030_281, w_015_067, w_023_138);
  not1 I030_282(w_030_282, w_001_618);
  or2  I030_287(w_030_287, w_029_004, w_024_146);
  or2  I030_288(w_030_288, w_015_447, w_026_068);
  and2 I030_294(w_030_294, w_000_078, w_005_035);
  nand2 I030_305(w_030_305, w_027_373, w_003_073);
  nand2 I030_308(w_030_308, w_000_191, w_001_129);
  nand2 I030_311(w_030_311, w_025_195, w_004_022);
  and2 I030_312(w_030_312, w_007_553, w_006_293);
  and2 I030_314(w_030_314, w_018_141, w_007_199);
  and2 I030_318(w_030_318, w_025_239, w_008_689);
  not1 I030_324(w_030_324, w_019_279);
  nand2 I030_335(w_030_335, w_026_382, w_020_129);
  not1 I030_340(w_030_340, w_003_145);
  and2 I030_341(w_030_341, w_000_342, w_012_191);
  or2  I030_342(w_030_342, w_008_567, w_012_270);
  nand2 I030_347(w_030_347, w_011_092, w_011_090);
  or2  I030_353(w_030_353, w_020_112, w_002_483);
  nand2 I030_357(w_030_357, w_003_224, w_005_023);
  or2  I030_358(w_030_358, w_011_007, w_008_122);
  or2  I030_360(w_030_360, w_023_400, w_005_362);
  not1 I030_362(w_030_362, w_020_027);
  and2 I030_364(w_030_364, w_010_115, w_009_004);
  and2 I030_367(w_030_367, w_023_104, w_027_600);
  or2  I030_371(w_030_371, w_001_637, w_018_091);
  not1 I030_380(w_030_380, w_018_026);
  or2  I030_385(w_030_385, w_009_039, w_014_013);
  and2 I030_386(w_030_386, w_012_126, w_027_779);
  or2  I030_387(w_030_387, w_007_042, w_005_319);
  and2 I030_390(w_030_390, w_026_054, w_021_341);
  and2 I030_391(w_030_391, w_020_069, w_007_549);
  and2 I030_399(w_030_399, w_012_297, w_022_090);
  and2 I030_401(w_030_401, w_020_084, w_013_459);
  nand2 I030_405(w_030_405, w_028_682, w_008_230);
  nand2 I030_408(w_030_408, w_004_025, w_008_920);
  not1 I030_409(w_030_409, w_028_885);
  not1 I030_410(w_030_410, w_009_029);
  and2 I030_412(w_030_412, w_019_092, w_004_022);
  or2  I030_415(w_030_415, w_007_190, w_021_319);
  not1 I030_418(w_030_418, w_023_576);
  and2 I030_420(w_030_420, w_024_244, w_024_523);
  or2  I030_423(w_030_423, w_013_204, w_022_472);
  nand2 I030_424(w_030_424, w_011_288, w_010_646);
  and2 I030_433(w_030_433, w_019_265, w_026_024);
  or2  I030_435(w_030_435, w_022_244, w_007_004);
  or2  I030_438(w_030_438, w_014_021, w_021_243);
  or2  I030_444(w_030_444, w_011_556, w_017_009);
  or2  I030_445(w_030_445, w_000_582, w_024_293);
  nand2 I030_450(w_030_450, w_009_037, w_008_553);
  not1 I030_461(w_030_461, w_004_023);
  not1 I030_462(w_030_462, w_011_003);
  not1 I030_463(w_030_463, w_028_652);
  or2  I030_468(w_030_468, w_028_638, w_023_215);
  not1 I030_473(w_030_473, w_026_310);
  not1 I030_477(w_030_477, w_022_506);
  not1 I030_478(w_030_478, w_007_398);
  nand2 I030_480(w_030_480, w_006_207, w_029_123);
  or2  I030_481(w_030_481, w_011_433, w_005_342);
  or2  I030_483(w_030_483, w_025_223, w_000_445);
  not1 I030_484(w_030_484, w_027_600);
  nand2 I030_487(w_030_487, w_023_049, w_008_482);
  not1 I030_490(w_030_490, w_016_064);
  or2  I030_491(w_030_491, w_018_048, w_010_137);
  and2 I030_495(w_030_495, w_022_364, w_006_257);
  not1 I031_002(w_031_002, w_016_255);
  or2  I031_003(w_031_003, w_014_504, w_021_018);
  nand2 I031_004(w_031_004, w_005_026, w_012_544);
  nand2 I031_010(w_031_010, w_021_179, w_000_085);
  nand2 I031_011(w_031_011, w_003_008, w_004_005);
  not1 I031_015(w_031_015, w_004_024);
  and2 I031_016(w_031_016, w_011_253, w_017_002);
  or2  I031_017(w_031_017, w_015_227, w_022_432);
  nand2 I031_019(w_031_019, w_006_221, w_024_191);
  and2 I031_023(w_031_023, w_004_034, w_027_011);
  not1 I031_025(w_031_025, w_009_001);
  or2  I031_027(w_031_027, w_027_707, w_001_089);
  not1 I031_030(w_031_030, w_020_096);
  or2  I031_031(w_031_031, w_013_251, w_024_229);
  nand2 I031_035(w_031_035, w_000_967, w_004_029);
  not1 I031_043(w_031_043, w_011_370);
  or2  I031_045(w_031_045, w_008_759, w_012_193);
  and2 I031_050(w_031_050, w_006_297, w_028_296);
  or2  I031_055(w_031_055, w_011_063, w_030_405);
  nand2 I031_057(w_031_057, w_015_426, w_003_067);
  nand2 I031_071(w_031_071, w_004_010, w_029_089);
  nand2 I031_078(w_031_078, w_000_274, w_009_000);
  nand2 I031_082(w_031_082, w_013_268, w_023_108);
  or2  I031_085(w_031_085, w_020_098, w_026_274);
  and2 I031_087(w_031_087, w_013_417, w_001_632);
  not1 I031_089(w_031_089, w_009_013);
  nand2 I031_090(w_031_090, w_000_540, w_027_535);
  not1 I031_091(w_031_091, w_013_050);
  nand2 I031_094(w_031_094, w_007_265, w_022_101);
  or2  I031_095(w_031_095, w_007_411, w_020_107);
  not1 I031_103(w_031_103, w_025_108);
  nand2 I031_118(w_031_118, w_012_112, w_008_302);
  not1 I031_121(w_031_121, w_019_274);
  not1 I031_123(w_031_123, w_019_043);
  or2  I031_130(w_031_130, w_029_021, w_028_613);
  nand2 I031_135(w_031_135, w_005_028, w_020_063);
  or2  I031_150(w_031_150, w_020_063, w_003_123);
  or2  I031_154(w_031_154, w_003_193, w_006_249);
  and2 I031_161(w_031_161, w_023_448, w_003_178);
  or2  I031_167(w_031_167, w_025_346, w_020_035);
  not1 I031_171(w_031_171, w_007_015);
  not1 I031_178(w_031_178, w_002_150);
  nand2 I031_183(w_031_183, w_023_679, w_017_004);
  nand2 I031_187(w_031_187, w_026_376, w_020_071);
  not1 I031_194(w_031_194, w_027_401);
  not1 I031_196(w_031_196, w_022_383);
  not1 I031_198(w_031_198, w_001_020);
  nand2 I031_199(w_031_199, w_008_718, w_011_309);
  nand2 I031_204(w_031_204, w_018_130, w_010_095);
  or2  I031_210(w_031_210, w_003_179, w_026_125);
  and2 I031_211(w_031_211, w_005_276, w_010_240);
  or2  I031_212(w_031_212, w_000_383, w_021_353);
  or2  I031_215(w_031_215, w_020_033, w_023_071);
  nand2 I031_216(w_031_216, w_028_024, w_011_018);
  nand2 I031_219(w_031_219, w_028_631, w_015_112);
  or2  I031_224(w_031_224, w_011_309, w_016_219);
  nand2 I031_227(w_031_227, w_029_011, w_028_876);
  nand2 I031_229(w_031_229, w_025_223, w_000_692);
  nand2 I031_232(w_031_232, w_025_630, w_023_547);
  and2 I031_234(w_031_234, w_004_014, w_010_057);
  or2  I031_235(w_031_235, w_023_611, w_018_181);
  nand2 I031_240(w_031_240, w_022_067, w_003_066);
  not1 I031_241(w_031_241, w_011_133);
  nand2 I031_243(w_031_243, w_014_139, w_016_060);
  nand2 I031_244(w_031_244, w_014_035, w_014_183);
  and2 I031_246(w_031_246, w_000_744, w_003_048);
  nand2 I031_247(w_031_247, w_023_668, w_021_277);
  not1 I031_251(w_031_251, w_002_101);
  not1 I031_261(w_031_261, w_006_052);
  not1 I031_270(w_031_270, w_021_066);
  or2  I031_277(w_031_277, w_016_345, w_000_348);
  and2 I031_280(w_031_280, w_007_187, w_020_006);
  or2  I031_288(w_031_288, w_016_452, w_000_383);
  or2  I031_293(w_031_293, w_021_275, w_017_006);
  not1 I031_294(w_031_294, w_018_089);
  and2 I031_296(w_031_296, w_000_384, w_003_149);
  or2  I031_297(w_031_297, w_020_048, w_008_575);
  not1 I031_298(w_031_298, w_005_149);
  nand2 I031_299(w_031_299, w_010_570, w_029_075);
  or2  I031_302(w_031_302, w_027_672, w_025_131);
  and2 I031_303(w_031_303, w_028_764, w_008_690);
  and2 I031_306(w_031_306, w_025_015, w_003_084);
  nand2 I031_308(w_031_308, w_017_024, w_027_606);
  or2  I031_310(w_031_310, w_001_655, w_029_087);
  not1 I031_312(w_031_312, w_003_223);
  and2 I031_314(w_031_314, w_010_029, w_016_260);
  or2  I031_319(w_031_319, w_020_032, w_026_172);
  or2  I031_324(w_031_324, w_002_186, w_026_176);
  and2 I031_329(w_031_329, w_011_160, w_022_124);
  or2  I031_332(w_031_332, w_014_051, w_029_075);
  and2 I031_333(w_031_333, w_006_272, w_004_037);
  nand2 I031_340(w_031_340, w_019_319, w_029_188);
  or2  I031_345(w_031_345, w_014_346, w_012_093);
  nand2 I031_347(w_031_347, w_006_296, w_011_072);
  not1 I031_355(w_031_355, w_016_226);
  and2 I031_362(w_031_362, w_026_247, w_020_007);
  or2  I031_364(w_031_364, w_016_348, w_026_388);
  nand2 I031_365(w_031_365, w_018_192, w_024_266);
  nand2 I031_367(w_031_367, w_006_252, w_016_024);
  or2  I031_368(w_031_368, w_020_069, w_022_165);
  or2  I031_373(w_031_373, w_001_860, w_001_005);
  and2 I031_374(w_031_374, w_005_303, w_029_040);
  nand2 I031_382(w_031_382, w_023_295, w_001_307);
  or2  I031_391(w_031_391, w_030_030, w_006_034);
  or2  I031_399(w_031_399, w_005_338, w_026_295);
  not1 I031_406(w_031_406, w_014_351);
  and2 I031_409(w_031_409, w_003_148, w_030_269);
  and2 I031_410(w_031_410, w_021_024, w_012_531);
  not1 I031_413(w_031_413, w_014_186);
  and2 I031_420(w_031_420, w_029_162, w_019_259);
  and2 I031_421(w_031_421, w_023_468, w_022_457);
  or2  I031_438(w_031_438, w_000_708, w_004_008);
  nand2 I031_442(w_031_442, w_008_388, w_009_044);
  nand2 I031_443(w_031_443, w_003_163, w_012_299);
  and2 I031_446(w_031_446, w_014_228, w_009_003);
  nand2 I031_454(w_031_454, w_015_089, w_021_014);
  or2  I032_003(w_032_003, w_021_025, w_028_785);
  nand2 I032_007(w_032_007, w_018_051, w_026_297);
  or2  I032_010(w_032_010, w_030_075, w_003_001);
  nand2 I032_012(w_032_012, w_028_599, w_029_084);
  and2 I032_014(w_032_014, w_031_446, w_012_044);
  or2  I032_020(w_032_020, w_030_360, w_027_339);
  nand2 I032_023(w_032_023, w_028_648, w_027_087);
  and2 I032_031(w_032_031, w_026_340, w_019_040);
  nand2 I032_033(w_032_033, w_022_119, w_018_031);
  and2 I032_047(w_032_047, w_031_224, w_016_316);
  not1 I032_051(w_032_051, w_009_057);
  nand2 I032_057(w_032_057, w_005_417, w_026_365);
  nand2 I032_060(w_032_060, w_023_024, w_008_654);
  and2 I032_064(w_032_064, w_021_105, w_017_018);
  not1 I032_074(w_032_074, w_000_980);
  or2  I032_092(w_032_092, w_011_201, w_016_492);
  not1 I032_095(w_032_095, w_007_187);
  not1 I032_096(w_032_096, w_002_045);
  not1 I032_098(w_032_098, w_020_029);
  or2  I032_100(w_032_100, w_010_128, w_003_220);
  not1 I032_107(w_032_107, w_013_455);
  nand2 I032_113(w_032_113, w_020_058, w_029_163);
  or2  I032_116(w_032_116, w_029_202, w_016_137);
  not1 I032_119(w_032_119, w_027_336);
  not1 I032_121(w_032_121, w_015_368);
  and2 I032_124(w_032_124, w_002_363, w_030_433);
  and2 I032_126(w_032_126, w_022_275, w_008_030);
  or2  I032_127(w_032_127, w_026_065, w_004_028);
  or2  I032_130(w_032_130, w_007_375, w_022_337);
  or2  I032_144(w_032_144, w_028_241, w_018_069);
  and2 I032_146(w_032_146, w_004_005, w_018_108);
  nand2 I032_148(w_032_148, w_002_020, w_004_001);
  or2  I032_151(w_032_151, w_012_226, w_027_628);
  not1 I032_161(w_032_161, w_011_130);
  and2 I032_162(w_032_162, w_012_300, w_012_329);
  and2 I032_169(w_032_169, w_017_011, w_031_288);
  nand2 I032_170(w_032_170, w_030_409, w_022_097);
  and2 I032_175(w_032_175, w_030_035, w_010_058);
  and2 I032_178(w_032_178, w_002_126, w_018_102);
  and2 I032_179(w_032_179, w_007_165, w_031_078);
  and2 I032_180(w_032_180, w_002_208, w_020_046);
  or2  I032_187(w_032_187, w_017_009, w_026_294);
  nand2 I032_188(w_032_188, w_030_282, w_028_875);
  and2 I032_204(w_032_204, w_020_104, w_017_006);
  not1 I032_210(w_032_210, w_024_364);
  or2  I032_212(w_032_212, w_024_546, w_000_873);
  not1 I032_225(w_032_225, w_017_012);
  not1 I032_227(w_032_227, w_011_045);
  not1 I032_232(w_032_232, w_015_146);
  nand2 I032_233(w_032_233, w_000_485, w_014_451);
  and2 I032_234(w_032_234, w_025_169, w_017_000);
  or2  I032_237(w_032_237, w_030_201, w_022_267);
  and2 I032_238(w_032_238, w_020_038, w_010_260);
  or2  I032_259(w_032_259, w_013_073, w_019_403);
  not1 I032_267(w_032_267, w_026_407);
  not1 I032_268(w_032_268, w_000_803);
  or2  I032_289(w_032_289, w_021_328, w_000_511);
  nand2 I032_292(w_032_292, w_010_086, w_015_470);
  or2  I032_297(w_032_297, w_014_353, w_021_013);
  and2 I032_298(w_032_298, w_019_416, w_007_070);
  nand2 I032_307(w_032_307, w_014_124, w_024_238);
  nand2 I032_308(w_032_308, w_009_000, w_010_780);
  not1 I032_315(w_032_315, w_007_247);
  or2  I032_322(w_032_322, w_003_155, w_004_007);
  or2  I032_332(w_032_332, w_001_101, w_017_007);
  not1 I032_336(w_032_336, w_023_140);
  nand2 I032_347(w_032_347, w_028_020, w_022_210);
  nand2 I032_354(w_032_354, w_011_310, w_006_150);
  and2 I032_362(w_032_362, w_031_135, w_023_358);
  not1 I032_365(w_032_365, w_001_041);
  or2  I032_370(w_032_370, w_001_683, w_006_218);
  nand2 I032_372(w_032_372, w_002_326, w_004_009);
  not1 I032_376(w_032_376, w_009_029);
  or2  I032_378(w_032_378, w_022_323, w_005_174);
  not1 I032_380(w_032_380, w_013_309);
  nand2 I032_383(w_032_383, w_007_336, w_013_302);
  nand2 I032_397(w_032_397, w_025_591, w_027_353);
  nand2 I032_406(w_032_406, w_006_143, w_006_266);
  and2 I032_416(w_032_416, w_013_242, w_026_181);
  nand2 I032_421(w_032_421, w_021_259, w_019_146);
  not1 I032_424(w_032_424, w_002_476);
  and2 I032_449(w_032_449, w_027_085, w_011_624);
  not1 I032_454(w_032_454, w_009_006);
  not1 I032_455(w_032_455, w_017_020);
  or2  I032_466(w_032_466, w_024_334, w_007_005);
  not1 I032_477(w_032_477, w_020_049);
  not1 I032_498(w_032_498, w_005_400);
  nand2 I032_499(w_032_499, w_018_186, w_018_172);
  not1 I032_523(w_032_523, w_024_426);
  and2 I032_546(w_032_546, w_004_036, w_016_064);
  and2 I032_548(w_032_548, w_021_123, w_013_112);
  or2  I032_554(w_032_554, w_005_325, w_014_356);
  nand2 I032_556(w_032_556, w_023_274, w_022_294);
  or2  I032_570(w_032_570, w_009_008, w_002_133);
  or2  I032_585(w_032_585, w_013_281, w_031_089);
  and2 I032_588(w_032_588, w_002_257, w_025_233);
  not1 I032_591(w_032_591, w_013_381);
  not1 I032_593(w_032_593, w_023_241);
  not1 I032_594(w_032_594, w_029_073);
  not1 I032_596(w_032_596, w_010_641);
  or2  I032_602(w_032_602, w_025_147, w_012_441);
  and2 I032_603(w_032_603, w_022_433, w_008_779);
  or2  I032_636(w_032_636, w_012_474, w_028_436);
  or2  I032_649(w_032_649, w_000_140, w_031_374);
  nand2 I032_654(w_032_654, w_011_143, w_008_690);
  not1 I032_655(w_032_655, w_008_049);
  or2  I032_658(w_032_658, w_022_128, w_010_466);
  and2 I032_668(w_032_668, w_005_264, w_016_473);
  and2 I032_692(w_032_692, w_019_129, w_016_049);
  not1 I032_705(w_032_705, w_011_268);
  not1 I032_707(w_032_707, w_006_024);
  not1 I032_715(w_032_715, w_028_811);
  and2 I032_716(w_032_716, w_002_022, w_022_453);
  and2 I032_732(w_032_732, w_005_440, w_016_034);
  and2 I032_738(w_032_738, w_014_346, w_005_092);
  or2  I032_753(w_032_753, w_017_008, w_000_919);
  not1 I032_759(w_032_759, w_007_229);
  and2 I032_762(w_032_762, w_013_286, w_011_374);
  and2 I032_765(w_032_765, w_010_152, w_006_119);
  nand2 I032_777(w_032_777, w_029_044, w_017_022);
  or2  I032_778(w_032_778, w_013_031, w_014_141);
  or2  I032_790(w_032_790, w_020_052, w_010_125);
  nand2 I032_803(w_032_803, w_028_078, w_001_710);
  nand2 I032_804(w_032_804, w_028_313, w_009_021);
  or2  I032_807(w_032_807, w_009_055, w_029_196);
  not1 I032_810(w_032_810, w_000_568);
  nand2 I033_004(w_033_004, w_017_008, w_006_036);
  nand2 I033_006(w_033_006, w_001_581, w_024_034);
  nand2 I033_007(w_033_007, w_024_393, w_004_018);
  nand2 I033_011(w_033_011, w_018_030, w_016_052);
  nand2 I033_015(w_033_015, w_027_128, w_032_130);
  or2  I033_016(w_033_016, w_024_345, w_003_020);
  not1 I033_030(w_033_030, w_030_072);
  not1 I033_031(w_033_031, w_008_272);
  not1 I033_037(w_033_037, w_023_181);
  not1 I033_038(w_033_038, w_027_768);
  or2  I033_040(w_033_040, w_023_166, w_005_276);
  or2  I033_041(w_033_041, w_003_199, w_014_286);
  and2 I033_042(w_033_042, w_006_043, w_031_015);
  or2  I033_043(w_033_043, w_018_186, w_004_013);
  and2 I033_045(w_033_045, w_020_045, w_023_252);
  not1 I033_049(w_033_049, w_012_306);
  nand2 I033_050(w_033_050, w_010_339, w_019_024);
  nand2 I033_052(w_033_052, w_014_469, w_017_023);
  or2  I033_053(w_033_053, w_008_806, w_021_222);
  and2 I033_067(w_033_067, w_024_259, w_024_189);
  and2 I033_071(w_033_071, w_021_330, w_016_083);
  and2 I033_074(w_033_074, w_022_246, w_020_077);
  or2  I033_084(w_033_084, w_023_093, w_031_355);
  not1 I033_099(w_033_099, w_018_097);
  and2 I033_116(w_033_116, w_011_225, w_007_163);
  and2 I033_124(w_033_124, w_014_330, w_002_255);
  or2  I033_135(w_033_135, w_022_372, w_027_035);
  or2  I033_145(w_033_145, w_004_026, w_013_377);
  nand2 I033_174(w_033_174, w_017_002, w_013_319);
  nand2 I033_182(w_033_182, w_008_773, w_011_079);
  nand2 I033_190(w_033_190, w_025_068, w_005_256);
  and2 I033_192(w_033_192, w_010_278, w_007_423);
  not1 I033_193(w_033_193, w_031_089);
  nand2 I033_195(w_033_195, w_022_105, w_021_060);
  nand2 I033_196(w_033_196, w_009_031, w_006_210);
  not1 I033_202(w_033_202, w_025_033);
  not1 I033_208(w_033_208, w_013_457);
  and2 I033_210(w_033_210, w_008_534, w_006_078);
  or2  I033_218(w_033_218, w_025_654, w_000_358);
  or2  I033_221(w_033_221, w_008_073, w_021_219);
  nand2 I033_232(w_033_232, w_017_017, w_004_024);
  and2 I033_247(w_033_247, w_018_075, w_001_065);
  or2  I033_254(w_033_254, w_016_064, w_023_002);
  not1 I033_257(w_033_257, w_011_603);
  not1 I033_267(w_033_267, w_013_243);
  not1 I033_268(w_033_268, w_008_861);
  and2 I033_283(w_033_283, w_012_038, w_024_090);
  nand2 I033_294(w_033_294, w_029_020, w_027_257);
  or2  I033_296(w_033_296, w_003_013, w_032_376);
  nand2 I033_301(w_033_301, w_016_141, w_017_015);
  or2  I033_307(w_033_307, w_032_454, w_010_712);
  nand2 I033_311(w_033_311, w_032_023, w_016_125);
  nand2 I033_314(w_033_314, w_025_274, w_001_689);
  and2 I033_315(w_033_315, w_028_440, w_006_215);
  not1 I033_319(w_033_319, w_030_031);
  and2 I033_325(w_033_325, w_005_108, w_001_330);
  nand2 I033_326(w_033_326, w_006_296, w_021_137);
  nand2 I033_339(w_033_339, w_010_576, w_012_325);
  and2 I033_345(w_033_345, w_005_083, w_031_235);
  nand2 I033_352(w_033_352, w_029_111, w_026_108);
  nand2 I033_354(w_033_354, w_006_272, w_018_010);
  not1 I033_358(w_033_358, w_022_032);
  nand2 I033_361(w_033_361, w_008_437, w_010_551);
  nand2 I033_372(w_033_372, w_016_084, w_017_005);
  not1 I033_384(w_033_384, w_008_654);
  not1 I033_386(w_033_386, w_013_412);
  and2 I033_391(w_033_391, w_008_263, w_031_167);
  and2 I033_397(w_033_397, w_028_220, w_031_421);
  and2 I033_402(w_033_402, w_009_025, w_001_030);
  not1 I033_405(w_033_405, w_004_037);
  nand2 I033_406(w_033_406, w_022_054, w_020_118);
  nand2 I033_407(w_033_407, w_018_141, w_013_025);
  nand2 I033_414(w_033_414, w_005_346, w_007_249);
  or2  I033_416(w_033_416, w_005_066, w_008_118);
  not1 I033_420(w_033_420, w_026_247);
  and2 I033_428(w_033_428, w_001_378, w_025_003);
  nand2 I033_435(w_033_435, w_007_207, w_002_217);
  nand2 I033_437(w_033_437, w_002_214, w_023_240);
  nand2 I033_454(w_033_454, w_016_418, w_004_011);
  and2 I033_467(w_033_467, w_015_042, w_012_244);
  or2  I033_471(w_033_471, w_017_003, w_023_092);
  and2 I033_493(w_033_493, w_015_027, w_023_278);
  or2  I033_497(w_033_497, w_020_010, w_031_299);
  and2 I033_499(w_033_499, w_020_023, w_001_502);
  and2 I033_511(w_033_511, w_019_288, w_028_573);
  not1 I033_525(w_033_525, w_001_263);
  not1 I033_535(w_033_535, w_021_137);
  or2  I033_546(w_033_546, w_026_075, w_003_018);
  or2  I033_547(w_033_547, w_004_034, w_009_028);
  nand2 I033_548(w_033_548, w_018_157, w_021_045);
  nand2 I033_549(w_033_549, w_009_053, w_026_364);
  or2  I033_568(w_033_568, w_015_024, w_031_130);
  and2 I033_569(w_033_569, w_013_112, w_030_324);
  and2 I033_571(w_033_571, w_027_143, w_021_283);
  or2  I033_594(w_033_594, w_021_257, w_026_181);
  nand2 I033_597(w_033_597, w_011_317, w_017_016);
  not1 I033_598(w_033_598, w_022_046);
  and2 I033_601(w_033_601, w_003_103, w_006_004);
  not1 I033_610(w_033_610, w_011_535);
  or2  I033_613(w_033_613, w_021_342, w_022_161);
  nand2 I033_629(w_033_629, w_017_015, w_028_877);
  not1 I033_630(w_033_630, w_007_537);
  nand2 I033_645(w_033_645, w_008_702, w_015_608);
  and2 I033_675(w_033_675, w_015_585, w_007_345);
  not1 I033_679(w_033_679, w_015_493);
  nand2 I033_691(w_033_691, w_021_039, w_014_076);
  and2 I033_692(w_033_692, w_017_000, w_024_089);
  and2 I033_699(w_033_699, w_010_246, w_027_222);
  and2 I033_700(w_033_700, w_029_077, w_006_131);
  nand2 I033_709(w_033_709, w_025_246, w_000_968);
  and2 I033_718(w_033_718, w_001_195, w_001_543);
  or2  I033_721(w_033_721, w_003_008, w_005_008);
  nand2 I033_723(w_033_723, w_026_210, w_030_353);
  nand2 I033_726(w_033_726, w_025_202, w_006_101);
  nand2 I033_736(w_033_736, w_021_155, w_000_666);
  not1 I033_739(w_033_739, w_008_608);
  not1 I033_751(w_033_751, w_013_030);
  and2 I033_763(w_033_763, w_021_294, w_028_042);
  or2  I033_771(w_033_771, w_028_567, w_007_081);
  not1 I033_773(w_033_773, w_010_598);
  or2  I033_778(w_033_778, w_007_475, w_021_012);
  or2  I033_788(w_033_788, w_007_217, w_019_011);
  nand2 I033_805(w_033_805, w_023_013, w_014_479);
  nand2 I033_815(w_033_815, w_000_749, w_002_344);
  not1 I033_834(w_033_834, w_016_053);
  and2 I033_849(w_033_849, w_008_259, w_011_014);
  not1 I033_856(w_033_856, w_027_042);
  and2 I033_862(w_033_862, w_000_981, w_005_091);
  not1 I033_878(w_033_878, w_010_307);
  and2 I033_897(w_033_897, w_016_067, w_016_378);
  or2  I033_902(w_033_902, w_019_014, w_028_135);
  or2  I033_905(w_033_905, w_019_404, w_029_189);
  not1 I033_909(w_033_909, w_024_034);
  and2 I034_001(w_034_001, w_004_013, w_033_208);
  and2 I034_005(w_034_005, w_026_338, w_011_004);
  nand2 I034_012(w_034_012, w_011_281, w_017_002);
  or2  I034_013(w_034_013, w_002_172, w_005_154);
  and2 I034_018(w_034_018, w_033_815, w_002_229);
  nand2 I034_022(w_034_022, w_021_195, w_032_096);
  or2  I034_023(w_034_023, w_028_070, w_006_048);
  or2  I034_028(w_034_028, w_014_025, w_006_155);
  or2  I034_031(w_034_031, w_008_792, w_005_305);
  not1 I034_032(w_034_032, w_005_427);
  nand2 I034_033(w_034_033, w_011_355, w_011_110);
  and2 I034_034(w_034_034, w_013_002, w_008_423);
  and2 I034_041(w_034_041, w_008_155, w_011_437);
  or2  I034_042(w_034_042, w_016_038, w_033_084);
  and2 I034_043(w_034_043, w_013_034, w_015_592);
  or2  I034_044(w_034_044, w_030_076, w_009_039);
  or2  I034_045(w_034_045, w_011_657, w_026_400);
  or2  I034_054(w_034_054, w_015_098, w_027_208);
  and2 I034_060(w_034_060, w_027_189, w_010_113);
  not1 I034_063(w_034_063, w_010_049);
  nand2 I034_068(w_034_068, w_024_347, w_019_103);
  or2  I034_076(w_034_076, w_021_143, w_011_071);
  and2 I034_087(w_034_087, w_015_743, w_007_004);
  not1 I034_088(w_034_088, w_006_142);
  and2 I034_089(w_034_089, w_018_113, w_030_274);
  and2 I034_091(w_034_091, w_016_302, w_014_243);
  or2  I034_092(w_034_092, w_007_497, w_024_283);
  and2 I034_093(w_034_093, w_005_030, w_028_234);
  and2 I034_096(w_034_096, w_019_170, w_028_043);
  and2 I034_099(w_034_099, w_007_395, w_032_227);
  or2  I034_100(w_034_100, w_027_077, w_016_004);
  and2 I034_101(w_034_101, w_032_810, w_000_300);
  nand2 I034_103(w_034_103, w_029_124, w_015_619);
  nand2 I034_104(w_034_104, w_017_010, w_029_186);
  nand2 I034_113(w_034_113, w_027_699, w_022_320);
  nand2 I034_115(w_034_115, w_004_013, w_012_284);
  not1 I034_116(w_034_116, w_019_308);
  not1 I034_122(w_034_122, w_003_057);
  and2 I034_123(w_034_123, w_022_234, w_020_047);
  not1 I034_124(w_034_124, w_020_107);
  nand2 I034_127(w_034_127, w_032_074, w_018_156);
  or2  I034_130(w_034_130, w_022_352, w_009_032);
  not1 I034_136(w_034_136, w_032_289);
  not1 I034_137(w_034_137, w_019_025);
  nand2 I034_138(w_034_138, w_004_007, w_002_388);
  and2 I034_145(w_034_145, w_005_042, w_001_744);
  and2 I034_149(w_034_149, w_022_336, w_027_348);
  or2  I034_154(w_034_154, w_013_445, w_029_070);
  nand2 I034_160(w_034_160, w_001_096, w_014_595);
  or2  I034_164(w_034_164, w_013_142, w_011_026);
  nand2 I034_177(w_034_177, w_008_553, w_029_038);
  and2 I034_184(w_034_184, w_026_379, w_015_699);
  or2  I034_194(w_034_194, w_033_135, w_027_525);
  and2 I034_197(w_034_197, w_013_098, w_003_001);
  or2  I034_206(w_034_206, w_030_308, w_023_302);
  and2 I034_210(w_034_210, w_005_268, w_011_186);
  and2 I034_211(w_034_211, w_008_400, w_006_302);
  and2 I034_214(w_034_214, w_016_004, w_002_303);
  or2  I034_217(w_034_217, w_023_529, w_008_714);
  and2 I034_220(w_034_220, w_011_236, w_033_006);
  nand2 I034_227(w_034_227, w_004_028, w_002_289);
  or2  I034_234(w_034_234, w_010_547, w_031_194);
  nand2 I034_235(w_034_235, w_032_126, w_011_661);
  or2  I034_241(w_034_241, w_025_050, w_009_037);
  nand2 I034_242(w_034_242, w_028_326, w_028_028);
  or2  I034_250(w_034_250, w_008_899, w_011_192);
  nand2 I034_260(w_034_260, w_004_037, w_033_268);
  and2 I034_266(w_034_266, w_033_354, w_027_080);
  nand2 I034_270(w_034_270, w_001_674, w_033_116);
  or2  I034_296(w_034_296, w_028_735, w_013_321);
  nand2 I034_317(w_034_317, w_019_135, w_010_094);
  or2  I034_334(w_034_334, w_028_882, w_017_003);
  and2 I034_344(w_034_344, w_030_478, w_008_458);
  not1 I034_351(w_034_351, w_025_050);
  and2 I034_414(w_034_414, w_020_067, w_017_010);
  nand2 I034_422(w_034_422, w_010_070, w_011_420);
  or2  I034_429(w_034_429, w_014_222, w_008_154);
  not1 I034_431(w_034_431, w_018_111);
  not1 I034_433(w_034_433, w_003_164);
  nand2 I034_435(w_034_435, w_026_009, w_000_434);
  or2  I034_446(w_034_446, w_016_407, w_021_281);
  or2  I034_451(w_034_451, w_017_007, w_026_247);
  nand2 I034_458(w_034_458, w_003_040, w_017_022);
  not1 I034_478(w_034_478, w_011_093);
  nand2 I034_483(w_034_483, w_021_314, w_020_029);
  and2 I034_495(w_034_495, w_023_073, w_020_130);
  and2 I034_501(w_034_501, w_029_063, w_001_020);
  or2  I034_527(w_034_527, w_032_116, w_032_354);
  or2  I034_534(w_034_534, w_020_111, w_030_385);
  or2  I034_539(w_034_539, w_011_209, w_016_232);
  and2 I034_554(w_034_554, w_016_114, w_005_452);
  nand2 I034_555(w_034_555, w_031_373, w_011_159);
  or2  I034_567(w_034_567, w_020_104, w_028_817);
  not1 I034_573(w_034_573, w_002_074);
  nand2 I034_579(w_034_579, w_005_531, w_011_306);
  not1 I034_583(w_034_583, w_028_439);
  or2  I034_588(w_034_588, w_001_356, w_008_780);
  not1 I034_596(w_034_596, w_018_141);
  nand2 I034_618(w_034_618, w_019_219, w_006_150);
  or2  I034_640(w_034_640, w_020_046, w_030_491);
  and2 I034_666(w_034_666, w_029_047, w_020_137);
  not1 I034_672(w_034_672, w_033_296);
  nand2 I034_681(w_034_681, w_002_309, w_014_464);
  nand2 I034_684(w_034_684, w_023_670, w_006_246);
  not1 I034_691(w_034_691, w_032_602);
  or2  I034_693(w_034_693, w_028_442, w_010_197);
  not1 I034_721(w_034_721, w_021_283);
  not1 I034_725(w_034_725, w_006_230);
  nand2 I034_729(w_034_729, w_023_138, w_010_123);
  or2  I034_775(w_034_775, w_013_281, w_013_353);
  and2 I034_785(w_034_785, w_013_249, w_022_057);
  nand2 I034_792(w_034_792, w_014_163, w_023_175);
  and2 I034_798(w_034_798, w_004_031, w_013_017);
  or2  I034_801(w_034_801, w_019_072, w_027_080);
  and2 I034_805(w_034_805, w_030_239, w_002_210);
  not1 I034_806(w_034_806, w_025_542);
  or2  I035_003(w_035_003, w_032_148, w_029_118);
  nand2 I035_006(w_035_006, w_032_297, w_021_045);
  or2  I035_009(w_035_009, w_034_640, w_026_058);
  and2 I035_015(w_035_015, w_017_017, w_009_014);
  not1 I035_024(w_035_024, w_022_159);
  not1 I035_025(w_035_025, w_012_423);
  not1 I035_032(w_035_032, w_017_016);
  or2  I035_041(w_035_041, w_018_104, w_029_149);
  or2  I035_051(w_035_051, w_029_086, w_003_048);
  or2  I035_054(w_035_054, w_007_089, w_007_163);
  not1 I035_072(w_035_072, w_013_428);
  not1 I035_074(w_035_074, w_026_007);
  or2  I035_078(w_035_078, w_019_185, w_000_129);
  and2 I035_081(w_035_081, w_009_032, w_031_123);
  not1 I035_083(w_035_083, w_033_679);
  not1 I035_089(w_035_089, w_026_091);
  and2 I035_092(w_035_092, w_017_004, w_004_033);
  nand2 I035_102(w_035_102, w_022_073, w_017_017);
  not1 I035_114(w_035_114, w_021_352);
  not1 I035_120(w_035_120, w_009_014);
  not1 I035_121(w_035_121, w_009_018);
  or2  I035_127(w_035_127, w_015_011, w_030_046);
  and2 I035_129(w_035_129, w_000_697, w_009_046);
  and2 I035_132(w_035_132, w_021_070, w_015_689);
  nand2 I035_134(w_035_134, w_033_174, w_002_360);
  not1 I035_135(w_035_135, w_025_153);
  nand2 I035_142(w_035_142, w_000_970, w_033_535);
  or2  I035_145(w_035_145, w_011_254, w_027_054);
  or2  I035_150(w_035_150, w_034_013, w_032_007);
  or2  I035_152(w_035_152, w_003_122, w_025_233);
  or2  I035_156(w_035_156, w_029_148, w_018_081);
  not1 I035_160(w_035_160, w_017_016);
  nand2 I035_163(w_035_163, w_028_218, w_016_065);
  not1 I035_167(w_035_167, w_014_180);
  and2 I035_169(w_035_169, w_010_065, w_000_555);
  not1 I035_170(w_035_170, w_027_234);
  and2 I035_179(w_035_179, w_011_564, w_004_038);
  nand2 I035_184(w_035_184, w_002_188, w_000_714);
  or2  I035_191(w_035_191, w_027_429, w_004_015);
  or2  I035_192(w_035_192, w_004_001, w_001_524);
  or2  I035_195(w_035_195, w_031_364, w_002_457);
  or2  I035_199(w_035_199, w_012_167, w_012_385);
  and2 I035_212(w_035_212, w_010_054, w_016_225);
  or2  I035_214(w_035_214, w_000_832, w_031_229);
  or2  I035_220(w_035_220, w_006_226, w_029_218);
  or2  I035_225(w_035_225, w_026_305, w_026_399);
  or2  I035_230(w_035_230, w_005_121, w_029_010);
  nand2 I035_245(w_035_245, w_014_237, w_006_274);
  not1 I035_258(w_035_258, w_025_294);
  and2 I035_261(w_035_261, w_005_113, w_008_497);
  and2 I035_265(w_035_265, w_034_351, w_034_130);
  nand2 I035_268(w_035_268, w_028_087, w_032_031);
  or2  I035_274(w_035_274, w_022_281, w_019_230);
  not1 I035_277(w_035_277, w_003_132);
  not1 I035_286(w_035_286, w_004_018);
  nand2 I035_292(w_035_292, w_029_118, w_007_053);
  and2 I035_297(w_035_297, w_005_031, w_012_435);
  not1 I035_304(w_035_304, w_007_275);
  and2 I035_307(w_035_307, w_002_294, w_005_288);
  or2  I035_313(w_035_313, w_012_434, w_006_262);
  not1 I035_323(w_035_323, w_027_177);
  nand2 I035_324(w_035_324, w_017_011, w_033_736);
  or2  I035_326(w_035_326, w_032_466, w_009_055);
  not1 I035_335(w_035_335, w_023_137);
  and2 I035_346(w_035_346, w_002_248, w_033_016);
  or2  I035_351(w_035_351, w_009_024, w_012_137);
  not1 I035_370(w_035_370, w_032_594);
  not1 I035_374(w_035_374, w_031_329);
  not1 I035_382(w_035_382, w_017_004);
  or2  I035_397(w_035_397, w_025_510, w_024_495);
  not1 I035_400(w_035_400, w_022_276);
  nand2 I035_415(w_035_415, w_028_076, w_031_347);
  not1 I035_429(w_035_429, w_008_215);
  not1 I035_460(w_035_460, w_006_274);
  nand2 I035_467(w_035_467, w_007_076, w_023_269);
  nand2 I035_473(w_035_473, w_034_012, w_010_414);
  or2  I035_479(w_035_479, w_013_209, w_010_111);
  nand2 I035_480(w_035_480, w_032_362, w_024_267);
  or2  I035_487(w_035_487, w_022_105, w_014_235);
  nand2 I035_492(w_035_492, w_000_739, w_034_234);
  and2 I035_518(w_035_518, w_007_438, w_008_840);
  and2 I035_524(w_035_524, w_016_040, w_024_192);
  not1 I035_527(w_035_527, w_007_083);
  nand2 I035_532(w_035_532, w_020_042, w_001_083);
  or2  I035_535(w_035_535, w_033_319, w_017_006);
  nand2 I035_539(w_035_539, w_003_046, w_032_051);
  or2  I035_540(w_035_540, w_008_129, w_014_306);
  nand2 I035_554(w_035_554, w_026_308, w_011_141);
  and2 I035_563(w_035_563, w_015_760, w_030_438);
  nand2 I035_574(w_035_574, w_002_000, w_029_101);
  not1 I035_578(w_035_578, w_008_629);
  not1 I035_588(w_035_588, w_014_162);
  or2  I035_592(w_035_592, w_018_190, w_013_128);
  or2  I035_598(w_035_598, w_032_010, w_018_084);
  or2  I035_607(w_035_607, w_030_041, w_025_308);
  not1 I035_612(w_035_612, w_001_182);
  or2  I035_616(w_035_616, w_008_077, w_012_166);
  nand2 I035_622(w_035_622, w_007_552, w_025_183);
  not1 I035_629(w_035_629, w_021_157);
  nand2 I035_631(w_035_631, w_013_239, w_000_982);
  nand2 I035_633(w_035_633, w_012_026, w_025_232);
  not1 I035_650(w_035_652, w_035_651);
  or2  I035_651(w_035_653, w_008_613, w_035_652);
  and2 I035_652(w_035_654, w_035_653, w_016_370);
  and2 I035_653(w_035_655, w_017_002, w_035_654);
  and2 I035_654(w_035_656, w_035_655, w_002_110);
  and2 I035_655(w_035_657, w_030_166, w_035_656);
  nand2 I035_656(w_035_658, w_035_657, w_001_666);
  not1 I035_657(w_035_659, w_035_658);
  and2 I035_658(w_035_660, w_008_746, w_035_659);
  or2  I035_659(w_035_651, w_007_437, w_035_660);
  and2 I036_005(w_036_005, w_034_005, w_015_037);
  nand2 I036_008(w_036_008, w_033_699, w_019_165);
  not1 I036_009(w_036_009, w_023_136);
  not1 I036_013(w_036_013, w_011_025);
  or2  I036_016(w_036_016, w_029_035, w_034_227);
  nand2 I036_018(w_036_018, w_035_429, w_010_037);
  or2  I036_019(w_036_019, w_026_361, w_031_443);
  or2  I036_021(w_036_021, w_011_261, w_005_297);
  or2  I036_023(w_036_023, w_027_172, w_019_279);
  or2  I036_031(w_036_031, w_024_194, w_020_086);
  and2 I036_036(w_036_036, w_025_160, w_010_208);
  not1 I036_040(w_036_040, w_012_426);
  nand2 I036_042(w_036_042, w_022_100, w_002_340);
  and2 I036_043(w_036_043, w_004_011, w_025_022);
  not1 I036_046(w_036_046, w_004_021);
  or2  I036_052(w_036_052, w_030_357, w_025_454);
  and2 I036_056(w_036_056, w_013_172, w_015_170);
  not1 I036_061(w_036_061, w_026_012);
  not1 I036_066(w_036_066, w_003_010);
  and2 I036_068(w_036_068, w_023_444, w_010_012);
  not1 I036_069(w_036_069, w_022_144);
  and2 I036_070(w_036_070, w_020_112, w_014_058);
  nand2 I036_071(w_036_071, w_028_482, w_002_001);
  not1 I036_073(w_036_073, w_012_299);
  not1 I036_080(w_036_080, w_002_021);
  nand2 I036_082(w_036_082, w_015_714, w_015_669);
  and2 I036_084(w_036_084, w_020_041, w_018_129);
  or2  I036_085(w_036_085, w_007_350, w_034_194);
  or2  I036_089(w_036_089, w_033_568, w_026_046);
  nand2 I036_090(w_036_090, w_006_185, w_016_211);
  nand2 I036_092(w_036_092, w_016_113, w_028_027);
  and2 I036_093(w_036_093, w_007_115, w_016_471);
  nand2 I036_095(w_036_095, w_023_387, w_015_206);
  or2  I036_097(w_036_097, w_013_399, w_002_303);
  not1 I036_102(w_036_102, w_003_057);
  and2 I036_103(w_036_103, w_021_164, w_027_776);
  nand2 I036_105(w_036_105, w_008_246, w_026_095);
  or2  I036_111(w_036_111, w_028_132, w_016_452);
  not1 I036_112(w_036_112, w_024_276);
  and2 I036_113(w_036_113, w_016_050, w_012_204);
  not1 I036_115(w_036_115, w_022_503);
  or2  I036_122(w_036_122, w_032_127, w_010_211);
  nand2 I036_123(w_036_123, w_006_195, w_012_318);
  and2 I036_125(w_036_125, w_030_005, w_031_413);
  or2  I036_131(w_036_131, w_028_615, w_003_158);
  nand2 I036_132(w_036_132, w_013_012, w_010_591);
  not1 I036_134(w_036_134, w_001_038);
  or2  I036_138(w_036_138, w_032_804, w_030_435);
  not1 I036_143(w_036_143, w_018_126);
  or2  I036_145(w_036_145, w_028_745, w_029_129);
  and2 I036_146(w_036_146, w_030_217, w_009_056);
  nand2 I036_147(w_036_147, w_027_412, w_018_057);
  and2 I036_149(w_036_149, w_003_061, w_023_109);
  nand2 I036_151(w_036_151, w_017_000, w_004_038);
  nand2 I036_153(w_036_153, w_002_110, w_002_012);
  not1 I036_154(w_036_154, w_020_137);
  and2 I036_156(w_036_156, w_029_050, w_023_359);
  and2 I036_158(w_036_158, w_006_109, w_008_863);
  not1 I036_166(w_036_166, w_019_102);
  not1 I036_171(w_036_171, w_011_257);
  or2  I036_175(w_036_175, w_033_405, w_030_380);
  or2  I036_177(w_036_177, w_021_181, w_024_244);
  not1 I036_185(w_036_185, w_015_629);
  and2 I036_193(w_036_193, w_028_161, w_025_297);
  not1 I036_197(w_036_197, w_017_009);
  or2  I036_199(w_036_199, w_021_158, w_021_248);
  or2  I036_201(w_036_201, w_014_020, w_019_310);
  or2  I036_205(w_036_205, w_018_194, w_013_133);
  or2  I036_209(w_036_209, w_011_526, w_011_050);
  not1 I036_217(w_036_217, w_031_210);
  and2 I036_222(w_036_222, w_035_346, w_002_355);
  or2  I036_228(w_036_228, w_033_386, w_013_480);
  and2 I036_233(w_036_233, w_016_318, w_022_155);
  or2  I036_234(w_036_234, w_027_055, w_026_249);
  not1 I036_237(w_036_237, w_009_065);
  and2 I036_238(w_036_238, w_002_491, w_011_225);
  and2 I036_239(w_036_239, w_025_465, w_008_893);
  not1 I036_247(w_036_247, w_007_287);
  and2 I036_249(w_036_249, w_025_554, w_003_110);
  not1 I036_260(w_036_260, w_007_369);
  or2  I036_262(w_036_262, w_009_027, w_002_168);
  not1 I036_266(w_036_266, w_017_017);
  or2  I036_271(w_036_271, w_009_009, w_020_020);
  and2 I036_273(w_036_273, w_031_362, w_009_024);
  or2  I036_276(w_036_276, w_020_006, w_027_343);
  and2 I036_277(w_036_277, w_023_197, w_011_336);
  not1 I036_278(w_036_278, w_000_105);
  and2 I036_282(w_036_282, w_034_043, w_017_006);
  nand2 I036_283(w_036_283, w_025_658, w_035_170);
  nand2 I036_284(w_036_286, w_004_009, w_036_285);
  nand2 I036_285(w_036_287, w_035_274, w_036_286);
  and2 I036_286(w_036_288, w_036_287, w_028_281);
  nand2 I036_287(w_036_289, w_036_288, w_001_264);
  or2  I036_288(w_036_290, w_016_370, w_036_289);
  and2 I036_289(w_036_285, w_036_290, w_026_361);
  not1 I037_000(w_037_000, w_016_181);
  nand2 I037_001(w_037_001, w_026_100, w_002_302);
  or2  I037_004(w_037_004, w_029_118, w_020_064);
  or2  I037_005(w_037_005, w_020_122, w_029_209);
  nand2 I037_006(w_037_006, w_011_267, w_029_071);
  or2  I037_008(w_037_008, w_013_437, w_021_044);
  or2  I037_009(w_037_009, w_008_517, w_033_232);
  not1 I037_011(w_037_011, w_007_177);
  nand2 I037_012(w_037_012, w_005_112, w_011_678);
  not1 I037_013(w_037_013, w_023_253);
  or2  I037_014(w_037_014, w_018_008, w_008_898);
  not1 I037_016(w_037_016, w_031_240);
  not1 I037_017(w_037_017, w_006_205);
  not1 I037_019(w_037_019, w_014_474);
  and2 I037_020(w_037_020, w_035_167, w_002_284);
  not1 I037_022(w_037_022, w_010_311);
  or2  I037_024(w_037_024, w_035_163, w_020_067);
  or2  I037_025(w_037_025, w_013_016, w_009_056);
  not1 I037_026(w_037_026, w_001_531);
  not1 I037_027(w_037_027, w_000_700);
  not1 I037_032(w_037_032, w_005_574);
  or2  I037_036(w_037_036, w_008_734, w_027_207);
  and2 I037_039(w_037_039, w_013_259, w_020_073);
  nand2 I037_040(w_037_040, w_028_222, w_026_307);
  and2 I037_041(w_037_041, w_018_038, w_036_132);
  or2  I037_043(w_037_043, w_036_149, w_028_206);
  and2 I037_047(w_037_047, w_004_015, w_024_473);
  or2  I037_049(w_037_049, w_031_345, w_026_139);
  and2 I037_051(w_037_051, w_035_479, w_006_214);
  not1 I037_052(w_037_052, w_011_361);
  not1 I037_055(w_037_055, w_028_827);
  nand2 I037_061(w_037_061, w_030_463, w_022_286);
  and2 I037_063(w_037_063, w_019_021, w_019_347);
  or2  I037_064(w_037_064, w_001_207, w_028_581);
  or2  I037_066(w_037_066, w_006_000, w_028_004);
  not1 I037_067(w_037_067, w_028_371);
  and2 I037_070(w_037_070, w_031_299, w_020_126);
  nand2 I037_073(w_037_073, w_004_015, w_023_177);
  nand2 I037_074(w_037_074, w_014_241, w_036_154);
  not1 I037_076(w_037_076, w_022_402);
  nand2 I037_077(w_037_077, w_017_001, w_027_114);
  not1 I037_079(w_037_079, w_007_187);
  or2  I037_081(w_037_081, w_029_084, w_000_752);
  and2 I037_085(w_037_085, w_028_793, w_028_294);
  not1 I037_090(w_037_090, w_024_029);
  nand2 I037_091(w_037_091, w_013_037, w_021_221);
  and2 I037_095(w_037_095, w_012_177, w_005_412);
  or2  I037_096(w_037_096, w_014_157, w_022_519);
  nand2 I037_097(w_037_097, w_024_496, w_020_091);
  not1 I037_098(w_037_098, w_005_141);
  or2  I037_099(w_037_099, w_036_070, w_033_283);
  or2  I037_103(w_037_103, w_022_162, w_004_007);
  nand2 I037_105(w_037_105, w_016_062, w_009_006);
  nand2 I037_106(w_037_106, w_001_087, w_030_189);
  not1 I037_107(w_037_107, w_016_028);
  or2  I037_109(w_037_109, w_027_087, w_020_027);
  and2 I037_111(w_037_111, w_028_128, w_008_922);
  and2 I037_112(w_037_112, w_032_178, w_032_707);
  or2  I037_113(w_037_113, w_003_022, w_014_043);
  and2 I037_114(w_037_114, w_022_426, w_035_467);
  nand2 I037_115(w_037_115, w_028_246, w_032_372);
  not1 I037_116(w_037_116, w_027_431);
  nand2 I037_119(w_037_119, w_034_478, w_024_364);
  or2  I037_122(w_037_122, w_030_011, w_007_027);
  nand2 I037_124(w_037_124, w_005_002, w_020_025);
  and2 I037_127(w_037_127, w_023_470, w_016_003);
  and2 I037_128(w_037_128, w_018_019, w_002_073);
  or2  I037_130(w_037_130, w_008_116, w_030_265);
  not1 I037_131(w_037_131, w_013_298);
  or2  I037_133(w_037_133, w_033_195, w_017_006);
  or2  I037_140(w_037_140, w_017_010, w_023_520);
  and2 I037_141(w_037_141, w_020_123, w_029_047);
  nand2 I037_142(w_037_142, w_000_277, w_028_258);
  not1 I037_145(w_037_145, w_015_191);
  nand2 I037_147(w_037_147, w_016_367, w_010_002);
  not1 I037_148(w_037_148, w_002_052);
  not1 I037_149(w_037_149, w_017_011);
  nand2 I037_152(w_037_152, w_029_216, w_006_022);
  nand2 I037_154(w_037_154, w_026_388, w_006_023);
  and2 I037_162(w_037_162, w_021_026, w_032_759);
  or2  I037_163(w_037_163, w_007_313, w_034_124);
  and2 I037_164(w_037_164, w_005_281, w_029_062);
  and2 I037_165(w_037_165, w_024_225, w_035_480);
  not1 I037_171(w_037_171, w_015_052);
  and2 I037_176(w_037_176, w_027_075, w_012_384);
  not1 I037_180(w_037_180, w_019_299);
  and2 I037_183(w_037_183, w_016_466, w_030_364);
  not1 I037_187(w_037_187, w_005_132);
  nand2 I037_189(w_037_189, w_033_525, w_002_186);
  and2 I037_190(w_037_190, w_031_198, w_004_020);
  not1 I038_009(w_038_009, w_005_045);
  and2 I038_012(w_038_012, w_005_185, w_028_359);
  and2 I038_015(w_038_015, w_007_238, w_024_316);
  not1 I038_028(w_038_028, w_020_002);
  and2 I038_031(w_038_031, w_033_405, w_009_024);
  and2 I038_035(w_038_035, w_011_065, w_016_221);
  not1 I038_037(w_038_037, w_031_261);
  nand2 I038_038(w_038_038, w_002_437, w_012_003);
  nand2 I038_041(w_038_041, w_021_201, w_021_120);
  and2 I038_046(w_038_046, w_025_347, w_021_314);
  and2 I038_047(w_038_047, w_014_311, w_015_538);
  not1 I038_049(w_038_049, w_019_068);
  and2 I038_050(w_038_050, w_023_457, w_030_386);
  and2 I038_057(w_038_057, w_029_166, w_030_205);
  and2 I038_094(w_038_094, w_021_079, w_018_129);
  or2  I038_101(w_038_101, w_008_411, w_021_048);
  nand2 I038_114(w_038_114, w_024_000, w_010_157);
  nand2 I038_117(w_038_117, w_030_481, w_016_387);
  or2  I038_118(w_038_118, w_000_624, w_020_008);
  nand2 I038_119(w_038_119, w_024_133, w_015_345);
  not1 I038_122(w_038_122, w_015_166);
  nand2 I038_123(w_038_123, w_037_127, w_034_041);
  nand2 I038_135(w_038_135, w_006_024, w_030_410);
  and2 I038_148(w_038_148, w_030_253, w_035_304);
  nand2 I038_149(w_038_149, w_037_019, w_022_026);
  and2 I038_156(w_038_156, w_017_021, w_017_008);
  or2  I038_157(w_038_157, w_015_021, w_002_346);
  nand2 I038_168(w_038_168, w_028_081, w_017_017);
  nand2 I038_172(w_038_172, w_002_417, w_000_182);
  and2 I038_173(w_038_173, w_028_043, w_015_418);
  nand2 I038_177(w_038_177, w_012_371, w_016_276);
  nand2 I038_180(w_038_180, w_025_093, w_030_003);
  and2 I038_186(w_038_186, w_025_018, w_027_794);
  or2  I038_188(w_038_188, w_026_110, w_035_199);
  or2  I038_190(w_038_190, w_013_300, w_037_190);
  or2  I038_194(w_038_194, w_013_003, w_013_090);
  nand2 I038_202(w_038_202, w_028_487, w_001_443);
  not1 I038_206(w_038_206, w_017_008);
  and2 I038_224(w_038_224, w_010_596, w_009_041);
  nand2 I038_227(w_038_227, w_011_458, w_032_347);
  and2 I038_235(w_038_235, w_032_365, w_016_021);
  or2  I038_238(w_038_238, w_006_257, w_004_005);
  or2  I038_277(w_038_277, w_004_021, w_023_352);
  and2 I038_303(w_038_303, w_014_434, w_034_666);
  or2  I038_305(w_038_305, w_008_514, w_026_048);
  and2 I038_324(w_038_324, w_024_455, w_015_476);
  nand2 I038_335(w_038_335, w_000_163, w_012_338);
  nand2 I038_345(w_038_345, w_019_101, w_010_359);
  or2  I038_388(w_038_388, w_016_191, w_024_037);
  or2  I038_413(w_038_413, w_036_102, w_006_031);
  not1 I038_432(w_038_432, w_026_393);
  nand2 I038_447(w_038_447, w_022_049, w_028_475);
  not1 I038_448(w_038_448, w_011_137);
  or2  I038_459(w_038_459, w_034_022, w_005_114);
  or2  I038_469(w_038_469, w_015_314, w_020_083);
  or2  I038_489(w_038_489, w_036_158, w_003_086);
  not1 I038_521(w_038_521, w_029_039);
  not1 I038_526(w_038_526, w_022_169);
  and2 I038_543(w_038_543, w_022_516, w_004_019);
  not1 I038_548(w_038_548, w_001_259);
  and2 I038_559(w_038_559, w_033_099, w_032_397);
  nand2 I038_560(w_038_560, w_019_248, w_024_307);
  nand2 I038_562(w_038_562, w_015_138, w_036_070);
  not1 I038_565(w_038_565, w_001_482);
  or2  I038_573(w_038_573, w_020_098, w_025_115);
  or2  I038_591(w_038_591, w_024_103, w_013_325);
  and2 I038_612(w_038_612, w_012_535, w_011_006);
  nand2 I038_621(w_038_621, w_026_039, w_015_146);
  and2 I038_625(w_038_625, w_031_043, w_023_472);
  nand2 I038_637(w_038_637, w_021_039, w_001_820);
  not1 I038_640(w_038_640, w_019_051);
  not1 I038_644(w_038_644, w_030_255);
  and2 I038_648(w_038_648, w_024_343, w_012_010);
  nand2 I038_665(w_038_665, w_032_074, w_025_011);
  and2 I038_689(w_038_689, w_013_479, w_031_229);
  not1 I038_694(w_038_694, w_000_983);
  not1 I038_696(w_038_696, w_007_428);
  or2  I038_701(w_038_701, w_021_084, w_003_093);
  and2 I038_709(w_038_709, w_023_513, w_014_542);
  or2  I038_713(w_038_713, w_025_275, w_013_466);
  and2 I038_735(w_038_735, w_024_560, w_027_478);
  not1 I038_747(w_038_747, w_007_319);
  not1 I038_748(w_038_748, w_002_317);
  and2 I038_762(w_038_762, w_026_226, w_021_159);
  or2  I038_764(w_038_764, w_027_624, w_011_232);
  and2 I039_002(w_039_002, w_015_442, w_015_117);
  nand2 I039_003(w_039_003, w_014_188, w_019_335);
  or2  I039_005(w_039_005, w_003_075, w_022_117);
  not1 I039_007(w_039_007, w_010_550);
  not1 I039_008(w_039_008, w_006_229);
  and2 I039_010(w_039_010, w_030_468, w_013_078);
  and2 I039_013(w_039_013, w_025_181, w_035_598);
  nand2 I039_017(w_039_017, w_035_179, w_032_161);
  and2 I039_023(w_039_023, w_003_100, w_025_506);
  not1 I039_031(w_039_031, w_006_216);
  or2  I039_033(w_039_033, w_024_574, w_020_007);
  nand2 I039_036(w_039_036, w_029_193, w_004_010);
  not1 I039_037(w_039_037, w_020_128);
  and2 I039_040(w_039_040, w_026_091, w_018_158);
  nand2 I039_047(w_039_047, w_035_083, w_010_588);
  nand2 I039_049(w_039_049, w_004_009, w_027_796);
  not1 I039_051(w_039_051, w_020_071);
  nand2 I039_056(w_039_056, w_004_036, w_026_381);
  nand2 I039_057(w_039_057, w_033_709, w_027_445);
  not1 I039_062(w_039_062, w_031_043);
  not1 I039_066(w_039_066, w_004_014);
  or2  I039_067(w_039_067, w_002_350, w_008_494);
  and2 I039_074(w_039_074, w_013_421, w_037_074);
  not1 I039_089(w_039_089, w_010_717);
  not1 I039_096(w_039_096, w_033_691);
  or2  I039_103(w_039_103, w_026_068, w_031_004);
  or2  I039_116(w_039_116, w_016_416, w_019_002);
  and2 I039_119(w_039_119, w_030_028, w_026_061);
  or2  I039_122(w_039_122, w_014_482, w_014_013);
  not1 I039_125(w_039_125, w_036_066);
  nand2 I039_128(w_039_128, w_008_050, w_010_025);
  nand2 I039_129(w_039_129, w_013_370, w_023_154);
  or2  I039_136(w_039_136, w_031_030, w_000_968);
  and2 I039_144(w_039_144, w_024_486, w_020_114);
  and2 I039_145(w_039_145, w_013_327, w_010_192);
  not1 I039_146(w_039_146, w_007_419);
  not1 I039_149(w_039_149, w_007_463);
  nand2 I039_153(w_039_153, w_035_539, w_038_762);
  and2 I039_162(w_039_162, w_027_299, w_002_291);
  or2  I039_164(w_039_164, w_033_723, w_035_616);
  nand2 I039_170(w_039_170, w_005_082, w_021_039);
  or2  I039_175(w_039_175, w_017_024, w_017_026);
  nand2 I039_180(w_039_180, w_014_346, w_022_305);
  and2 I039_183(w_039_183, w_009_053, w_038_035);
  or2  I039_184(w_039_184, w_008_621, w_004_023);
  or2  I039_187(w_039_187, w_024_319, w_024_228);
  nand2 I039_188(w_039_188, w_028_049, w_035_326);
  and2 I039_189(w_039_189, w_016_448, w_027_145);
  and2 I039_190(w_039_190, w_015_532, w_029_103);
  or2  I039_197(w_039_197, w_004_021, w_021_033);
  nand2 I039_201(w_039_201, w_016_129, w_026_358);
  and2 I039_204(w_039_204, w_006_244, w_024_574);
  and2 I039_228(w_039_228, w_013_044, w_036_156);
  and2 I039_232(w_039_232, w_026_035, w_026_089);
  not1 I039_234(w_039_234, w_034_721);
  not1 I039_235(w_039_235, w_031_229);
  nand2 I039_243(w_039_243, w_000_982, w_026_356);
  and2 I039_250(w_039_250, w_021_348, w_024_012);
  nand2 I039_253(w_039_253, w_019_124, w_022_307);
  and2 I039_259(w_039_259, w_014_087, w_035_132);
  and2 I039_265(w_039_265, w_005_324, w_026_282);
  not1 I039_268(w_039_268, w_010_118);
  and2 I039_277(w_039_277, w_007_400, w_012_437);
  not1 I039_284(w_039_284, w_019_213);
  and2 I039_288(w_039_288, w_002_372, w_025_396);
  nand2 I039_289(w_039_289, w_013_387, w_007_281);
  or2  I039_299(w_039_299, w_005_016, w_038_447);
  and2 I039_303(w_039_303, w_002_246, w_009_026);
  or2  I039_305(w_039_305, w_030_044, w_010_367);
  and2 I039_309(w_039_309, w_026_399, w_009_000);
  nand2 I039_310(w_039_310, w_019_275, w_008_853);
  nand2 I039_312(w_039_312, w_013_148, w_028_146);
  and2 I039_332(w_039_332, w_024_104, w_031_442);
  or2  I039_333(w_039_333, w_025_286, w_032_499);
  or2  I039_336(w_039_336, w_030_050, w_032_298);
  or2  I039_340(w_039_340, w_020_030, w_029_139);
  or2  I039_349(w_039_349, w_022_113, w_018_048);
  nand2 I039_362(w_039_362, w_025_251, w_032_119);
  nand2 I039_371(w_039_371, w_017_020, w_016_037);
  or2  I039_375(w_039_375, w_037_040, w_017_001);
  not1 I039_377(w_039_377, w_031_211);
  or2  I039_381(w_039_381, w_019_101, w_036_273);
  not1 I039_382(w_039_382, w_024_285);
  or2  I039_385(w_039_385, w_030_347, w_006_225);
  or2  I039_392(w_039_392, w_005_076, w_026_051);
  nand2 I039_395(w_039_395, w_025_665, w_036_042);
  nand2 I039_400(w_039_400, w_001_678, w_038_114);
  and2 I039_405(w_039_405, w_015_264, w_009_059);
  not1 I039_413(w_039_413, w_037_111);
  or2  I039_417(w_039_417, w_003_019, w_007_222);
  nand2 I039_427(w_039_427, w_034_101, w_007_189);
  or2  I039_431(w_039_431, w_014_613, w_011_299);
  and2 I039_443(w_039_443, w_002_291, w_038_277);
  not1 I039_444(w_039_444, w_031_235);
  nand2 I039_450(w_039_450, w_024_388, w_003_168);
  or2  I039_456(w_039_456, w_026_047, w_029_187);
  not1 I039_459(w_039_459, w_033_031);
  not1 I039_460(w_039_460, w_023_212);
  and2 I039_461(w_039_461, w_038_012, w_004_033);
  not1 I040_003(w_040_003, w_013_198);
  or2  I040_008(w_040_008, w_015_128, w_007_318);
  and2 I040_016(w_040_016, w_011_175, w_006_140);
  and2 I040_017(w_040_017, w_035_160, w_004_030);
  or2  I040_025(w_040_025, w_020_062, w_025_187);
  not1 I040_026(w_040_026, w_032_144);
  and2 I040_027(w_040_027, w_003_136, w_012_257);
  nand2 I040_029(w_040_029, w_003_140, w_028_108);
  and2 I040_033(w_040_033, w_029_030, w_016_425);
  nand2 I040_037(w_040_037, w_028_862, w_002_446);
  nand2 I040_043(w_040_043, w_000_571, w_005_003);
  and2 I040_048(w_040_048, w_036_112, w_005_023);
  and2 I040_057(w_040_057, w_004_037, w_011_173);
  nand2 I040_058(w_040_058, w_016_124, w_031_019);
  nand2 I040_060(w_040_060, w_024_267, w_036_177);
  not1 I040_066(w_040_066, w_003_037);
  nand2 I040_068(w_040_068, w_014_159, w_031_297);
  or2  I040_071(w_040_071, w_003_155, w_007_238);
  not1 I040_075(w_040_075, w_019_322);
  not1 I040_083(w_040_083, w_025_468);
  or2  I040_084(w_040_084, w_008_131, w_005_174);
  not1 I040_089(w_040_089, w_008_225);
  not1 I040_095(w_040_095, w_039_184);
  nand2 I040_098(w_040_098, w_012_322, w_027_222);
  not1 I040_102(w_040_102, w_039_116);
  not1 I040_103(w_040_103, w_039_450);
  nand2 I040_104(w_040_104, w_025_041, w_036_084);
  nand2 I040_105(w_040_105, w_000_758, w_002_055);
  not1 I040_110(w_040_110, w_008_038);
  or2  I040_111(w_040_111, w_010_009, w_026_370);
  not1 I040_112(w_040_112, w_022_537);
  nand2 I040_113(w_040_113, w_020_091, w_010_008);
  not1 I040_115(w_040_115, w_032_336);
  nand2 I040_116(w_040_116, w_005_283, w_002_277);
  or2  I040_117(w_040_117, w_012_397, w_014_054);
  and2 I040_122(w_040_122, w_013_074, w_024_341);
  or2  I040_126(w_040_126, w_025_269, w_010_035);
  or2  I040_127(w_040_127, w_031_234, w_000_901);
  or2  I040_128(w_040_128, w_032_554, w_019_004);
  not1 I040_131(w_040_131, w_029_215);
  or2  I040_132(w_040_132, w_013_180, w_006_097);
  nand2 I040_140(w_040_140, w_021_082, w_002_457);
  and2 I040_141(w_040_141, w_037_154, w_015_652);
  or2  I040_142(w_040_142, w_020_133, w_038_665);
  not1 I040_148(w_040_148, w_011_122);
  or2  I040_149(w_040_149, w_015_004, w_014_518);
  and2 I040_151(w_040_151, w_013_453, w_035_152);
  and2 I040_152(w_040_152, w_002_092, w_025_480);
  nand2 I040_155(w_040_155, w_037_124, w_026_310);
  not1 I040_156(w_040_156, w_002_258);
  not1 I040_158(w_040_158, w_032_406);
  not1 I040_159(w_040_159, w_024_194);
  or2  I040_167(w_040_167, w_000_788, w_034_044);
  or2  I040_168(w_040_168, w_022_066, w_026_206);
  and2 I040_169(w_040_169, w_029_114, w_025_158);
  and2 I040_170(w_040_170, w_031_227, w_033_700);
  or2  I040_173(w_040_173, w_020_135, w_006_308);
  or2  I040_175(w_040_175, w_011_398, w_012_237);
  or2  I040_176(w_040_176, w_016_100, w_031_154);
  not1 I040_178(w_040_178, w_015_541);
  not1 I040_182(w_040_182, w_006_121);
  not1 I040_186(w_040_186, w_002_055);
  nand2 I040_194(w_040_194, w_004_013, w_015_636);
  nand2 I040_201(w_040_201, w_031_302, w_006_013);
  or2  I040_204(w_040_204, w_010_050, w_006_308);
  nand2 I040_207(w_040_207, w_010_134, w_007_390);
  and2 I040_210(w_040_210, w_021_076, w_007_234);
  nand2 I040_215(w_040_215, w_000_105, w_005_277);
  not1 I040_217(w_040_217, w_023_659);
  and2 I040_219(w_040_219, w_011_107, w_007_166);
  not1 I040_224(w_040_224, w_004_008);
  or2  I040_230(w_040_230, w_020_064, w_027_576);
  or2  I040_235(w_040_235, w_016_356, w_010_162);
  not1 I040_237(w_040_237, w_022_043);
  nand2 I040_243(w_040_243, w_005_055, w_019_015);
  or2  I040_245(w_040_245, w_030_358, w_020_014);
  not1 I040_248(w_040_248, w_032_655);
  nand2 I040_250(w_040_250, w_007_149, w_008_629);
  and2 I040_252(w_040_252, w_005_037, w_026_048);
  and2 I040_254(w_040_254, w_024_302, w_034_136);
  and2 I040_257(w_040_257, w_030_305, w_035_524);
  not1 I040_259(w_040_259, w_009_000);
  nand2 I040_264(w_040_264, w_000_481, w_014_125);
  nand2 I040_272(w_040_272, w_009_037, w_032_175);
  nand2 I040_274(w_040_274, w_002_152, w_022_428);
  nand2 I040_294(w_040_294, w_010_365, w_025_056);
  or2  I040_298(w_040_298, w_029_130, w_037_006);
  or2  I040_302(w_040_302, w_009_054, w_020_012);
  not1 I040_305(w_040_305, w_024_236);
  or2  I040_306(w_040_306, w_037_064, w_004_019);
  or2  I040_308(w_040_308, w_038_031, w_030_288);
  not1 I040_314(w_040_314, w_028_360);
  not1 I040_316(w_040_316, w_002_188);
  or2  I040_320(w_040_320, w_028_403, w_028_358);
  not1 I040_321(w_040_321, w_030_380);
  nand2 I040_322(w_040_322, w_022_426, w_002_414);
  nand2 I040_323(w_040_323, w_016_108, w_025_215);
  or2  I040_325(w_040_325, w_021_111, w_029_009);
  not1 I040_327(w_040_327, w_027_027);
  and2 I040_331(w_040_331, w_011_606, w_036_185);
  and2 I040_338(w_040_338, w_022_236, w_028_030);
  or2  I040_340(w_040_340, w_011_242, w_029_133);
  and2 I040_347(w_040_347, w_020_037, w_002_263);
  not1 I040_355(w_040_355, w_031_091);
  or2  I040_357(w_040_357, w_020_121, w_001_348);
  not1 I040_361(w_040_361, w_031_340);
  not1 I041_000(w_041_000, w_018_002);
  and2 I041_001(w_041_001, w_037_127, w_036_238);
  or2  I041_002(w_041_002, w_005_395, w_011_360);
  not1 I041_003(w_041_003, w_011_464);
  not1 I041_005(w_041_005, w_015_129);
  and2 I041_007(w_041_007, w_035_524, w_027_762);
  and2 I041_008(w_041_008, w_023_242, w_026_183);
  nand2 I041_009(w_041_009, w_034_596, w_018_120);
  not1 I041_010(w_041_010, w_032_380);
  or2  I041_011(w_041_011, w_040_323, w_031_312);
  or2  I041_012(w_041_012, w_007_044, w_023_037);
  not1 I041_014(w_041_014, w_019_084);
  and2 I041_015(w_041_015, w_026_419, w_004_007);
  not1 I041_016(w_041_016, w_020_045);
  not1 I041_017(w_041_017, w_014_582);
  not1 I041_018(w_041_018, w_017_000);
  nand2 I041_019(w_041_019, w_001_896, w_029_133);
  nand2 I041_020(w_041_020, w_011_030, w_028_012);
  not1 I041_022(w_041_022, w_021_039);
  and2 I041_023(w_041_023, w_001_004, w_000_609);
  or2  I041_026(w_041_026, w_008_174, w_019_241);
  or2  I041_027(w_041_027, w_030_231, w_012_338);
  and2 I041_028(w_041_028, w_026_097, w_010_006);
  nand2 I041_031(w_041_031, w_013_480, w_013_186);
  nand2 I041_032(w_041_032, w_019_042, w_001_549);
  not1 I041_033(w_041_033, w_020_013);
  and2 I041_035(w_041_035, w_014_540, w_023_664);
  and2 I041_036(w_041_036, w_017_002, w_025_005);
  or2  I041_037(w_041_037, w_011_486, w_026_407);
  and2 I041_039(w_041_039, w_015_618, w_022_183);
  and2 I041_043(w_041_043, w_036_113, w_007_080);
  not1 I041_044(w_041_044, w_007_218);
  not1 I041_045(w_041_045, w_020_019);
  and2 I041_047(w_041_047, w_034_001, w_033_435);
  and2 I041_048(w_041_048, w_019_329, w_019_060);
  and2 I041_049(w_041_049, w_010_140, w_020_134);
  nand2 I041_050(w_041_050, w_009_041, w_021_236);
  and2 I041_052(w_041_052, w_004_014, w_038_094);
  or2  I041_054(w_041_054, w_031_306, w_007_378);
  not1 I041_055(w_041_055, w_023_383);
  and2 I041_057(w_041_057, w_030_033, w_027_683);
  nand2 I041_058(w_041_058, w_011_262, w_015_221);
  nand2 I041_060(w_041_060, w_008_002, w_014_008);
  or2  I041_061(w_041_061, w_023_255, w_036_249);
  not1 I041_062(w_041_062, w_017_004);
  and2 I041_068(w_041_068, w_002_377, w_015_341);
  nand2 I041_070(w_041_070, w_001_211, w_008_446);
  or2  I041_071(w_041_071, w_024_364, w_028_237);
  nand2 I041_073(w_041_073, w_030_409, w_010_060);
  not1 I041_075(w_041_075, w_034_031);
  nand2 I041_076(w_041_076, w_023_277, w_038_748);
  and2 I041_077(w_041_077, w_007_194, w_014_128);
  not1 I041_078(w_041_078, w_001_005);
  and2 I041_079(w_041_079, w_040_207, w_023_197);
  or2  I041_082(w_041_082, w_023_622, w_039_400);
  or2  I041_083(w_041_083, w_024_491, w_028_647);
  nand2 I041_084(w_041_084, w_035_192, w_012_163);
  and2 I041_085(w_041_085, w_015_072, w_035_351);
  not1 I041_086(w_041_086, w_019_170);
  or2  I041_089(w_041_089, w_025_557, w_025_077);
  and2 I041_091(w_041_091, w_003_085, w_024_522);
  not1 I041_094(w_041_094, w_021_086);
  and2 I041_096(w_041_096, w_033_805, w_022_163);
  not1 I041_097(w_041_097, w_016_393);
  not1 I041_098(w_041_098, w_028_107);
  not1 I041_099(w_041_099, w_038_148);
  nand2 I041_100(w_041_100, w_021_075, w_036_008);
  nand2 I041_101(w_041_101, w_001_365, w_004_010);
  not1 I041_102(w_041_102, w_024_265);
  and2 I041_104(w_041_104, w_015_160, w_039_017);
  and2 I041_106(w_041_106, w_006_289, w_004_025);
  or2  I041_107(w_041_107, w_025_094, w_021_166);
  not1 I041_111(w_041_111, w_013_339);
  and2 I041_112(w_041_112, w_012_516, w_036_143);
  not1 I041_113(w_041_113, w_040_048);
  and2 I041_114(w_041_114, w_027_173, w_015_718);
  not1 I041_115(w_041_115, w_037_016);
  and2 I041_116(w_041_116, w_005_502, w_036_177);
  and2 I041_117(w_041_117, w_028_013, w_016_275);
  and2 I041_118(w_041_118, w_011_635, w_000_776);
  and2 I041_119(w_041_119, w_012_092, w_037_006);
  nand2 I041_120(w_041_120, w_039_067, w_034_099);
  or2  I041_121(w_041_121, w_008_169, w_034_160);
  not1 I041_122(w_041_122, w_017_019);
  or2  I042_001(w_042_001, w_015_018, w_010_200);
  not1 I042_002(w_042_002, w_024_056);
  nand2 I042_003(w_042_003, w_011_209, w_030_152);
  and2 I042_004(w_042_004, w_018_123, w_009_042);
  or2  I042_005(w_042_005, w_016_290, w_025_498);
  not1 I042_006(w_042_006, w_024_122);
  not1 I042_011(w_042_011, w_006_324);
  or2  I042_012(w_042_012, w_037_109, w_005_020);
  not1 I042_013(w_042_013, w_025_009);
  not1 I042_014(w_042_014, w_033_428);
  nand2 I042_016(w_042_016, w_005_352, w_036_247);
  nand2 I042_017(w_042_017, w_033_361, w_025_535);
  or2  I042_018(w_042_018, w_018_177, w_007_535);
  or2  I042_021(w_042_021, w_005_386, w_006_153);
  nand2 I042_024(w_042_024, w_017_024, w_024_267);
  nand2 I042_026(w_042_026, w_010_694, w_014_292);
  not1 I042_028(w_042_028, w_040_075);
  or2  I042_031(w_042_031, w_009_004, w_011_276);
  not1 I042_033(w_042_033, w_029_009);
  and2 I042_041(w_042_041, w_037_024, w_023_054);
  and2 I042_042(w_042_042, w_007_144, w_009_054);
  and2 I042_043(w_042_043, w_030_194, w_021_055);
  and2 I042_045(w_042_045, w_011_304, w_003_216);
  nand2 I042_046(w_042_046, w_030_275, w_010_518);
  nand2 I042_050(w_042_050, w_020_061, w_041_047);
  not1 I042_052(w_042_052, w_004_011);
  or2  I042_055(w_042_055, w_002_267, w_041_018);
  not1 I042_056(w_042_056, w_026_294);
  not1 I042_057(w_042_057, w_000_775);
  nand2 I042_059(w_042_059, w_023_178, w_007_192);
  nand2 I042_064(w_042_064, w_007_539, w_009_061);
  not1 I042_065(w_042_065, w_019_149);
  or2  I042_066(w_042_066, w_000_442, w_001_324);
  and2 I042_067(w_042_067, w_035_184, w_009_009);
  and2 I042_068(w_042_068, w_023_215, w_012_438);
  not1 I042_069(w_042_069, w_038_015);
  nand2 I042_070(w_042_070, w_041_071, w_022_236);
  nand2 I042_074(w_042_074, w_008_397, w_024_283);
  nand2 I042_077(w_042_077, w_003_151, w_039_201);
  not1 I042_078(w_042_078, w_025_203);
  and2 I042_081(w_042_081, w_023_127, w_030_342);
  or2  I042_083(w_042_083, w_029_135, w_030_186);
  and2 I042_084(w_042_084, w_028_235, w_002_471);
  nand2 I042_094(w_042_094, w_027_134, w_026_048);
  not1 I042_097(w_042_097, w_030_484);
  and2 I042_098(w_042_098, w_012_538, w_041_086);
  nand2 I042_099(w_042_099, w_016_038, w_037_043);
  nand2 I042_103(w_042_103, w_029_040, w_020_000);
  and2 I042_108(w_042_108, w_031_244, w_022_146);
  or2  I042_110(w_042_110, w_014_470, w_035_220);
  not1 I042_114(w_042_114, w_029_217);
  not1 I043_000(w_043_000, w_042_114);
  and2 I043_001(w_043_001, w_030_495, w_036_068);
  and2 I043_002(w_043_002, w_040_264, w_037_180);
  nand2 I043_003(w_043_003, w_021_352, w_025_144);
  and2 I043_004(w_043_004, w_007_509, w_012_396);
  not1 I043_005(w_043_005, w_039_253);
  not1 I043_006(w_043_006, w_026_088);
  and2 I043_007(w_043_007, w_008_490, w_020_032);
  and2 I043_009(w_043_009, w_007_078, w_016_363);
  nand2 I043_010(w_043_010, w_000_498, w_022_489);
  not1 I043_011(w_043_011, w_005_026);
  nand2 I043_013(w_043_013, w_019_064, w_025_295);
  and2 I043_014(w_043_014, w_026_374, w_020_115);
  not1 I043_015(w_043_015, w_019_043);
  not1 I043_016(w_043_016, w_027_681);
  not1 I043_017(w_043_017, w_014_137);
  not1 I043_018(w_043_018, w_000_119);
  nand2 I043_019(w_043_019, w_003_216, w_025_228);
  not1 I043_020(w_043_020, w_027_195);
  and2 I043_021(w_043_021, w_018_151, w_024_289);
  and2 I043_022(w_043_022, w_024_052, w_027_050);
  or2  I043_023(w_043_023, w_007_407, w_041_094);
  and2 I043_024(w_043_024, w_005_421, w_019_321);
  not1 I043_025(w_043_025, w_011_182);
  nand2 I043_027(w_043_027, w_027_344, w_008_568);
  and2 I043_028(w_043_028, w_027_118, w_016_142);
  not1 I043_029(w_043_029, w_040_066);
  or2  I043_031(w_043_031, w_020_064, w_000_853);
  nand2 I043_032(w_043_032, w_001_553, w_030_045);
  or2  I043_035(w_043_035, w_041_027, w_024_529);
  and2 I043_036(w_043_036, w_036_239, w_000_014);
  not1 I043_038(w_043_038, w_009_053);
  or2  I043_039(w_043_039, w_010_018, w_023_118);
  not1 I043_040(w_043_040, w_006_317);
  nand2 I043_041(w_043_041, w_004_004, w_016_161);
  or2  I043_042(w_043_042, w_006_201, w_016_349);
  nand2 I043_043(w_043_043, w_009_017, w_039_057);
  not1 I043_044(w_043_044, w_030_019);
  or2  I043_045(w_043_045, w_033_597, w_033_040);
  not1 I043_046(w_043_046, w_035_245);
  or2  I043_047(w_043_047, w_010_401, w_034_028);
  and2 I043_048(w_043_048, w_038_621, w_014_305);
  not1 I043_049(w_043_049, w_021_119);
  or2  I043_051(w_043_051, w_017_012, w_014_030);
  or2  I043_052(w_043_052, w_014_155, w_027_647);
  not1 I043_053(w_043_053, w_021_025);
  not1 I043_054(w_043_054, w_020_074);
  and2 I043_055(w_043_055, w_039_033, w_026_215);
  not1 I043_057(w_043_057, w_037_091);
  not1 I043_058(w_043_058, w_013_006);
  not1 I043_059(w_043_059, w_028_015);
  and2 I043_060(w_043_060, w_022_065, w_033_416);
  and2 I043_061(w_043_061, w_012_055, w_041_091);
  or2  I043_062(w_043_062, w_030_203, w_019_050);
  and2 I043_063(w_043_063, w_013_223, w_032_803);
  or2  I043_064(w_043_064, w_002_264, w_023_325);
  and2 I043_065(w_043_065, w_036_093, w_015_254);
  nand2 I044_007(w_044_007, w_031_094, w_013_276);
  not1 I044_012(w_044_012, w_040_089);
  nand2 I044_014(w_044_014, w_035_324, w_039_204);
  nand2 I044_015(w_044_015, w_020_016, w_019_335);
  nand2 I044_017(w_044_017, w_022_297, w_002_449);
  or2  I044_024(w_044_024, w_017_013, w_039_259);
  nand2 I044_031(w_044_031, w_033_301, w_010_430);
  and2 I044_033(w_044_033, w_017_015, w_024_051);
  nand2 I044_036(w_044_036, w_003_030, w_000_796);
  not1 I044_037(w_044_037, w_039_377);
  or2  I044_038(w_044_038, w_028_492, w_043_010);
  nand2 I044_039(w_044_039, w_001_033, w_002_397);
  nand2 I044_040(w_044_040, w_039_288, w_031_199);
  and2 I044_043(w_044_043, w_006_105, w_034_501);
  or2  I044_047(w_044_047, w_006_325, w_041_100);
  not1 I044_048(w_044_048, w_004_000);
  not1 I044_049(w_044_049, w_010_344);
  and2 I044_051(w_044_051, w_037_001, w_018_156);
  not1 I044_055(w_044_055, w_018_115);
  not1 I044_058(w_044_058, w_006_304);
  or2  I044_061(w_044_061, w_010_507, w_001_018);
  not1 I044_063(w_044_063, w_027_007);
  and2 I044_067(w_044_067, w_026_431, w_003_061);
  or2  I044_070(w_044_070, w_026_274, w_031_310);
  or2  I044_075(w_044_075, w_036_134, w_043_051);
  not1 I044_083(w_044_083, w_025_557);
  not1 I044_093(w_044_093, w_000_889);
  not1 I044_105(w_044_105, w_030_335);
  nand2 I044_107(w_044_107, w_014_348, w_023_578);
  and2 I044_110(w_044_110, w_001_147, w_019_121);
  not1 I044_114(w_044_114, w_043_006);
  nand2 I044_118(w_044_118, w_010_580, w_009_019);
  not1 I044_120(w_044_120, w_001_199);
  nand2 I044_128(w_044_128, w_015_083, w_030_248);
  not1 I044_133(w_044_133, w_001_769);
  or2  I044_139(w_044_139, w_040_186, w_006_169);
  or2  I044_140(w_044_140, w_007_063, w_012_303);
  not1 I044_142(w_044_142, w_020_072);
  or2  I044_145(w_044_145, w_039_349, w_026_269);
  not1 I044_155(w_044_155, w_041_098);
  nand2 I044_156(w_044_156, w_038_177, w_033_210);
  or2  I044_159(w_044_159, w_021_298, w_011_650);
  or2  I044_162(w_044_162, w_012_071, w_028_102);
  nand2 I044_166(w_044_166, w_006_145, w_042_052);
  or2  I044_172(w_044_172, w_028_762, w_017_026);
  and2 I044_174(w_044_174, w_027_236, w_005_124);
  not1 I044_175(w_044_175, w_019_371);
  not1 I044_181(w_044_181, w_040_357);
  and2 I044_183(w_044_183, w_025_516, w_032_121);
  and2 I044_184(w_044_184, w_035_127, w_035_245);
  and2 I044_188(w_044_188, w_023_153, w_016_112);
  and2 I044_193(w_044_193, w_038_180, w_028_625);
  and2 I044_194(w_044_194, w_020_072, w_015_759);
  and2 I044_198(w_044_198, w_043_031, w_001_743);
  not1 I044_199(w_044_199, w_011_604);
  or2  I044_203(w_044_203, w_014_560, w_017_006);
  nand2 I044_216(w_044_216, w_020_040, w_025_033);
  and2 I044_219(w_044_219, w_039_144, w_021_209);
  not1 I044_220(w_044_220, w_010_670);
  nand2 I044_223(w_044_223, w_016_381, w_020_015);
  and2 I044_227(w_044_227, w_036_073, w_034_270);
  or2  I044_231(w_044_231, w_020_130, w_019_157);
  not1 I044_232(w_044_232, w_021_029);
  not1 I044_234(w_044_234, w_004_035);
  and2 I044_261(w_044_261, w_037_051, w_014_485);
  not1 I044_263(w_044_263, w_022_193);
  or2  I044_273(w_044_273, w_031_368, w_003_102);
  nand2 I044_274(w_044_274, w_039_153, w_039_250);
  or2  I044_276(w_044_276, w_000_454, w_014_500);
  nand2 I044_278(w_044_278, w_021_053, w_041_043);
  nand2 I044_292(w_044_292, w_015_359, w_007_365);
  nand2 I044_296(w_044_296, w_015_443, w_025_039);
  nand2 I044_304(w_044_304, w_034_296, w_043_003);
  or2  I044_310(w_044_310, w_015_541, w_013_434);
  not1 I044_312(w_044_312, w_030_193);
  not1 I044_314(w_044_314, w_021_307);
  not1 I044_315(w_044_315, w_020_067);
  or2  I044_323(w_044_323, w_003_137, w_007_342);
  not1 I044_338(w_044_338, w_013_265);
  nand2 I044_341(w_044_341, w_004_026, w_041_016);
  nand2 I044_343(w_044_343, w_010_177, w_038_335);
  not1 I044_347(w_044_347, w_003_163);
  not1 I044_348(w_044_348, w_021_310);
  nand2 I044_356(w_044_356, w_040_152, w_035_051);
  not1 I044_360(w_044_360, w_003_071);
  or2  I044_365(w_044_365, w_009_008, w_038_764);
  not1 I044_371(w_044_371, w_000_956);
  and2 I044_378(w_044_378, w_001_140, w_028_470);
  or2  I044_384(w_044_384, w_024_539, w_005_238);
  not1 I044_386(w_044_386, w_043_027);
  and2 I044_391(w_044_391, w_028_318, w_022_081);
  not1 I044_392(w_044_392, w_038_238);
  nand2 I045_001(w_045_001, w_008_280, w_002_056);
  not1 I045_004(w_045_004, w_037_032);
  nand2 I045_005(w_045_005, w_008_803, w_017_022);
  nand2 I045_006(w_045_006, w_004_004, w_005_218);
  or2  I045_013(w_045_013, w_025_087, w_002_130);
  or2  I045_016(w_045_016, w_038_521, w_010_389);
  or2  I045_018(w_045_018, w_015_036, w_008_826);
  and2 I045_021(w_045_021, w_035_225, w_040_029);
  or2  I045_029(w_045_029, w_007_250, w_014_533);
  and2 I045_043(w_045_043, w_025_247, w_006_017);
  or2  I045_053(w_045_053, w_028_345, w_002_334);
  nand2 I045_067(w_045_067, w_043_019, w_015_465);
  not1 I045_074(w_045_074, w_033_511);
  not1 I045_076(w_045_076, w_000_520);
  or2  I045_079(w_045_079, w_025_132, w_036_082);
  nand2 I045_092(w_045_092, w_031_085, w_019_019);
  nand2 I045_093(w_045_093, w_028_065, w_033_041);
  and2 I045_102(w_045_102, w_017_012, w_034_483);
  nand2 I045_105(w_045_105, w_001_051, w_026_303);
  and2 I045_106(w_045_106, w_029_038, w_027_143);
  and2 I045_108(w_045_108, w_041_113, w_044_061);
  nand2 I045_110(w_045_110, w_014_322, w_036_066);
  and2 I045_111(w_045_111, w_015_211, w_031_196);
  and2 I045_123(w_045_123, w_014_401, w_012_299);
  nand2 I045_127(w_045_127, w_021_252, w_016_102);
  or2  I045_128(w_045_128, w_033_043, w_034_145);
  not1 I045_141(w_045_141, w_020_130);
  and2 I045_142(w_045_142, w_041_037, w_028_144);
  or2  I045_145(w_045_145, w_010_229, w_007_306);
  and2 I045_149(w_045_149, w_044_310, w_039_375);
  or2  I045_151(w_045_151, w_014_152, w_024_407);
  and2 I045_153(w_045_153, w_017_010, w_043_025);
  or2  I045_160(w_045_160, w_006_227, w_020_045);
  or2  I045_165(w_045_165, w_039_180, w_044_175);
  not1 I045_170(w_045_170, w_041_001);
  not1 I045_175(w_045_175, w_007_255);
  and2 I045_179(w_045_179, w_001_780, w_036_071);
  and2 I045_192(w_045_192, w_004_032, w_007_361);
  not1 I045_193(w_045_193, w_008_886);
  and2 I045_203(w_045_203, w_010_111, w_043_052);
  or2  I045_206(w_045_206, w_010_397, w_021_256);
  and2 I045_214(w_045_214, w_027_819, w_030_163);
  and2 I045_223(w_045_223, w_015_092, w_005_095);
  not1 I045_226(w_045_226, w_037_022);
  or2  I045_227(w_045_227, w_029_140, w_020_092);
  or2  I045_229(w_045_229, w_041_100, w_008_918);
  or2  I045_243(w_045_243, w_001_391, w_039_033);
  nand2 I045_252(w_045_252, w_033_196, w_004_036);
  or2  I045_253(w_045_253, w_003_123, w_000_239);
  not1 I045_255(w_045_255, w_018_051);
  not1 I045_258(w_045_258, w_024_072);
  not1 I045_271(w_045_271, w_037_116);
  and2 I045_277(w_045_277, w_026_309, w_027_625);
  nand2 I045_281(w_045_281, w_005_254, w_003_149);
  nand2 I045_294(w_045_294, w_006_328, w_039_136);
  nand2 I045_296(w_045_296, w_016_406, w_039_309);
  nand2 I045_315(w_045_315, w_005_373, w_039_277);
  nand2 I045_323(w_045_323, w_040_095, w_011_537);
  and2 I045_324(w_045_324, w_013_181, w_000_283);
  not1 I045_328(w_045_328, w_027_813);
  not1 I045_339(w_045_339, w_017_021);
  and2 I045_340(w_045_340, w_020_102, w_012_373);
  or2  I045_341(w_045_341, w_007_413, w_041_104);
  and2 I045_348(w_045_348, w_002_494, w_030_287);
  or2  I045_353(w_045_353, w_037_020, w_017_008);
  and2 I045_382(w_045_382, w_018_098, w_014_053);
  and2 I045_411(w_045_411, w_016_209, w_009_034);
  or2  I045_415(w_045_415, w_017_016, w_025_571);
  not1 I045_421(w_045_421, w_008_562);
  and2 I045_440(w_045_440, w_028_162, w_000_265);
  not1 I045_443(w_045_443, w_030_016);
  nand2 I045_467(w_045_467, w_040_305, w_008_392);
  nand2 I045_474(w_045_474, w_034_483, w_034_691);
  nand2 I045_500(w_045_500, w_008_488, w_030_004);
  or2  I045_503(w_045_503, w_010_448, w_025_238);
  not1 I045_505(w_045_505, w_002_129);
  and2 I045_506(w_045_506, w_011_456, w_030_049);
  or2  I045_511(w_045_511, w_000_025, w_013_239);
  and2 I045_531(w_045_531, w_033_856, w_034_684);
  not1 I045_534(w_045_534, w_037_004);
  not1 I045_548(w_045_548, w_034_725);
  not1 I045_549(w_045_549, w_011_101);
  and2 I045_560(w_045_560, w_022_398, w_042_042);
  not1 I045_563(w_045_563, w_000_223);
  not1 I045_564(w_045_564, w_043_019);
  nand2 I045_567(w_045_567, w_010_141, w_027_083);
  or2  I045_593(w_045_593, w_026_246, w_007_159);
  or2  I045_629(w_045_629, w_039_243, w_006_180);
  or2  I045_633(w_045_633, w_042_098, w_035_169);
  nand2 I045_662(w_045_662, w_021_035, w_023_242);
  not1 I045_667(w_045_667, w_032_322);
  and2 I045_692(w_045_692, w_013_316, w_024_136);
  or2  I046_000(w_046_000, w_018_084, w_016_381);
  nand2 I046_006(w_046_006, w_018_117, w_016_129);
  or2  I046_012(w_046_012, w_004_028, w_016_185);
  or2  I046_029(w_046_029, w_017_026, w_001_818);
  or2  I046_035(w_046_035, w_006_323, w_042_003);
  not1 I046_048(w_046_048, w_029_126);
  nand2 I046_052(w_046_052, w_015_172, w_020_044);
  not1 I046_059(w_046_059, w_021_307);
  and2 I046_062(w_046_062, w_027_300, w_019_111);
  nand2 I046_067(w_046_067, w_021_322, w_003_172);
  nand2 I046_070(w_046_070, w_004_013, w_011_050);
  or2  I046_076(w_046_076, w_035_114, w_034_054);
  not1 I046_091(w_046_091, w_022_322);
  or2  I046_097(w_046_097, w_004_021, w_032_098);
  not1 I046_098(w_046_098, w_002_144);
  or2  I046_115(w_046_115, w_045_294, w_012_252);
  not1 I046_120(w_046_120, w_011_017);
  and2 I046_122(w_046_122, w_004_007, w_006_119);
  or2  I046_141(w_046_141, w_024_183, w_045_500);
  and2 I046_143(w_046_143, w_004_027, w_024_217);
  and2 I046_148(w_046_148, w_040_025, w_023_134);
  not1 I046_156(w_046_156, w_015_744);
  not1 I046_157(w_046_157, w_008_226);
  and2 I046_158(w_046_158, w_013_442, w_028_088);
  or2  I046_171(w_046_171, w_005_078, w_018_184);
  nand2 I046_176(w_046_176, w_026_075, w_040_257);
  and2 I046_178(w_046_178, w_006_303, w_005_299);
  nand2 I046_179(w_046_179, w_002_000, w_028_323);
  and2 I046_181(w_046_181, w_006_091, w_016_367);
  or2  I046_182(w_046_182, w_002_123, w_024_588);
  and2 I046_184(w_046_184, w_015_216, w_006_034);
  or2  I046_185(w_046_185, w_011_245, w_026_435);
  not1 I046_194(w_046_194, w_030_314);
  or2  I046_195(w_046_195, w_032_113, w_012_088);
  and2 I046_212(w_046_212, w_026_326, w_033_902);
  not1 I046_294(w_046_294, w_007_437);
  not1 I046_300(w_046_300, w_028_768);
  nand2 I046_305(w_046_305, w_020_066, w_030_408);
  and2 I046_310(w_046_310, w_026_045, w_033_414);
  or2  I046_324(w_046_324, w_020_095, w_007_073);
  and2 I046_327(w_046_327, w_027_433, w_012_185);
  or2  I046_328(w_046_328, w_014_223, w_028_648);
  or2  I046_333(w_046_333, w_033_569, w_033_052);
  not1 I046_342(w_046_342, w_012_471);
  and2 I046_367(w_046_367, w_013_047, w_001_342);
  nand2 I046_386(w_046_386, w_045_281, w_012_248);
  and2 I046_393(w_046_393, w_015_095, w_017_007);
  not1 I046_414(w_046_414, w_025_199);
  and2 I046_420(w_046_420, w_014_080, w_007_070);
  not1 I046_421(w_046_421, w_026_387);
  nand2 I046_422(w_046_422, w_044_338, w_026_094);
  or2  I046_461(w_046_461, w_005_102, w_008_633);
  and2 I046_467(w_046_467, w_001_786, w_031_118);
  or2  I046_479(w_046_479, w_036_092, w_009_006);
  not1 I046_488(w_046_488, w_013_009);
  and2 I046_497(w_046_497, w_038_038, w_001_039);
  not1 I046_501(w_046_501, w_031_010);
  nand2 I046_504(w_046_504, w_030_490, w_018_129);
  nand2 I046_510(w_046_510, w_043_015, w_040_159);
  nand2 I046_525(w_046_525, w_042_006, w_045_411);
  not1 I046_539(w_046_539, w_041_079);
  not1 I046_540(w_046_540, w_040_158);
  nand2 I046_545(w_046_545, w_020_083, w_013_317);
  or2  I046_546(w_046_546, w_008_134, w_017_004);
  or2  I046_559(w_046_559, w_015_021, w_043_064);
  or2  I046_572(w_046_572, w_040_148, w_045_165);
  and2 I046_614(w_046_614, w_030_401, w_032_804);
  and2 I046_627(w_046_627, w_040_169, w_010_111);
  or2  I046_642(w_046_642, w_020_039, w_034_227);
  and2 I046_660(w_046_660, w_041_003, w_033_897);
  nand2 I046_664(w_046_664, w_003_174, w_013_274);
  nand2 I046_669(w_046_669, w_043_022, w_036_018);
  and2 I046_673(w_046_673, w_003_043, w_003_225);
  and2 I046_674(w_046_674, w_031_071, w_021_063);
  not1 I046_689(w_046_689, w_034_123);
  and2 I046_697(w_046_697, w_010_027, w_001_713);
  nand2 I046_733(w_046_733, w_033_145, w_013_228);
  not1 I046_734(w_046_734, w_009_047);
  nand2 I046_767(w_046_767, w_013_308, w_044_232);
  and2 I047_001(w_047_001, w_012_511, w_045_348);
  and2 I047_006(w_047_006, w_032_292, w_017_004);
  or2  I047_033(w_047_033, w_031_296, w_011_137);
  not1 I047_056(w_047_056, w_021_156);
  or2  I047_062(w_047_062, w_013_198, w_025_290);
  or2  I047_066(w_047_066, w_046_504, w_035_089);
  not1 I047_067(w_047_067, w_002_388);
  or2  I047_082(w_047_082, w_003_092, w_002_369);
  nand2 I047_095(w_047_095, w_002_462, w_001_059);
  not1 I047_096(w_047_096, w_022_072);
  not1 I047_098(w_047_098, w_024_344);
  and2 I047_105(w_047_105, w_030_318, w_017_019);
  and2 I047_107(w_047_107, w_019_073, w_010_531);
  or2  I047_118(w_047_118, w_016_252, w_012_110);
  or2  I047_124(w_047_124, w_030_362, w_025_107);
  and2 I047_146(w_047_146, w_025_660, w_013_389);
  and2 I047_157(w_047_157, w_028_574, w_015_778);
  and2 I047_158(w_047_158, w_021_270, w_044_234);
  and2 I047_164(w_047_164, w_031_241, w_041_076);
  not1 I047_171(w_047_171, w_040_037);
  and2 I047_176(w_047_176, w_015_134, w_003_171);
  not1 I047_178(w_047_178, w_037_041);
  and2 I047_183(w_047_183, w_021_143, w_030_258);
  nand2 I047_187(w_047_187, w_017_022, w_043_000);
  or2  I047_188(w_047_188, w_000_721, w_046_115);
  and2 I047_190(w_047_190, w_000_804, w_029_071);
  not1 I047_203(w_047_203, w_010_452);
  nand2 I047_208(w_047_208, w_012_332, w_024_218);
  or2  I047_212(w_047_212, w_033_042, w_036_016);
  and2 I047_226(w_047_226, w_014_629, w_039_056);
  or2  I047_229(w_047_229, w_020_000, w_012_161);
  and2 I047_230(w_047_230, w_017_010, w_041_005);
  nand2 I047_232(w_047_232, w_009_047, w_027_668);
  and2 I047_238(w_047_238, w_032_591, w_008_815);
  not1 I047_244(w_047_244, w_001_199);
  and2 I047_245(w_047_245, w_003_042, w_039_125);
  and2 I047_247(w_047_247, w_016_404, w_044_347);
  or2  I047_257(w_047_257, w_040_060, w_022_282);
  or2  I047_262(w_047_262, w_011_044, w_014_128);
  nand2 I047_272(w_047_272, w_035_540, w_020_068);
  or2  I047_278(w_047_278, w_030_109, w_009_008);
  or2  I047_279(w_047_279, w_044_049, w_015_093);
  nand2 I047_281(w_047_281, w_007_507, w_044_017);
  or2  I047_288(w_047_288, w_004_035, w_010_628);
  nand2 I047_289(w_047_289, w_025_188, w_039_145);
  or2  I047_295(w_047_295, w_016_006, w_022_090);
  and2 I047_327(w_047_327, w_009_059, w_007_068);
  nand2 I047_332(w_047_332, w_015_164, w_009_052);
  or2  I047_339(w_047_339, w_046_510, w_039_031);
  or2  I047_348(w_047_348, w_028_013, w_033_849);
  and2 I047_357(w_047_357, w_019_345, w_022_376);
  or2  I047_364(w_047_364, w_013_335, w_009_012);
  or2  I047_379(w_047_379, w_010_715, w_033_493);
  nand2 I047_385(w_047_385, w_012_262, w_032_332);
  or2  I047_386(w_047_386, w_044_033, w_044_193);
  nand2 I047_396(w_047_396, w_042_103, w_007_401);
  or2  I047_401(w_047_401, w_044_360, w_011_156);
  or2  I047_404(w_047_404, w_009_032, w_020_075);
  and2 I047_427(w_047_427, w_003_097, w_003_083);
  nand2 I047_436(w_047_436, w_014_070, w_017_008);
  not1 I047_443(w_047_443, w_009_064);
  nand2 I047_448(w_047_448, w_007_200, w_018_124);
  nand2 I047_450(w_047_450, w_022_416, w_014_025);
  or2  I047_460(w_047_460, w_020_103, w_046_386);
  not1 I047_464(w_047_464, w_034_805);
  or2  I047_470(w_047_470, w_005_401, w_024_377);
  or2  I047_472(w_047_472, w_032_715, w_020_037);
  nand2 I047_474(w_047_474, w_026_124, w_040_250);
  nand2 I047_475(w_047_475, w_038_621, w_020_020);
  and2 I047_481(w_047_481, w_025_317, w_043_065);
  and2 I047_485(w_047_485, w_019_255, w_013_365);
  or2  I047_492(w_047_492, w_045_315, w_015_175);
  not1 I048_018(w_048_018, w_032_753);
  nand2 I048_023(w_048_023, w_004_002, w_039_312);
  not1 I048_029(w_048_029, w_010_506);
  nand2 I048_034(w_048_034, w_017_022, w_031_078);
  or2  I048_050(w_048_050, w_009_020, w_011_010);
  not1 I048_068(w_048_068, w_023_333);
  and2 I048_070(w_048_070, w_038_713, w_011_578);
  not1 I048_078(w_048_078, w_000_670);
  and2 I048_089(w_048_089, w_035_629, w_015_072);
  or2  I048_090(w_048_090, w_024_042, w_041_085);
  or2  I048_095(w_048_095, w_005_493, w_041_070);
  or2  I048_097(w_048_097, w_013_465, w_038_041);
  nand2 I048_101(w_048_101, w_044_348, w_028_186);
  nand2 I048_111(w_048_111, w_023_100, w_025_405);
  nand2 I048_114(w_048_114, w_043_019, w_002_199);
  and2 I048_116(w_048_116, w_042_097, w_000_752);
  not1 I048_118(w_048_118, w_046_012);
  nand2 I048_121(w_048_121, w_034_149, w_033_601);
  not1 I048_133(w_048_133, w_003_216);
  and2 I048_136(w_048_136, w_015_036, w_008_053);
  and2 I048_139(w_048_139, w_002_032, w_037_081);
  or2  I048_158(w_048_158, w_008_022, w_046_414);
  or2  I048_161(w_048_161, w_046_141, w_026_063);
  not1 I048_188(w_048_188, w_032_716);
  nand2 I048_189(w_048_189, w_010_114, w_043_016);
  nand2 I048_198(w_048_198, w_028_876, w_036_262);
  nand2 I048_201(w_048_201, w_024_142, w_040_113);
  or2  I048_203(w_048_203, w_014_375, w_014_033);
  not1 I048_205(w_048_205, w_011_412);
  not1 I048_218(w_048_218, w_012_382);
  and2 I048_227(w_048_227, w_030_198, w_041_015);
  nand2 I048_276(w_048_276, w_037_119, w_032_315);
  and2 I048_285(w_048_285, w_021_127, w_023_445);
  nand2 I048_296(w_048_296, w_010_267, w_022_278);
  and2 I048_308(w_048_308, w_002_307, w_017_026);
  not1 I048_313(w_048_313, w_008_377);
  nand2 I048_320(w_048_320, w_014_109, w_020_124);
  and2 I048_335(w_048_335, w_004_017, w_012_392);
  and2 I048_348(w_048_348, w_011_130, w_001_763);
  and2 I048_368(w_048_368, w_041_022, w_016_124);
  or2  I048_380(w_048_380, w_028_648, w_012_114);
  nand2 I048_384(w_048_384, w_005_165, w_047_289);
  and2 I048_385(w_048_385, w_001_734, w_022_258);
  or2  I048_410(w_048_410, w_018_144, w_032_020);
  not1 I048_412(w_048_412, w_026_321);
  or2  I048_418(w_048_418, w_013_244, w_023_405);
  not1 I048_427(w_048_427, w_008_466);
  not1 I048_445(w_048_445, w_014_383);
  or2  I048_448(w_048_448, w_006_191, w_013_152);
  not1 I048_450(w_048_450, w_010_156);
  and2 I048_458(w_048_458, w_017_001, w_018_117);
  not1 I048_479(w_048_479, w_000_018);
  not1 I048_490(w_048_490, w_031_025);
  or2  I048_493(w_048_493, w_019_197, w_042_108);
  not1 I048_517(w_048_517, w_022_383);
  nand2 I048_519(w_048_519, w_037_070, w_012_177);
  nand2 I048_525(w_048_525, w_030_282, w_042_011);
  not1 I048_542(w_048_542, w_032_370);
  not1 I048_552(w_048_552, w_046_098);
  not1 I048_559(w_048_559, w_015_547);
  not1 I048_575(w_048_575, w_012_416);
  or2  I048_591(w_048_591, w_040_131, w_030_244);
  nand2 I048_595(w_048_595, w_006_009, w_009_034);
  not1 I048_599(w_048_599, w_009_041);
  not1 I048_605(w_048_605, w_036_052);
  and2 I048_606(w_048_606, w_013_020, w_001_551);
  nand2 I048_620(w_048_620, w_012_061, w_013_324);
  nand2 I048_673(w_048_673, w_022_527, w_010_107);
  or2  I048_679(w_048_679, w_045_503, w_008_435);
  and2 I048_694(w_048_694, w_040_104, w_025_488);
  nand2 I048_706(w_048_706, w_047_229, w_001_353);
  nand2 I048_732(w_048_732, w_027_108, w_002_496);
  and2 I048_734(w_048_734, w_030_123, w_038_101);
  nand2 I048_738(w_048_738, w_038_188, w_005_264);
  not1 I048_748(w_048_748, w_030_151);
  nand2 I048_780(w_048_780, w_034_618, w_032_778);
  or2  I048_801(w_048_801, w_037_061, w_030_415);
  and2 I048_803(w_048_803, w_018_109, w_037_105);
  not1 I048_816(w_048_816, w_014_516);
  nand2 I049_003(w_049_003, w_017_017, w_035_592);
  and2 I049_018(w_049_018, w_008_822, w_015_235);
  not1 I049_041(w_049_041, w_017_009);
  or2  I049_044(w_049_044, w_012_263, w_001_523);
  or2  I049_069(w_049_069, w_018_182, w_003_015);
  or2  I049_071(w_049_071, w_028_527, w_021_091);
  not1 I049_075(w_049_075, w_034_334);
  nand2 I049_078(w_049_078, w_000_728, w_047_492);
  not1 I049_147(w_049_147, w_029_202);
  or2  I049_190(w_049_190, w_036_040, w_032_692);
  or2  I049_192(w_049_192, w_048_133, w_036_085);
  nand2 I049_194(w_049_194, w_048_410, w_026_056);
  nand2 I049_210(w_049_210, w_040_215, w_001_514);
  nand2 I049_217(w_049_217, w_024_138, w_007_348);
  and2 I049_218(w_049_218, w_029_042, w_010_817);
  and2 I049_220(w_049_220, w_024_183, w_022_256);
  nand2 I049_245(w_049_245, w_007_399, w_014_057);
  or2  I049_246(w_049_246, w_034_693, w_016_376);
  and2 I049_247(w_049_247, w_037_076, w_038_206);
  and2 I049_250(w_049_250, w_013_382, w_044_107);
  nand2 I049_259(w_049_259, w_043_009, w_005_289);
  and2 I049_270(w_049_270, w_040_175, w_015_782);
  not1 I049_298(w_049_298, w_030_145);
  and2 I049_307(w_049_307, w_035_081, w_046_070);
  and2 I049_309(w_049_309, w_038_612, w_004_006);
  nand2 I049_321(w_049_321, w_015_027, w_020_126);
  not1 I049_327(w_049_327, w_006_237);
  nand2 I049_329(w_049_329, w_035_054, w_046_212);
  and2 I049_334(w_049_334, w_039_164, w_010_501);
  nand2 I049_338(w_049_338, w_003_222, w_011_129);
  or2  I049_341(w_049_341, w_024_166, w_029_120);
  nand2 I049_343(w_049_343, w_045_110, w_001_247);
  not1 I049_358(w_049_358, w_046_488);
  not1 I049_363(w_049_363, w_015_159);
  or2  I049_383(w_049_383, w_022_097, w_040_235);
  not1 I049_397(w_049_397, w_001_324);
  or2  I049_412(w_049_412, w_022_543, w_001_701);
  or2  I049_414(w_049_414, w_004_032, w_011_263);
  nand2 I049_445(w_049_445, w_037_013, w_032_668);
  and2 I049_454(w_049_454, w_029_038, w_026_317);
  nand2 I049_459(w_049_459, w_026_001, w_034_096);
  not1 I049_470(w_049_470, w_006_050);
  or2  I049_478(w_049_478, w_016_218, w_009_061);
  not1 I049_516(w_049_516, w_039_122);
  nand2 I049_521(w_049_521, w_024_084, w_020_057);
  and2 I049_525(w_049_525, w_013_129, w_000_851);
  or2  I049_534(w_049_534, w_022_360, w_041_119);
  and2 I049_541(w_049_541, w_042_024, w_026_217);
  and2 I049_548(w_049_548, w_025_250, w_023_553);
  nand2 I049_587(w_049_587, w_040_224, w_040_060);
  or2  I049_602(w_049_602, w_027_546, w_046_310);
  and2 I049_607(w_049_607, w_002_226, w_032_654);
  and2 I049_619(w_049_619, w_029_183, w_048_116);
  nand2 I049_623(w_049_623, w_029_047, w_031_308);
  nand2 I049_629(w_049_629, w_001_360, w_019_191);
  or2  I049_633(w_049_633, w_028_397, w_024_145);
  or2  I049_649(w_049_649, w_030_053, w_037_097);
  not1 I049_651(w_049_651, w_026_039);
  not1 I049_654(w_049_654, w_008_218);
  or2  I049_657(w_049_657, w_002_356, w_038_235);
  or2  I049_690(w_049_690, w_028_349, w_000_574);
  not1 I049_691(w_049_691, w_043_043);
  not1 I049_706(w_049_706, w_040_325);
  or2  I049_739(w_049_739, w_009_021, w_028_546);
  not1 I049_742(w_049_742, w_017_027);
  and2 I049_750(w_049_750, w_044_024, w_028_366);
  not1 I049_786(w_049_786, w_019_064);
  nand2 I049_797(w_049_797, w_006_082, w_045_440);
  or2  I049_828(w_049_828, w_026_436, w_013_418);
  nand2 I049_835(w_049_835, w_041_091, w_040_033);
  nand2 I049_855(w_049_855, w_019_269, w_022_205);
  or2  I049_879(w_049_879, w_018_093, w_040_152);
  nand2 I049_883(w_049_883, w_042_094, w_046_048);
  not1 I049_886(w_049_886, w_034_076);
  or2  I049_913(w_049_913, w_040_327, w_039_013);
  nand2 I049_925(w_049_925, w_037_165, w_020_106);
  and2 I049_930(w_049_930, w_014_554, w_010_716);
  nand2 I049_936(w_049_936, w_026_328, w_023_020);
  not1 I049_943(w_049_943, w_016_228);
  or2  I049_944(w_049_944, w_009_022, w_015_210);
  and2 I049_965(w_049_965, w_015_118, w_041_052);
  or2  I050_002(w_050_002, w_040_252, w_045_382);
  not1 I050_003(w_050_003, w_042_066);
  or2  I050_005(w_050_005, w_026_106, w_029_154);
  nand2 I050_035(w_050_035, w_048_188, w_026_340);
  or2  I050_037(w_050_037, w_002_193, w_004_016);
  not1 I050_038(w_050_038, w_013_362);
  or2  I050_039(w_050_039, w_041_028, w_012_409);
  and2 I050_044(w_050_044, w_034_235, w_009_034);
  or2  I050_058(w_050_058, w_002_245, w_010_573);
  not1 I050_059(w_050_059, w_034_555);
  not1 I050_068(w_050_068, w_030_242);
  or2  I050_083(w_050_083, w_043_046, w_021_320);
  or2  I050_086(w_050_086, w_038_149, w_036_138);
  and2 I050_088(w_050_088, w_036_115, w_033_247);
  or2  I050_100(w_050_100, w_033_267, w_028_482);
  nand2 I050_102(w_050_102, w_015_131, w_044_067);
  nand2 I050_111(w_050_111, w_020_012, w_023_184);
  not1 I050_141(w_050_141, w_001_091);
  not1 I050_147(w_050_147, w_045_506);
  nand2 I050_152(w_050_152, w_033_778, w_035_382);
  or2  I050_159(w_050_159, w_003_140, w_013_297);
  or2  I050_166(w_050_166, w_046_143, w_046_664);
  or2  I050_186(w_050_186, w_045_341, w_000_850);
  nand2 I050_192(w_050_192, w_039_189, w_016_354);
  or2  I050_195(w_050_195, w_022_455, w_028_066);
  or2  I050_198(w_050_198, w_048_385, w_002_188);
  or2  I050_200(w_050_200, w_048_599, w_014_270);
  and2 I050_215(w_050_215, w_028_496, w_044_145);
  nand2 I050_229(w_050_229, w_001_780, w_035_120);
  nand2 I050_231(w_050_231, w_046_305, w_014_147);
  or2  I050_237(w_050_237, w_015_187, w_017_027);
  nand2 I050_244(w_050_244, w_026_158, w_040_115);
  or2  I050_247(w_050_247, w_039_066, w_045_175);
  and2 I050_248(w_050_248, w_023_530, w_034_044);
  not1 I050_250(w_050_250, w_014_289);
  and2 I050_255(w_050_255, w_012_265, w_010_756);
  nand2 I050_264(w_050_264, w_030_367, w_017_025);
  nand2 I050_282(w_050_282, w_000_637, w_023_459);
  nand2 I050_289(w_050_289, w_016_465, w_022_088);
  nand2 I050_294(w_050_294, w_029_117, w_022_429);
  not1 I050_299(w_050_299, w_032_225);
  nand2 I050_301(w_050_301, w_043_040, w_017_018);
  and2 I050_311(w_050_311, w_014_031, w_047_485);
  and2 I050_322(w_050_322, w_041_012, w_003_159);
  or2  I050_323(w_050_323, w_028_062, w_045_127);
  nand2 I050_344(w_050_344, w_026_323, w_018_067);
  and2 I050_353(w_050_353, w_019_279, w_044_219);
  nand2 I050_361(w_050_361, w_003_180, w_014_320);
  and2 I050_365(w_050_365, w_035_142, w_037_005);
  or2  I050_366(w_050_366, w_009_044, w_027_776);
  not1 I050_369(w_050_369, w_014_218);
  not1 I050_370(w_050_370, w_030_002);
  or2  I050_371(w_050_371, w_014_291, w_026_408);
  not1 I050_376(w_050_376, w_005_056);
  or2  I050_386(w_050_386, w_033_723, w_040_306);
  and2 I050_389(w_050_389, w_008_161, w_032_212);
  not1 I050_395(w_050_395, w_045_252);
  not1 I050_396(w_050_396, w_013_479);
  not1 I050_401(w_050_401, w_035_145);
  and2 I050_407(w_050_407, w_022_243, w_011_394);
  nand2 I050_409(w_050_409, w_013_241, w_012_387);
  or2  I050_413(w_050_413, w_041_033, w_019_291);
  not1 I050_423(w_050_423, w_016_208);
  not1 I050_438(w_050_438, w_016_207);
  not1 I050_469(w_050_469, w_040_151);
  nand2 I051_002(w_051_002, w_015_395, w_033_067);
  or2  I051_023(w_051_023, w_009_030, w_026_098);
  and2 I051_031(w_051_031, w_004_009, w_007_299);
  and2 I051_037(w_051_037, w_019_342, w_022_002);
  and2 I051_046(w_051_046, w_006_063, w_030_420);
  nand2 I051_047(w_051_047, w_025_542, w_000_965);
  not1 I051_050(w_051_050, w_027_006);
  and2 I051_060(w_051_060, w_027_041, w_023_015);
  or2  I051_066(w_051_066, w_035_078, w_030_423);
  or2  I051_069(w_051_069, w_004_029, w_045_340);
  nand2 I051_071(w_051_071, w_000_813, w_007_042);
  nand2 I051_075(w_051_075, w_029_064, w_038_194);
  and2 I051_094(w_051_094, w_023_666, w_037_103);
  not1 I051_102(w_051_102, w_001_072);
  nand2 I051_108(w_051_108, w_006_009, w_026_054);
  nand2 I051_114(w_051_114, w_026_361, w_018_025);
  nand2 I051_115(w_051_115, w_019_138, w_003_125);
  nand2 I051_118(w_051_118, w_043_001, w_010_232);
  nand2 I051_123(w_051_123, w_045_564, w_031_413);
  or2  I051_129(w_051_129, w_035_487, w_013_228);
  and2 I051_134(w_051_134, w_021_259, w_000_963);
  not1 I051_138(w_051_138, w_013_028);
  not1 I051_142(w_051_142, w_032_187);
  not1 I051_161(w_051_161, w_044_133);
  not1 I051_165(w_051_165, w_018_064);
  or2  I051_167(w_051_167, w_047_188, w_022_388);
  and2 I051_178(w_051_178, w_034_242, w_020_128);
  nand2 I051_179(w_051_179, w_034_115, w_019_191);
  and2 I051_184(w_051_184, w_046_767, w_043_063);
  and2 I051_196(w_051_196, w_042_108, w_024_590);
  not1 I051_204(w_051_204, w_049_217);
  or2  I051_223(w_051_223, w_003_132, w_043_052);
  or2  I051_240(w_051_240, w_017_000, w_025_206);
  not1 I051_249(w_051_249, w_034_164);
  not1 I051_255(w_051_255, w_010_734);
  nand2 I051_286(w_051_286, w_018_092, w_018_038);
  or2  I051_288(w_051_288, w_035_415, w_013_064);
  not1 I051_290(w_051_290, w_027_124);
  not1 I051_299(w_051_299, w_033_834);
  not1 I051_306(w_051_306, w_009_011);
  nand2 I051_307(w_051_307, w_035_032, w_036_175);
  and2 I051_308(w_051_308, w_043_020, w_010_012);
  nand2 I051_313(w_051_313, w_022_291, w_041_049);
  nand2 I051_314(w_051_314, w_045_193, w_004_023);
  and2 I051_317(w_051_317, w_041_073, w_037_152);
  not1 I051_318(w_051_318, w_020_083);
  or2  I051_320(w_051_320, w_026_025, w_038_543);
  nand2 I051_327(w_051_327, w_041_035, w_004_014);
  or2  I051_336(w_051_336, w_005_173, w_004_020);
  nand2 I051_339(w_051_339, w_037_063, w_009_005);
  and2 I051_342(w_051_342, w_002_218, w_033_038);
  not1 I051_356(w_051_356, w_022_319);
  and2 I051_360(w_051_360, w_014_282, w_028_052);
  or2  I051_370(w_051_370, w_037_176, w_021_039);
  not1 I051_372(w_051_372, w_025_208);
  and2 I051_381(w_051_381, w_011_226, w_044_296);
  nand2 I051_382(w_051_382, w_016_390, w_033_402);
  nand2 I051_384(w_051_384, w_037_014, w_012_124);
  or2  I051_392(w_051_392, w_031_004, w_010_053);
  not1 I051_404(w_051_404, w_037_183);
  or2  I051_409(w_051_409, w_037_113, w_033_571);
  or2  I051_413(w_051_413, w_029_036, w_010_010);
  nand2 I051_417(w_051_417, w_015_098, w_048_089);
  and2 I051_420(w_051_420, w_011_200, w_014_380);
  and2 I051_438(w_051_438, w_011_505, w_023_614);
  and2 I051_439(w_051_439, w_014_095, w_021_065);
  and2 I051_457(w_051_457, w_007_427, w_049_041);
  not1 I051_517(w_051_517, w_046_697);
  not1 I051_527(w_051_527, w_030_052);
  not1 I051_540(w_051_540, w_006_287);
  nand2 I052_002(w_052_002, w_036_023, w_030_158);
  not1 I052_004(w_052_004, w_046_076);
  not1 I052_006(w_052_006, w_009_004);
  or2  I052_007(w_052_007, w_020_020, w_019_332);
  nand2 I052_008(w_052_008, w_016_422, w_011_523);
  nand2 I052_009(w_052_009, w_023_206, w_033_406);
  not1 I052_012(w_052_012, w_046_029);
  and2 I052_013(w_052_013, w_031_050, w_018_101);
  not1 I052_015(w_052_015, w_028_276);
  or2  I052_016(w_052_016, w_027_526, w_046_097);
  nand2 I052_017(w_052_017, w_043_062, w_026_228);
  and2 I052_022(w_052_022, w_034_429, w_026_421);
  and2 I052_023(w_052_023, w_048_519, w_035_024);
  not1 I052_026(w_052_026, w_009_048);
  or2  I052_029(w_052_029, w_033_763, w_023_015);
  or2  I052_030(w_052_030, w_009_015, w_025_656);
  not1 I052_031(w_052_031, w_041_078);
  and2 I052_034(w_052_034, w_051_179, w_041_008);
  nand2 I052_035(w_052_035, w_050_044, w_032_151);
  or2  I052_036(w_052_036, w_032_210, w_034_045);
  or2  I052_037(w_052_037, w_035_051, w_032_649);
  and2 I052_041(w_052_041, w_010_040, w_010_543);
  or2  I052_046(w_052_046, w_018_125, w_017_001);
  nand2 I052_049(w_052_049, w_014_446, w_008_319);
  nand2 I052_051(w_052_051, w_026_298, w_035_145);
  and2 I052_053(w_052_053, w_018_052, w_001_435);
  not1 I052_058(w_052_058, w_034_446);
  not1 I052_059(w_052_059, w_051_223);
  not1 I052_060(w_052_060, w_010_804);
  and2 I052_062(w_052_062, w_023_110, w_029_174);
  not1 I052_064(w_052_064, w_034_317);
  or2  I052_067(w_052_067, w_019_093, w_019_297);
  and2 I052_068(w_052_068, w_025_640, w_028_112);
  nand2 I052_071(w_052_071, w_012_525, w_024_437);
  or2  I052_073(w_052_073, w_008_209, w_008_959);
  nand2 I052_078(w_052_078, w_000_455, w_028_462);
  and2 I052_080(w_052_080, w_004_014, w_029_106);
  nand2 I052_082(w_052_082, w_035_633, w_011_655);
  nand2 I052_099(w_052_099, w_020_081, w_040_294);
  not1 I052_100(w_052_100, w_049_220);
  or2  I052_101(w_052_101, w_026_264, w_051_413);
  and2 I052_102(w_052_102, w_009_044, w_023_503);
  and2 I052_106(w_052_106, w_028_854, w_031_121);
  and2 I052_108(w_052_108, w_027_717, w_024_000);
  and2 I052_109(w_052_109, w_023_099, w_014_344);
  nand2 I052_115(w_052_115, w_006_173, w_019_255);
  nand2 I052_117(w_052_117, w_009_040, w_024_122);
  nand2 I052_120(w_052_120, w_008_126, w_001_226);
  nand2 I052_121(w_052_121, w_004_024, w_000_767);
  nand2 I052_125(w_052_125, w_027_171, w_000_106);
  nand2 I052_126(w_052_126, w_023_558, w_001_488);
  nand2 I052_128(w_052_128, w_010_738, w_008_217);
  and2 I052_129(w_052_129, w_020_114, w_051_050);
  or2  I052_132(w_052_132, w_002_208, w_044_220);
  not1 I052_133(w_052_133, w_000_272);
  not1 I052_135(w_052_135, w_019_248);
  nand2 I052_137(w_052_137, w_049_548, w_001_260);
  not1 I052_143(w_052_143, w_038_202);
  not1 I052_144(w_052_144, w_016_079);
  nand2 I052_145(w_052_145, w_030_073, w_032_232);
  and2 I052_147(w_052_147, w_003_072, w_000_527);
  or2  I052_148(w_052_148, w_008_182, w_033_905);
  or2  I052_150(w_052_150, w_029_148, w_007_377);
  nand2 I052_152(w_052_152, w_016_142, w_032_449);
  and2 I052_153(w_052_153, w_021_335, w_038_009);
  not1 I052_160(w_052_160, w_024_401);
  and2 I052_162(w_052_162, w_038_277, w_014_248);
  or2  I052_164(w_052_164, w_029_089, w_018_157);
  and2 I052_165(w_052_165, w_014_577, w_043_036);
  not1 I053_002(w_053_002, w_006_007);
  nand2 I053_005(w_053_005, w_048_445, w_003_035);
  and2 I053_012(w_053_012, w_026_332, w_024_024);
  nand2 I053_019(w_053_019, w_052_162, w_023_051);
  or2  I053_022(w_053_022, w_052_165, w_021_059);
  nand2 I053_030(w_053_030, w_029_173, w_048_450);
  and2 I053_036(w_053_036, w_001_070, w_028_211);
  not1 I053_042(w_053_042, w_005_395);
  nand2 I053_053(w_053_053, w_020_046, w_025_519);
  or2  I053_055(w_053_055, w_051_370, w_005_002);
  and2 I053_058(w_053_058, w_051_320, w_027_227);
  not1 I053_069(w_053_069, w_024_082);
  or2  I053_070(w_053_070, w_016_195, w_003_160);
  not1 I053_081(w_053_081, w_048_205);
  or2  I053_089(w_053_089, w_048_285, w_031_332);
  nand2 I053_092(w_053_092, w_009_010, w_052_059);
  and2 I053_102(w_053_102, w_028_511, w_015_106);
  or2  I053_109(w_053_109, w_013_032, w_025_292);
  or2  I053_112(w_053_112, w_002_432, w_002_158);
  or2  I053_145(w_053_145, w_003_176, w_049_454);
  not1 I053_151(w_053_151, w_039_336);
  and2 I053_175(w_053_175, w_012_276, w_025_282);
  not1 I053_181(w_053_181, w_034_018);
  not1 I053_193(w_053_193, w_043_014);
  not1 I053_230(w_053_230, w_016_305);
  or2  I053_236(w_053_236, w_048_348, w_011_266);
  not1 I053_238(w_053_238, w_024_128);
  not1 I053_289(w_053_289, w_005_361);
  nand2 I053_292(w_053_292, w_018_146, w_036_217);
  or2  I053_297(w_053_297, w_051_318, w_034_672);
  and2 I053_300(w_053_300, w_040_302, w_051_457);
  not1 I053_310(w_053_310, w_028_472);
  and2 I053_341(w_053_341, w_046_184, w_015_026);
  or2  I053_346(w_053_346, w_031_438, w_012_157);
  not1 I053_364(w_053_364, w_012_136);
  or2  I053_377(w_053_377, w_045_548, w_011_178);
  and2 I053_388(w_053_388, w_034_197, w_038_009);
  nand2 I053_391(w_053_391, w_031_057, w_025_239);
  and2 I053_400(w_053_400, w_050_100, w_000_453);
  not1 I053_404(w_053_404, w_037_096);
  and2 I053_425(w_053_425, w_017_008, w_009_016);
  not1 I053_437(w_053_437, w_033_721);
  nand2 I053_456(w_053_456, w_030_387, w_003_219);
  nand2 I053_492(w_053_492, w_006_170, w_050_068);
  nand2 I053_515(w_053_515, w_009_022, w_043_021);
  not1 I053_526(w_053_526, w_045_128);
  nand2 I053_528(w_053_528, w_025_514, w_021_123);
  and2 I053_533(w_053_533, w_041_102, w_052_162);
  nand2 I053_551(w_053_551, w_015_643, w_013_421);
  not1 I053_562(w_053_562, w_034_116);
  or2  I053_575(w_053_575, w_032_146, w_043_035);
  nand2 I053_582(w_053_582, w_046_525, w_032_585);
  nand2 I053_587(w_053_587, w_025_003, w_027_007);
  and2 I053_592(w_053_592, w_006_288, w_007_276);
  not1 I053_616(w_053_616, w_043_051);
  not1 I053_645(w_053_645, w_032_162);
  or2  I053_647(w_053_647, w_023_559, w_011_154);
  and2 I053_654(w_053_654, w_020_043, w_007_537);
  not1 I053_655(w_053_655, w_045_252);
  and2 I053_676(w_053_676, w_031_183, w_006_111);
  nand2 I053_677(w_053_677, w_003_013, w_046_176);
  not1 I053_707(w_053_707, w_013_161);
  and2 I053_729(w_053_729, w_011_564, w_024_351);
  nand2 I053_733(w_053_733, w_016_437, w_012_451);
  or2  I053_735(w_053_735, w_011_281, w_002_373);
  or2  I053_760(w_053_760, w_027_466, w_004_028);
  not1 I053_763(w_053_763, w_026_377);
  and2 I053_816(w_053_816, w_047_379, w_014_217);
  or2  I053_824(w_053_824, w_041_023, w_026_296);
  and2 I053_835(w_053_835, w_036_102, w_010_321);
  not1 I053_837(w_053_837, w_026_326);
  nand2 I054_008(w_054_008, w_028_544, w_017_007);
  and2 I054_009(w_054_009, w_017_017, w_040_210);
  not1 I054_014(w_054_014, w_027_067);
  not1 I054_015(w_054_015, w_001_611);
  nand2 I054_016(w_054_016, w_003_034, w_020_098);
  not1 I054_017(w_054_017, w_033_345);
  and2 I054_020(w_054_020, w_034_042, w_033_007);
  not1 I054_023(w_054_023, w_041_057);
  nand2 I054_029(w_054_029, w_037_149, w_010_054);
  or2  I054_034(w_054_034, w_025_125, w_002_175);
  nand2 I054_035(w_054_035, w_028_890, w_041_009);
  nand2 I054_041(w_054_041, w_027_259, w_018_143);
  not1 I054_054(w_054_054, w_000_953);
  and2 I054_058(w_054_058, w_042_084, w_017_003);
  or2  I054_060(w_054_060, w_024_287, w_033_004);
  nand2 I054_077(w_054_077, w_013_002, w_019_027);
  or2  I054_079(w_054_079, w_013_263, w_039_385);
  not1 I054_080(w_054_080, w_038_345);
  not1 I054_081(w_054_081, w_022_280);
  nand2 I054_084(w_054_084, w_012_266, w_011_102);
  not1 I054_085(w_054_085, w_022_185);
  not1 I054_086(w_054_086, w_039_405);
  nand2 I054_089(w_054_089, w_039_201, w_053_012);
  or2  I054_102(w_054_102, w_017_014, w_033_030);
  nand2 I054_110(w_054_110, w_040_320, w_040_068);
  not1 I054_112(w_054_112, w_042_045);
  and2 I054_116(w_054_116, w_023_139, w_022_033);
  or2  I054_126(w_054_126, w_000_980, w_004_030);
  and2 I054_128(w_054_128, w_036_276, w_017_025);
  and2 I054_134(w_054_134, w_016_423, w_012_080);
  not1 I054_141(w_054_141, w_022_198);
  not1 I054_147(w_054_147, w_031_391);
  and2 I054_152(w_054_152, w_017_024, w_005_257);
  not1 I054_160(w_054_160, w_031_365);
  or2  I054_163(w_054_163, w_047_481, w_003_019);
  not1 I054_165(w_054_165, w_014_252);
  or2  I054_167(w_054_167, w_020_080, w_010_329);
  and2 I054_170(w_054_170, w_051_129, w_023_172);
  not1 I054_179(w_054_179, w_034_093);
  or2  I054_180(w_054_180, w_010_110, w_022_446);
  nand2 I054_185(w_054_185, w_015_130, w_041_121);
  nand2 I054_191(w_054_191, w_024_171, w_050_039);
  not1 I054_195(w_054_195, w_041_002);
  not1 I054_196(w_054_196, w_051_288);
  and2 I054_200(w_054_200, w_025_530, w_008_244);
  and2 I054_201(w_054_201, w_041_073, w_030_080);
  and2 I054_203(w_054_203, w_031_023, w_040_048);
  nand2 I054_209(w_054_209, w_036_228, w_005_001);
  and2 I054_210(w_054_210, w_053_092, w_018_093);
  not1 I054_214(w_054_214, w_003_201);
  not1 I054_215(w_054_215, w_016_104);
  nand2 I054_216(w_054_216, w_049_412, w_051_249);
  nand2 I054_217(w_054_217, w_047_158, w_047_157);
  nand2 I054_218(w_054_218, w_042_028, w_004_006);
  or2  I054_221(w_054_221, w_049_534, w_046_545);
  and2 I054_227(w_054_227, w_002_430, w_038_747);
  not1 I054_234(w_054_234, w_001_620);
  or2  I054_240(w_054_240, w_038_559, w_014_315);
  not1 I054_246(w_054_246, w_028_017);
  nand2 I054_249(w_054_249, w_006_100, w_053_377);
  nand2 I054_251(w_054_251, w_006_316, w_033_629);
  not1 I054_253(w_054_253, w_045_229);
  or2  I054_255(w_054_255, w_010_807, w_022_260);
  not1 I055_000(w_055_000, w_004_010);
  and2 I055_001(w_055_001, w_049_298, w_041_122);
  not1 I055_010(w_055_010, w_024_404);
  and2 I055_011(w_055_011, w_032_556, w_052_106);
  not1 I055_017(w_055_017, w_013_097);
  nand2 I055_022(w_055_022, w_010_413, w_005_085);
  or2  I055_033(w_055_033, w_050_005, w_046_122);
  nand2 I055_035(w_055_035, w_014_168, w_049_147);
  or2  I055_055(w_055_055, w_020_099, w_038_172);
  or2  I055_065(w_055_065, w_026_131, w_000_292);
  and2 I055_071(w_055_071, w_054_015, w_031_319);
  or2  I055_080(w_055_080, w_043_021, w_044_384);
  nand2 I055_081(w_055_081, w_016_337, w_001_136);
  nand2 I055_105(w_055_105, w_054_041, w_007_343);
  or2  I055_129(w_055_129, w_005_193, w_012_431);
  nand2 I055_138(w_055_138, w_002_234, w_051_115);
  nand2 I055_159(w_055_159, w_045_206, w_052_058);
  and2 I055_163(w_055_163, w_028_119, w_025_008);
  and2 I055_174(w_055_174, w_012_330, w_043_019);
  or2  I055_176(w_055_176, w_014_085, w_008_949);
  nand2 I055_183(w_055_183, w_039_392, w_029_160);
  not1 I055_192(w_055_192, w_007_237);
  and2 I055_194(w_055_194, w_030_444, w_016_422);
  nand2 I055_210(w_055_210, w_026_235, w_027_565);
  not1 I055_223(w_055_223, w_040_112);
  nand2 I055_233(w_055_233, w_016_048, w_003_068);
  and2 I055_245(w_055_245, w_010_773, w_031_374);
  nand2 I055_250(w_055_250, w_041_054, w_042_017);
  not1 I055_261(w_055_261, w_045_005);
  and2 I055_311(w_055_311, w_023_499, w_000_201);
  or2  I055_319(w_055_319, w_026_280, w_026_142);
  or2  I055_336(w_055_336, w_002_046, w_000_612);
  not1 I055_358(w_055_358, w_006_051);
  not1 I055_375(w_055_375, w_034_241);
  not1 I055_398(w_055_398, w_021_190);
  and2 I055_474(w_055_474, w_037_027, w_011_004);
  not1 I055_500(w_055_500, w_043_007);
  and2 I055_503(w_055_503, w_017_027, w_026_014);
  nand2 I055_529(w_055_529, w_036_023, w_004_005);
  or2  I055_548(w_055_548, w_047_212, w_023_234);
  nand2 I055_574(w_055_574, w_030_196, w_050_301);
  and2 I055_593(w_055_593, w_014_405, w_041_113);
  not1 I055_594(w_055_594, w_021_194);
  and2 I055_596(w_055_596, w_016_208, w_014_434);
  not1 I055_603(w_055_603, w_025_105);
  or2  I055_607(w_055_607, w_052_006, w_022_358);
  not1 I055_611(w_055_611, w_052_023);
  or2  I055_615(w_055_615, w_011_014, w_022_479);
  nand2 I055_664(w_055_664, w_020_013, w_012_197);
  or2  I055_688(w_055_688, w_053_089, w_008_482);
  nand2 I055_723(w_055_723, w_054_210, w_033_307);
  or2  I055_731(w_055_731, w_004_024, w_021_010);
  or2  I055_732(w_055_732, w_029_214, w_002_118);
  not1 I055_744(w_055_744, w_039_305);
  or2  I055_762(w_055_762, w_024_141, w_008_305);
  or2  I056_003(w_056_003, w_013_146, w_050_344);
  and2 I056_004(w_056_004, w_054_034, w_029_067);
  or2  I056_007(w_056_007, w_009_000, w_039_382);
  or2  I056_010(w_056_010, w_040_149, w_049_383);
  nand2 I056_012(w_056_012, w_010_332, w_026_264);
  or2  I056_022(w_056_022, w_047_295, w_044_039);
  nand2 I056_034(w_056_034, w_033_815, w_042_041);
  and2 I056_039(w_056_039, w_048_384, w_033_016);
  nand2 I056_045(w_056_045, w_010_426, w_007_067);
  or2  I056_048(w_056_048, w_034_123, w_030_340);
  or2  I056_065(w_056_065, w_046_642, w_039_371);
  not1 I056_077(w_056_077, w_015_124);
  nand2 I056_081(w_056_081, w_040_182, w_006_220);
  nand2 I056_086(w_056_086, w_040_259, w_026_353);
  not1 I056_088(w_056_088, w_041_049);
  and2 I056_092(w_056_092, w_017_001, w_051_372);
  not1 I056_096(w_056_096, w_044_075);
  or2  I056_099(w_056_099, w_030_046, w_049_691);
  nand2 I056_112(w_056_112, w_009_052, w_024_323);
  nand2 I056_125(w_056_125, w_044_067, w_030_461);
  not1 I056_128(w_056_128, w_026_180);
  or2  I056_166(w_056_166, w_037_055, w_027_826);
  nand2 I056_170(w_056_170, w_011_143, w_037_142);
  not1 I056_175(w_056_175, w_033_613);
  nand2 I056_177(w_056_177, w_003_115, w_030_480);
  not1 I056_187(w_056_187, w_041_101);
  and2 I056_188(w_056_188, w_000_215, w_040_084);
  or2  I056_190(w_056_190, w_007_020, w_035_578);
  or2  I056_193(w_056_193, w_045_106, w_024_426);
  and2 I056_196(w_056_196, w_037_016, w_048_803);
  nand2 I056_212(w_056_212, w_041_032, w_021_170);
  and2 I056_219(w_056_219, w_000_624, w_023_445);
  and2 I056_227(w_056_227, w_008_878, w_019_097);
  nand2 I056_228(w_056_228, w_043_065, w_015_124);
  not1 I056_231(w_056_231, w_051_223);
  nand2 I056_235(w_056_235, w_033_202, w_049_828);
  and2 I056_236(w_056_236, w_012_288, w_021_050);
  not1 I056_255(w_056_255, w_051_356);
  or2  I056_256(w_056_256, w_010_247, w_009_042);
  not1 I056_275(w_056_275, w_024_416);
  not1 I056_279(w_056_279, w_019_165);
  or2  I056_280(w_056_280, w_054_008, w_020_092);
  nand2 I056_284(w_056_284, w_001_360, w_028_715);
  or2  I056_285(w_056_285, w_034_104, w_000_749);
  nand2 I056_299(w_056_299, w_031_178, w_025_125);
  and2 I056_311(w_056_311, w_044_162, w_002_271);
  and2 I057_002(w_057_002, w_046_158, w_004_007);
  nand2 I057_008(w_057_008, w_012_413, w_029_136);
  and2 I057_010(w_057_010, w_054_110, w_014_308);
  nand2 I057_017(w_057_017, w_028_783, w_002_123);
  and2 I057_021(w_057_021, w_053_763, w_054_126);
  nand2 I057_023(w_057_023, w_022_010, w_016_275);
  not1 I057_024(w_057_024, w_044_120);
  and2 I057_031(w_057_031, w_017_026, w_040_116);
  and2 I057_039(w_057_039, w_050_250, w_006_149);
  not1 I057_041(w_057_041, w_048_095);
  not1 I057_043(w_057_043, w_022_174);
  and2 I057_050(w_057_050, w_055_261, w_004_030);
  or2  I057_051(w_057_051, w_022_325, w_038_565);
  or2  I057_063(w_057_063, w_007_417, w_016_128);
  and2 I057_067(w_057_067, w_037_012, w_007_078);
  not1 I057_091(w_057_091, w_003_086);
  not1 I057_092(w_057_092, w_026_308);
  or2  I057_102(w_057_102, w_054_201, w_005_060);
  and2 I057_113(w_057_113, w_024_229, w_001_363);
  and2 I057_121(w_057_121, w_023_309, w_014_435);
  and2 I057_122(w_057_122, w_054_152, w_003_038);
  not1 I057_145(w_057_145, w_015_003);
  not1 I057_154(w_057_154, w_053_533);
  and2 I057_157(w_057_157, w_001_156, w_042_001);
  not1 I057_167(w_057_167, w_007_328);
  nand2 I057_169(w_057_169, w_025_585, w_034_785);
  or2  I057_190(w_057_190, w_001_034, w_006_057);
  not1 I057_198(w_057_198, w_009_062);
  nand2 I057_200(w_057_200, w_018_196, w_037_180);
  not1 I057_202(w_057_202, w_041_118);
  not1 I057_209(w_057_209, w_037_008);
  not1 I057_210(w_057_210, w_008_764);
  or2  I057_233(w_057_233, w_029_123, w_015_365);
  nand2 I057_252(w_057_252, w_002_055, w_025_066);
  or2  I057_253(w_057_253, w_043_061, w_025_555);
  and2 I057_256(w_057_256, w_002_313, w_028_629);
  not1 I057_262(w_057_262, w_036_266);
  not1 I057_275(w_057_275, w_049_629);
  nand2 I057_305(w_057_305, w_032_716, w_006_095);
  and2 I057_311(w_057_311, w_017_025, w_008_951);
  not1 I057_316(w_057_316, w_035_631);
  nand2 I057_322(w_057_322, w_008_071, w_045_339);
  or2  I057_323(w_057_323, w_051_037, w_054_084);
  or2  I057_325(w_057_325, w_043_005, w_004_037);
  not1 I057_336(w_057_336, w_041_117);
  nand2 I057_337(w_057_337, w_056_128, w_023_621);
  not1 I057_350(w_057_350, w_043_060);
  and2 I057_353(w_057_353, w_030_390, w_034_214);
  nand2 I057_357(w_057_357, w_004_013, w_023_666);
  not1 I057_385(w_057_385, w_007_358);
  and2 I057_393(w_057_393, w_019_275, w_001_157);
  nand2 I057_397(w_057_397, w_030_206, w_026_231);
  nand2 I057_403(w_057_403, w_009_008, w_035_374);
  not1 I057_415(w_057_415, w_038_046);
  nand2 I057_417(w_057_417, w_001_038, w_012_102);
  and2 I057_425(w_057_425, w_048_136, w_054_116);
  or2  I057_435(w_057_435, w_005_454, w_018_096);
  nand2 I057_443(w_057_443, w_009_002, w_006_310);
  and2 I057_445(w_057_445, w_029_115, w_017_007);
  nand2 I057_467(w_057_467, w_031_294, w_044_292);
  or2  I058_002(w_058_002, w_008_247, w_008_760);
  nand2 I058_006(w_058_006, w_045_006, w_003_169);
  and2 I058_009(w_058_009, w_053_677, w_013_048);
  and2 I058_010(w_058_010, w_045_567, w_053_022);
  or2  I058_015(w_058_015, w_048_559, w_023_190);
  nand2 I058_040(w_058_040, w_029_050, w_036_260);
  not1 I058_050(w_058_050, w_026_368);
  nand2 I058_058(w_058_058, w_018_131, w_008_486);
  not1 I058_064(w_058_064, w_041_003);
  or2  I058_065(w_058_065, w_001_703, w_001_151);
  and2 I058_070(w_058_070, w_019_118, w_044_047);
  and2 I058_071(w_058_071, w_037_114, w_033_294);
  and2 I058_072(w_058_072, w_017_011, w_044_315);
  not1 I058_080(w_058_080, w_000_430);
  and2 I058_085(w_058_085, w_004_035, w_004_010);
  and2 I058_086(w_058_086, w_033_190, w_037_013);
  and2 I058_094(w_058_094, w_014_529, w_030_010);
  and2 I058_097(w_058_097, w_017_003, w_045_111);
  and2 I058_108(w_058_108, w_030_082, w_039_265);
  and2 I058_112(w_058_112, w_025_668, w_043_011);
  and2 I058_115(w_058_115, w_052_037, w_055_593);
  nand2 I058_123(w_058_123, w_011_155, w_001_259);
  not1 I058_128(w_058_128, w_045_593);
  nand2 I058_139(w_058_139, w_046_421, w_037_109);
  not1 I058_140(w_058_140, w_021_210);
  or2  I058_151(w_058_151, w_014_411, w_019_233);
  nand2 I058_154(w_058_154, w_017_001, w_019_200);
  not1 I058_155(w_058_155, w_027_272);
  nand2 I058_167(w_058_167, w_015_693, w_049_478);
  nand2 I058_172(w_058_172, w_015_096, w_002_333);
  and2 I058_176(w_058_176, w_024_014, w_014_115);
  not1 I058_177(w_058_177, w_006_187);
  or2  I058_179(w_058_179, w_027_091, w_016_496);
  nand2 I058_182(w_058_182, w_005_327, w_051_075);
  and2 I058_190(w_058_190, w_029_199, w_029_087);
  nand2 I058_191(w_058_191, w_016_323, w_048_201);
  nand2 I058_196(w_058_196, w_045_531, w_043_054);
  or2  I058_197(w_058_197, w_036_131, w_016_016);
  and2 I058_199(w_058_199, w_050_299, w_041_096);
  not1 I058_205(w_058_205, w_026_040);
  not1 I058_215(w_058_215, w_054_215);
  not1 I058_220(w_058_220, w_009_004);
  and2 I058_221(w_058_221, w_040_008, w_042_045);
  and2 I058_225(w_058_225, w_041_070, w_054_102);
  not1 I058_227(w_058_227, w_055_398);
  nand2 I058_233(w_058_233, w_023_157, w_035_518);
  nand2 I058_238(w_058_238, w_018_116, w_010_072);
  and2 I058_239(w_058_239, w_033_049, w_015_350);
  and2 I058_247(w_058_247, w_018_053, w_002_022);
  or2  I058_250(w_058_250, w_001_138, w_052_064);
  nand2 I058_281(w_058_281, w_057_102, w_003_033);
  and2 I058_292(w_058_292, w_030_391, w_003_028);
  not1 I058_302(w_058_302, w_057_256);
  and2 I058_317(w_058_317, w_052_129, w_046_195);
  and2 I058_320(w_058_320, w_024_592, w_015_025);
  or2  I058_324(w_058_324, w_052_017, w_039_003);
  and2 I058_335(w_058_335, w_047_095, w_020_129);
  not1 I058_341(w_058_341, w_049_883);
  and2 I058_347(w_058_347, w_020_028, w_032_596);
  not1 I058_360(w_058_360, w_021_259);
  not1 I059_018(w_059_018, w_058_335);
  and2 I059_028(w_059_028, w_044_015, w_058_058);
  not1 I059_030(w_059_030, w_047_448);
  nand2 I059_032(w_059_032, w_051_314, w_017_020);
  nand2 I059_044(w_059_044, w_005_201, w_028_210);
  nand2 I059_047(w_059_047, w_031_055, w_057_233);
  not1 I059_058(w_059_058, w_015_168);
  and2 I059_068(w_059_068, w_050_215, w_045_328);
  nand2 I059_076(w_059_076, w_040_057, w_006_147);
  and2 I059_090(w_059_090, w_037_047, w_039_146);
  or2  I059_092(w_059_092, w_002_290, w_027_016);
  or2  I059_094(w_059_094, w_029_202, w_057_336);
  and2 I059_097(w_059_097, w_010_052, w_051_108);
  and2 I059_105(w_059_105, w_039_459, w_027_736);
  not1 I059_116(w_059_116, w_057_417);
  nand2 I059_121(w_059_121, w_026_383, w_024_209);
  and2 I059_123(w_059_123, w_058_112, w_047_118);
  and2 I059_134(w_059_134, w_016_337, w_005_093);
  nand2 I059_135(w_059_135, w_029_119, w_018_118);
  and2 I059_138(w_059_138, w_033_124, w_055_311);
  or2  I059_142(w_059_142, w_036_043, w_015_713);
  and2 I059_143(w_059_143, w_009_033, w_054_214);
  and2 I059_145(w_059_145, w_036_197, w_004_013);
  and2 I059_146(w_059_146, w_049_246, w_022_039);
  and2 I059_147(w_059_147, w_000_554, w_055_176);
  not1 I059_149(w_059_149, w_055_250);
  or2  I059_151(w_059_151, w_052_100, w_006_000);
  nand2 I059_152(w_059_152, w_032_179, w_009_019);
  or2  I059_154(w_059_154, w_024_019, w_035_212);
  nand2 I059_164(w_059_164, w_003_096, w_006_221);
  nand2 I059_169(w_059_169, w_013_426, w_008_158);
  not1 I059_177(w_059_177, w_022_400);
  or2  I059_179(w_059_179, w_004_012, w_000_078);
  nand2 I059_180(w_059_180, w_029_061, w_055_174);
  not1 I059_192(w_059_192, w_021_006);
  and2 I059_193(w_059_193, w_042_069, w_020_016);
  nand2 I059_209(w_059_209, w_006_187, w_028_241);
  or2  I059_213(w_059_213, w_027_537, w_049_329);
  and2 I059_214(w_059_214, w_041_077, w_009_012);
  or2  I059_224(w_059_224, w_025_657, w_044_058);
  and2 I059_230(w_059_230, w_043_025, w_006_329);
  or2  I059_235(w_059_235, w_055_744, w_002_291);
  and2 I059_237(w_059_237, w_023_659, w_005_090);
  not1 I059_245(w_059_245, w_023_348);
  nand2 I059_247(w_059_247, w_042_064, w_007_437);
  nand2 I059_258(w_059_258, w_050_438, w_058_097);
  and2 I059_263(w_059_263, w_051_023, w_025_419);
  nand2 I059_264(w_059_264, w_037_099, w_007_203);
  nand2 I059_272(w_059_272, w_004_033, w_036_090);
  not1 I059_277(w_059_277, w_058_179);
  not1 I059_278(w_059_278, w_034_092);
  and2 I059_279(w_059_279, w_003_143, w_023_200);
  or2  I059_282(w_059_282, w_008_361, w_025_648);
  or2  I059_308(w_059_308, w_036_097, w_026_034);
  and2 I059_317(w_059_317, w_044_227, w_016_425);
  or2  I059_318(w_059_318, w_016_186, w_015_624);
  and2 I059_333(w_059_333, w_025_215, w_000_574);
  nand2 I060_012(w_060_012, w_012_256, w_054_081);
  not1 I060_018(w_060_018, w_051_299);
  and2 I060_024(w_060_024, w_012_101, w_032_204);
  nand2 I060_035(w_060_035, w_034_666, w_014_190);
  or2  I060_057(w_060_057, w_046_091, w_059_097);
  and2 I060_071(w_060_071, w_000_480, w_004_030);
  or2  I060_095(w_060_095, w_045_415, w_013_433);
  and2 I060_101(w_060_101, w_007_011, w_045_145);
  nand2 I060_105(w_060_105, w_052_007, w_039_125);
  and2 I060_120(w_060_120, w_047_262, w_024_268);
  and2 I060_134(w_060_134, w_013_450, w_023_429);
  not1 I060_142(w_060_142, w_054_255);
  and2 I060_153(w_060_153, w_001_229, w_048_070);
  nand2 I060_155(w_060_155, w_021_130, w_011_596);
  not1 I060_165(w_060_165, w_017_006);
  nand2 I060_171(w_060_171, w_059_164, w_026_266);
  not1 I060_173(w_060_173, w_039_431);
  not1 I060_178(w_060_178, w_004_021);
  or2  I060_183(w_060_183, w_052_102, w_058_139);
  and2 I060_185(w_060_185, w_005_024, w_052_030);
  and2 I060_189(w_060_189, w_009_000, w_007_219);
  nand2 I060_212(w_060_212, w_035_214, w_056_004);
  nand2 I060_213(w_060_213, w_046_324, w_041_007);
  and2 I060_215(w_060_215, w_011_056, w_045_192);
  and2 I060_229(w_060_229, w_051_327, w_040_331);
  or2  I060_240(w_060_240, w_047_247, w_033_182);
  nand2 I060_241(w_060_241, w_054_200, w_045_692);
  and2 I060_242(w_060_242, w_003_134, w_023_334);
  not1 I060_246(w_060_246, w_026_328);
  and2 I060_247(w_060_247, w_044_365, w_038_694);
  not1 I060_249(w_060_249, w_044_371);
  and2 I060_257(w_060_257, w_054_112, w_047_332);
  or2  I060_260(w_060_260, w_053_655, w_009_034);
  and2 I060_263(w_060_263, w_012_369, w_032_658);
  not1 I060_269(w_060_269, w_007_489);
  or2  I060_288(w_060_288, w_015_205, w_050_083);
  not1 I060_297(w_060_297, w_033_192);
  not1 I060_301(w_060_301, w_023_588);
  nand2 I060_305(w_060_305, w_046_156, w_012_042);
  not1 I060_307(w_060_307, w_052_078);
  nand2 I060_311(w_060_311, w_058_123, w_041_077);
  not1 I060_313(w_060_313, w_033_372);
  nand2 I060_316(w_060_316, w_007_097, w_010_583);
  and2 I060_320(w_060_320, w_055_732, w_045_467);
  and2 I060_323(w_060_323, w_034_087, w_035_003);
  or2  I060_331(w_060_331, w_031_187, w_059_143);
  or2  I060_341(w_060_341, w_011_223, w_036_111);
  nand2 I061_009(w_061_009, w_038_122, w_049_470);
  not1 I061_017(w_061_017, w_018_034);
  nand2 I061_023(w_061_023, w_005_233, w_051_069);
  not1 I061_033(w_061_033, w_026_073);
  not1 I061_034(w_061_034, w_019_359);
  nand2 I061_045(w_061_045, w_017_008, w_054_180);
  not1 I061_052(w_061_052, w_054_195);
  nand2 I061_055(w_061_055, w_033_071, w_010_798);
  or2  I061_063(w_061_063, w_036_080, w_040_027);
  or2  I061_069(w_061_069, w_051_196, w_021_064);
  not1 I061_070(w_061_070, w_050_088);
  or2  I061_071(w_061_071, w_027_225, w_042_059);
  not1 I061_078(w_061_078, w_031_150);
  not1 I061_095(w_061_095, w_044_312);
  not1 I061_123(w_061_123, w_056_175);
  nand2 I061_132(w_061_132, w_018_175, w_021_106);
  and2 I061_147(w_061_147, w_037_107, w_028_311);
  not1 I061_168(w_061_168, w_033_193);
  and2 I061_172(w_061_172, w_050_389, w_003_050);
  or2  I061_174(w_061_174, w_004_001, w_056_034);
  not1 I061_216(w_061_216, w_038_644);
  nand2 I061_221(w_061_221, w_052_060, w_025_613);
  or2  I061_222(w_061_222, w_025_036, w_044_024);
  or2  I061_235(w_061_235, w_046_461, w_027_797);
  not1 I061_238(w_061_238, w_054_029);
  nand2 I061_241(w_061_241, w_037_171, w_009_000);
  nand2 I061_245(w_061_245, w_021_245, w_021_163);
  or2  I061_247(w_061_247, w_057_154, w_055_319);
  not1 I061_250(w_061_250, w_003_171);
  and2 I061_254(w_061_254, w_027_497, w_028_848);
  not1 I061_255(w_061_255, w_002_160);
  or2  I061_257(w_061_257, w_037_016, w_017_016);
  nand2 I061_267(w_061_267, w_030_234, w_022_034);
  and2 I061_283(w_061_283, w_005_470, w_042_068);
  and2 I061_286(w_061_286, w_017_005, w_003_202);
  nand2 I061_298(w_061_298, w_009_000, w_028_087);
  nand2 I061_300(w_061_300, w_040_141, w_049_623);
  not1 I061_331(w_061_331, w_042_050);
  or2  I061_333(w_061_333, w_041_008, w_023_462);
  not1 I061_355(w_061_355, w_027_426);
  or2  I061_360(w_061_360, w_044_274, w_047_232);
  nand2 I061_377(w_061_377, w_004_002, w_031_085);
  nand2 I061_379(w_061_379, w_021_222, w_036_134);
  and2 I061_380(w_061_380, w_053_042, w_032_092);
  nand2 I061_394(w_061_394, w_007_195, w_002_068);
  and2 I061_403(w_061_403, w_039_460, w_024_292);
  or2  I061_410(w_061_410, w_058_140, w_007_165);
  or2  I061_414(w_061_414, w_046_674, w_026_395);
  not1 I061_432(w_061_432, w_037_145);
  not1 I061_433(w_061_433, w_033_315);
  and2 I061_461(w_061_461, w_041_017, w_006_275);
  and2 I061_478(w_061_478, w_052_152, w_060_018);
  and2 I061_490(w_061_490, w_057_435, w_024_398);
  nand2 I061_497(w_061_497, w_025_362, w_049_516);
  not1 I061_502(w_061_502, w_039_062);
  nand2 I061_528(w_061_528, w_028_171, w_060_215);
  or2  I061_560(w_061_560, w_025_314, w_027_101);
  and2 I062_021(w_062_021, w_030_064, w_013_416);
  nand2 I062_022(w_062_022, w_042_081, w_028_631);
  nand2 I062_029(w_062_029, w_038_324, w_059_245);
  and2 I062_031(w_062_031, w_022_307, w_059_094);
  or2  I062_032(w_062_032, w_014_282, w_055_500);
  nand2 I062_037(w_062_037, w_014_032, w_042_005);
  or2  I062_069(w_062_069, w_037_111, w_018_167);
  not1 I062_100(w_062_100, w_047_082);
  and2 I062_121(w_062_121, w_024_284, w_041_115);
  and2 I062_124(w_062_124, w_044_341, w_048_493);
  and2 I062_140(w_062_140, w_019_249, w_044_118);
  or2  I062_149(w_062_149, w_032_268, w_011_013);
  or2  I062_165(w_062_165, w_044_114, w_024_321);
  or2  I062_166(w_062_166, w_026_030, w_026_062);
  not1 I062_167(w_062_167, w_017_010);
  nand2 I062_174(w_062_174, w_053_582, w_023_603);
  or2  I062_228(w_062_228, w_034_433, w_017_025);
  nand2 I062_240(w_062_240, w_038_469, w_023_307);
  nand2 I062_251(w_062_251, w_022_439, w_023_416);
  nand2 I062_252(w_062_252, w_033_040, w_038_305);
  and2 I062_253(w_062_253, w_020_128, w_046_059);
  or2  I062_272(w_062_272, w_009_066, w_037_039);
  nand2 I062_280(w_062_280, w_025_047, w_058_205);
  and2 I062_292(w_062_292, w_000_559, w_045_421);
  nand2 I062_300(w_062_300, w_003_175, w_060_120);
  or2  I062_312(w_062_312, w_003_161, w_039_299);
  nand2 I062_314(w_062_314, w_024_515, w_004_002);
  nand2 I062_353(w_062_353, w_049_327, w_025_535);
  and2 I062_371(w_062_371, w_058_112, w_051_102);
  not1 I062_373(w_062_373, w_007_316);
  nand2 I062_374(w_062_374, w_028_899, w_002_173);
  nand2 I062_386(w_062_386, w_026_011, w_058_115);
  or2  I062_428(w_062_428, w_013_025, w_040_098);
  nand2 I062_432(w_062_432, w_041_031, w_021_099);
  nand2 I062_436(w_062_436, w_058_239, w_042_068);
  and2 I062_440(w_062_440, w_013_469, w_025_090);
  or2  I062_469(w_062_469, w_012_420, w_022_495);
  or2  I062_471(w_062_471, w_056_034, w_035_230);
  nand2 I062_474(w_062_474, w_032_546, w_042_094);
  or2  I062_478(w_062_478, w_054_216, w_028_590);
  and2 I062_479(w_062_479, w_057_415, w_024_555);
  nand2 I063_027(w_063_027, w_052_109, w_047_187);
  and2 I063_037(w_063_037, w_047_033, w_017_003);
  not1 I063_038(w_063_038, w_061_132);
  and2 I063_053(w_063_053, w_010_640, w_034_091);
  and2 I063_054(w_063_054, w_023_253, w_004_009);
  not1 I063_059(w_063_059, w_060_142);
  not1 I063_064(w_063_064, w_047_158);
  nand2 I063_071(w_063_071, w_007_244, w_061_410);
  or2  I063_081(w_063_081, w_011_146, w_059_105);
  and2 I063_083(w_063_083, w_047_096, w_053_562);
  not1 I063_084(w_063_084, w_022_315);
  not1 I063_085(w_063_085, w_034_583);
  and2 I063_098(w_063_098, w_045_511, w_020_104);
  nand2 I063_099(w_063_099, w_019_100, w_046_006);
  or2  I063_103(w_063_103, w_011_205, w_006_187);
  not1 I063_104(w_063_104, w_033_548);
  nand2 I063_107(w_063_107, w_041_099, w_052_147);
  or2  I063_110(w_063_110, w_003_155, w_044_031);
  and2 I063_119(w_063_119, w_003_090, w_053_400);
  or2  I063_130(w_063_130, w_055_375, w_053_575);
  and2 I063_133(w_063_133, w_034_023, w_034_177);
  or2  I063_135(w_063_135, w_049_835, w_051_138);
  nand2 I063_138(w_063_138, w_050_423, w_031_406);
  or2  I063_146(w_063_146, w_020_058, w_038_206);
  nand2 I063_162(w_063_162, w_001_187, w_028_494);
  nand2 I063_181(w_063_181, w_024_084, w_015_496);
  or2  I063_193(w_063_193, w_024_096, w_017_016);
  and2 I063_195(w_063_195, w_048_018, w_050_469);
  or2  I063_198(w_063_198, w_040_347, w_013_459);
  and2 I063_200(w_063_200, w_008_771, w_020_011);
  not1 I063_201(w_063_201, w_056_193);
  nand2 I063_204(w_063_204, w_014_527, w_000_488);
  nand2 I063_205(w_063_205, w_023_041, w_021_219);
  or2  I063_210(w_063_210, w_018_034, w_035_313);
  or2  I063_212(w_063_212, w_032_234, w_002_292);
  or2  I063_215(w_063_215, w_041_033, w_037_162);
  nand2 I063_216(w_063_216, w_052_099, w_055_183);
  and2 I063_217(w_063_217, w_022_243, w_010_170);
  nand2 I063_225(w_063_225, w_034_068, w_048_227);
  and2 I063_226(w_063_226, w_004_024, w_041_076);
  and2 I063_231(w_063_231, w_019_069, w_055_358);
  not1 I063_242(w_063_242, w_021_035);
  or2  I063_258(w_063_258, w_052_026, w_006_258);
  or2  I063_260(w_063_260, w_040_113, w_001_030);
  nand2 I063_266(w_063_266, w_027_543, w_040_178);
  or2  I063_274(w_063_274, w_014_275, w_004_023);
  and2 I063_286(w_063_286, w_008_461, w_025_280);
  or2  I063_287(w_063_287, w_024_570, w_031_382);
  not1 I063_290(w_063_290, w_046_497);
  or2  I063_293(w_063_293, w_022_286, w_010_736);
  and2 I063_303(w_063_303, w_014_006, w_055_065);
  and2 I063_315(w_063_315, w_010_346, w_036_036);
  nand2 I063_322(w_063_322, w_050_244, w_053_837);
  nand2 I063_353(w_063_353, w_028_468, w_009_062);
  not1 I063_357(w_063_357, w_038_735);
  not1 I063_360(w_063_360, w_014_181);
  nand2 I064_002(w_064_002, w_012_323, w_007_294);
  not1 I064_003(w_064_003, w_014_091);
  or2  I064_021(w_064_021, w_038_459, w_063_098);
  not1 I064_032(w_064_032, w_039_040);
  or2  I064_036(w_064_036, w_044_378, w_040_111);
  or2  I064_041(w_064_041, w_030_271, w_020_096);
  not1 I064_070(w_064_070, w_006_043);
  not1 I064_076(w_064_076, w_021_048);
  nand2 I064_086(w_064_086, w_032_124, w_038_190);
  not1 I064_091(w_064_091, w_008_601);
  nand2 I064_102(w_064_102, w_057_357, w_018_098);
  nand2 I064_131(w_064_131, w_031_333, w_046_420);
  not1 I064_138(w_064_138, w_044_172);
  nand2 I064_142(w_064_142, w_002_293, w_059_030);
  not1 I064_146(w_064_146, w_063_225);
  not1 I064_157(w_064_157, w_040_237);
  not1 I064_169(w_064_169, w_024_380);
  not1 I064_188(w_064_188, w_047_238);
  not1 I064_247(w_064_247, w_051_161);
  or2  I064_264(w_064_264, w_061_283, w_011_273);
  nand2 I064_271(w_064_271, w_029_011, w_050_159);
  and2 I064_277(w_064_277, w_058_094, w_039_031);
  or2  I064_311(w_064_311, w_042_070, w_054_249);
  not1 I064_338(w_064_338, w_035_134);
  nand2 I064_340(w_064_340, w_033_862, w_044_314);
  or2  I064_347(w_064_347, w_046_294, w_053_528);
  not1 I064_355(w_064_355, w_049_218);
  and2 I064_375(w_064_375, w_054_165, w_018_091);
  not1 I064_411(w_064_411, w_021_157);
  or2  I064_433(w_064_433, w_007_286, w_007_488);
  and2 I064_448(w_064_448, w_021_172, w_048_023);
  or2  I064_453(w_064_453, w_001_555, w_033_339);
  not1 I064_477(w_064_477, w_036_151);
  or2  I064_482(w_064_482, w_037_040, w_034_495);
  nand2 I064_493(w_064_493, w_047_176, w_044_133);
  nand2 I064_503(w_064_503, w_039_007, w_062_428);
  or2  I064_515(w_064_515, w_038_526, w_032_548);
  not1 I064_526(w_064_526, w_059_092);
  or2  I064_534(w_064_534, w_028_411, w_040_016);
  or2  I064_537(w_064_537, w_041_097, w_019_020);
  not1 I064_554(w_064_554, w_055_000);
  and2 I064_574(w_064_574, w_057_311, w_027_635);
  not1 I064_606(w_064_606, w_016_476);
  nand2 I064_610(w_064_610, w_028_092, w_015_021);
  not1 I064_630(w_064_630, w_018_116);
  not1 I064_637(w_064_637, w_037_187);
  nand2 I064_665(w_064_665, w_023_196, w_025_658);
  or2  I064_668(w_064_668, w_030_311, w_044_070);
  and2 I064_679(w_064_679, w_048_034, w_022_187);
  and2 I064_690(w_064_690, w_022_294, w_051_384);
  or2  I064_692(w_064_692, w_009_046, w_030_487);
  nand2 I064_695(w_064_695, w_051_404, w_001_253);
  and2 I064_727(w_064_727, w_031_212, w_054_209);
  nand2 I064_741(w_064_741, w_012_303, w_053_526);
  nand2 I064_749(w_064_749, w_016_074, w_058_167);
  not1 I064_750(w_064_750, w_060_185);
  or2  I064_789(w_064_789, w_005_252, w_040_029);
  nand2 I064_804(w_064_804, w_044_037, w_048_706);
  nand2 I064_806(w_064_806, w_045_193, w_047_470);
  and2 I064_832(w_064_832, w_001_548, w_016_290);
  or2  I065_006(w_065_006, w_043_024, w_007_532);
  not1 I065_013(w_065_013, w_056_112);
  nand2 I065_017(w_065_017, w_033_878, w_001_358);
  nand2 I065_051(w_065_051, w_008_035, w_009_055);
  not1 I065_091(w_065_091, w_012_058);
  or2  I065_094(w_065_094, w_062_374, w_002_001);
  or2  I065_095(w_065_095, w_050_002, w_008_499);
  nand2 I065_160(w_065_160, w_044_038, w_043_028);
  or2  I065_204(w_065_204, w_034_458, w_036_005);
  nand2 I065_223(w_065_223, w_004_021, w_030_450);
  and2 I065_251(w_065_251, w_055_081, w_036_222);
  not1 I065_279(w_065_279, w_021_220);
  not1 I065_305(w_065_305, w_064_411);
  and2 I065_312(w_065_312, w_026_032, w_019_085);
  and2 I065_333(w_065_333, w_002_148, w_007_265);
  not1 I065_363(w_065_363, w_019_320);
  not1 I065_373(w_065_373, w_046_559);
  or2  I065_380(w_065_380, w_006_203, w_048_816);
  or2  I065_422(w_065_422, w_048_552, w_002_134);
  not1 I065_423(w_065_423, w_057_353);
  and2 I065_433(w_065_433, w_008_586, w_043_044);
  and2 I065_509(w_065_509, w_012_491, w_042_012);
  nand2 I065_527(w_065_527, w_013_365, w_008_024);
  not1 I065_537(w_065_537, w_009_015);
  and2 I065_551(w_065_551, w_056_187, w_045_105);
  not1 I065_556(w_065_556, w_030_318);
  and2 I065_585(w_065_585, w_055_080, w_049_879);
  or2  I065_613(w_065_613, w_064_157, w_013_485);
  nand2 I065_631(w_065_631, w_025_382, w_048_479);
  not1 I065_652(w_065_652, w_059_047);
  and2 I065_665(w_065_665, w_004_023, w_006_086);
  nand2 I065_686(w_065_686, w_024_209, w_050_366);
  and2 I065_697(w_065_697, w_040_243, w_025_136);
  nand2 I065_711(w_065_711, w_001_362, w_031_090);
  not1 I065_732(w_065_732, w_004_010);
  and2 I065_740(w_065_740, w_008_355, w_035_195);
  or2  I065_742(w_065_742, w_013_181, w_055_594);
  nand2 I065_750(w_065_750, w_055_035, w_016_330);
  or2  I065_850(w_065_850, w_046_157, w_027_676);
  not1 I065_855(w_065_855, w_045_108);
  and2 I065_861(w_065_861, w_007_432, w_015_136);
  nand2 I065_883(w_065_883, w_030_182, w_005_219);
  or2  I065_895(w_065_895, w_054_035, w_014_058);
  not1 I065_914(w_065_914, w_045_067);
  or2  I065_920(w_065_920, w_003_147, w_048_335);
  nand2 I065_941(w_065_941, w_051_094, w_038_625);
  or2  I065_944(w_065_944, w_012_337, w_044_166);
  or2  I065_950(w_065_950, w_026_079, w_023_451);
  and2 I065_951(w_065_951, w_037_009, w_035_170);
  nand2 I065_972(w_065_972, w_042_083, w_001_778);
  and2 I065_978(w_065_978, w_014_167, w_028_219);
  and2 I066_014(w_066_014, w_062_292, w_007_012);
  nand2 I066_017(w_066_017, w_063_201, w_026_210);
  and2 I066_023(w_066_023, w_017_018, w_028_626);
  or2  I066_024(w_066_024, w_023_196, w_055_194);
  nand2 I066_037(w_066_037, w_060_213, w_009_047);
  not1 I066_039(w_066_039, w_005_179);
  not1 I066_051(w_066_051, w_045_141);
  and2 I066_054(w_066_054, w_063_226, w_032_188);
  and2 I066_058(w_066_058, w_016_467, w_011_657);
  nand2 I066_072(w_066_072, w_036_089, w_009_032);
  or2  I066_082(w_066_082, w_028_024, w_025_378);
  and2 I066_107(w_066_107, w_004_028, w_015_774);
  or2  I066_114(w_066_114, w_060_165, w_030_178);
  not1 I066_115(w_066_115, w_028_595);
  and2 I066_119(w_066_119, w_036_147, w_001_187);
  nand2 I066_124(w_066_124, w_028_368, w_035_078);
  and2 I066_141(w_066_141, w_047_245, w_035_540);
  or2  I066_146(w_066_146, w_021_220, w_037_098);
  not1 I066_187(w_066_187, w_008_156);
  or2  I066_202(w_066_202, w_049_654, w_040_204);
  and2 I066_209(w_066_209, w_008_236, w_044_323);
  or2  I066_210(w_066_210, w_016_047, w_064_355);
  nand2 I066_213(w_066_213, w_009_017, w_020_053);
  not1 I066_224(w_066_224, w_053_647);
  nand2 I066_249(w_066_249, w_001_655, w_026_243);
  nand2 I066_282(w_066_282, w_043_011, w_011_183);
  or2  I066_285(w_066_285, w_000_627, w_032_170);
  nand2 I066_295(w_066_295, w_065_740, w_007_277);
  nand2 I066_317(w_066_317, w_022_314, w_009_011);
  not1 I066_345(w_066_345, w_001_883);
  and2 I066_355(w_066_355, w_012_414, w_047_190);
  nand2 I066_359(w_066_359, w_003_080, w_053_297);
  and2 I066_368(w_066_368, w_058_215, w_036_021);
  not1 I066_371(w_066_371, w_057_021);
  nand2 I066_376(w_066_376, w_026_155, w_014_559);
  nand2 I066_392(w_066_392, w_041_055, w_040_355);
  and2 I066_399(w_066_399, w_056_275, w_039_303);
  or2  I066_400(w_066_400, w_035_006, w_040_230);
  and2 I066_414(w_066_414, w_033_773, w_031_247);
  or2  I066_465(w_066_465, w_003_095, w_046_342);
  nand2 I066_475(w_066_475, w_050_086, w_044_043);
  or2  I066_476(w_066_476, w_037_164, w_044_278);
  or2  I066_485(w_066_485, w_061_216, w_019_070);
  and2 I066_493(w_066_493, w_041_079, w_016_002);
  and2 I066_511(w_066_511, w_009_052, w_061_221);
  nand2 I067_029(w_067_029, w_061_250, w_059_192);
  nand2 I067_075(w_067_075, w_049_358, w_049_210);
  nand2 I067_077(w_067_077, w_026_149, w_011_314);
  not1 I067_085(w_067_085, w_009_064);
  not1 I067_121(w_067_121, w_037_130);
  and2 I067_148(w_067_148, w_056_280, w_008_361);
  not1 I067_151(w_067_151, w_004_011);
  or2  I067_168(w_067_168, w_064_138, w_015_238);
  and2 I067_178(w_067_178, w_040_128, w_029_046);
  or2  I067_200(w_067_200, w_011_168, w_046_614);
  nand2 I067_216(w_067_216, w_061_394, w_020_044);
  nand2 I067_218(w_067_218, w_018_121, w_008_358);
  nand2 I067_224(w_067_224, w_059_317, w_004_009);
  and2 I067_226(w_067_226, w_061_023, w_018_101);
  and2 I067_229(w_067_229, w_001_385, w_029_054);
  or2  I067_242(w_067_242, w_015_099, w_029_084);
  and2 I067_245(w_067_245, w_027_791, w_001_231);
  not1 I067_251(w_067_251, w_001_866);
  and2 I067_263(w_067_263, w_040_103, w_028_709);
  nand2 I067_265(w_067_265, w_015_175, w_052_128);
  not1 I067_283(w_067_283, w_005_360);
  and2 I067_294(w_067_294, w_064_102, w_026_218);
  and2 I067_334(w_067_334, w_037_052, w_023_148);
  nand2 I067_343(w_067_343, w_020_124, w_016_471);
  nand2 I067_363(w_067_363, w_024_105, w_037_025);
  nand2 I067_444(w_067_444, w_017_003, w_048_448);
  or2  I067_508(w_067_508, w_026_408, w_038_640);
  or2  I067_516(w_067_516, w_052_133, w_042_002);
  or2  I067_615(w_067_615, w_045_179, w_024_042);
  or2  I067_649(w_067_649, w_010_148, w_000_402);
  not1 I067_711(w_067_711, w_049_018);
  or2  I067_724(w_067_724, w_034_583, w_016_495);
  and2 I067_728(w_067_728, w_008_271, w_050_141);
  not1 I067_746(w_067_746, w_019_084);
  not1 I067_754(w_067_754, w_034_431);
  not1 I067_785(w_067_785, w_038_046);
  nand2 I067_786(w_067_786, w_010_667, w_040_316);
  and2 I067_804(w_067_804, w_042_108, w_025_103);
  or2  I067_816(w_067_816, w_027_162, w_043_035);
  nand2 I067_866(w_067_866, w_047_281, w_008_222);
  not1 I067_880(w_067_880, w_030_230);
  nand2 I067_905(w_067_905, w_030_252, w_016_043);
  and2 I067_920(w_067_920, w_058_215, w_013_416);
  nand2 I067_921(w_067_921, w_019_085, w_065_665);
  and2 I067_939(w_067_939, w_056_311, w_064_750);
  not1 I067_945(w_067_945, w_055_664);
  nand2 I068_005(w_068_005, w_043_001, w_009_004);
  not1 I068_010(w_068_010, w_027_470);
  or2  I068_011(w_068_011, w_001_568, w_053_230);
  not1 I068_013(w_068_013, w_050_237);
  or2  I068_018(w_068_018, w_007_345, w_032_169);
  not1 I068_024(w_068_024, w_031_410);
  nand2 I068_025(w_068_025, w_038_562, w_047_385);
  nand2 I068_039(w_068_039, w_035_297, w_033_788);
  or2  I068_049(w_068_049, w_013_174, w_061_078);
  or2  I068_056(w_068_056, w_063_216, w_014_021);
  not1 I068_068(w_068_068, w_016_289);
  not1 I068_069(w_068_069, w_025_061);
  or2  I068_081(w_068_081, w_014_080, w_006_004);
  or2  I068_091(w_068_091, w_017_027, w_034_093);
  or2  I068_093(w_068_093, w_000_858, w_026_401);
  and2 I068_108(w_068_108, w_040_321, w_067_151);
  or2  I068_128(w_068_128, w_025_026, w_041_083);
  and2 I068_138(w_068_138, w_017_027, w_017_007);
  and2 I068_141(w_068_141, w_039_234, w_062_471);
  nand2 I068_145(w_068_145, w_041_082, w_036_145);
  nand2 I068_150(w_068_150, w_049_247, w_053_456);
  nand2 I068_157(w_068_157, w_047_178, w_067_251);
  not1 I068_171(w_068_171, w_013_253);
  nand2 I068_175(w_068_175, w_028_201, w_055_336);
  and2 I068_178(w_068_178, w_038_049, w_046_035);
  or2  I068_187(w_068_187, w_058_335, w_023_132);
  or2  I068_191(w_068_191, w_043_023, w_048_780);
  not1 I068_194(w_068_194, w_001_100);
  and2 I068_198(w_068_198, w_064_086, w_019_229);
  nand2 I068_203(w_068_203, w_037_026, w_026_272);
  and2 I068_212(w_068_212, w_046_669, w_018_107);
  and2 I068_219(w_068_219, w_002_361, w_014_426);
  or2  I068_234(w_068_234, w_007_515, w_024_080);
  or2  I068_256(w_068_256, w_027_602, w_056_275);
  nand2 I068_258(w_068_258, w_051_439, w_059_224);
  not1 I068_275(w_068_275, w_053_175);
  and2 I068_283(w_068_283, w_009_026, w_067_343);
  nand2 I068_302(w_068_302, w_009_025, w_005_496);
  or2  I068_303(w_068_303, w_050_195, w_019_051);
  and2 I068_306(w_068_306, w_046_300, w_014_341);
  nand2 I068_307(w_068_307, w_014_271, w_064_188);
  or2  I068_309(w_068_309, w_016_179, w_026_175);
  not1 I068_313(w_068_313, w_031_246);
  and2 I068_315(w_068_315, w_059_058, w_031_030);
  or2  I068_327(w_068_327, w_045_258, w_056_285);
  not1 I068_329(w_068_329, w_013_010);
  not1 I069_000(w_069_000, w_021_093);
  nand2 I069_004(w_069_004, w_061_241, w_066_023);
  nand2 I069_005(w_069_005, w_037_187, w_007_031);
  not1 I069_014(w_069_014, w_035_467);
  and2 I069_017(w_069_017, w_049_706, w_068_011);
  not1 I069_018(w_069_018, w_047_257);
  not1 I069_022(w_069_022, w_043_060);
  nand2 I069_024(w_069_024, w_004_013, w_060_212);
  and2 I069_029(w_069_029, w_045_382, w_034_801);
  not1 I069_033(w_069_033, w_000_682);
  not1 I069_058(w_069_058, w_041_052);
  nand2 I069_067(w_069_067, w_024_259, w_043_000);
  and2 I069_070(w_069_070, w_012_003, w_016_271);
  and2 I069_081(w_069_081, w_060_134, w_045_271);
  or2  I069_084(w_069_084, w_061_052, w_004_025);
  nand2 I069_107(w_069_107, w_028_180, w_009_068);
  nand2 I069_108(w_069_108, w_034_539, w_058_347);
  nand2 I069_114(w_069_114, w_023_455, w_055_548);
  not1 I069_125(w_069_125, w_059_090);
  and2 I069_126(w_069_126, w_000_533, w_006_053);
  not1 I069_137(w_069_137, w_017_007);
  or2  I069_139(w_069_139, w_065_509, w_051_308);
  nand2 I069_143(w_069_143, w_007_019, w_058_360);
  not1 I069_144(w_069_144, w_012_207);
  or2  I069_145(w_069_145, w_051_420, w_002_189);
  nand2 I069_146(w_069_146, w_038_050, w_010_622);
  nand2 I069_149(w_069_149, w_053_236, w_056_255);
  not1 I069_151(w_069_151, w_045_277);
  not1 I069_159(w_069_159, w_031_420);
  not1 I069_163(w_069_163, w_009_011);
  and2 I070_026(w_070_026, w_000_131, w_065_013);
  and2 I070_027(w_070_027, w_057_393, w_061_497);
  and2 I070_053(w_070_053, w_002_117, w_054_014);
  nand2 I070_117(w_070_117, w_011_241, w_035_072);
  or2  I070_147(w_070_147, w_059_247, w_053_388);
  or2  I070_154(w_070_154, w_016_273, w_007_189);
  nand2 I070_204(w_070_204, w_062_300, w_044_356);
  and2 I070_234(w_070_234, w_048_595, w_017_009);
  or2  I070_256(w_070_256, w_036_171, w_012_116);
  or2  I070_261(w_070_261, w_016_175, w_068_327);
  not1 I070_289(w_070_289, w_062_167);
  nand2 I070_346(w_070_346, w_000_542, w_065_091);
  not1 I070_356(w_070_356, w_010_065);
  nand2 I070_381(w_070_381, w_000_442, w_014_119);
  nand2 I070_388(w_070_388, w_039_162, w_036_201);
  and2 I070_403(w_070_403, w_034_775, w_026_031);
  nand2 I070_446(w_070_446, w_052_013, w_064_477);
  or2  I070_464(w_070_464, w_066_024, w_041_107);
  not1 I070_484(w_070_484, w_029_073);
  not1 I070_488(w_070_488, w_012_170);
  not1 I070_493(w_070_493, w_030_196);
  or2  I070_528(w_070_528, w_039_051, w_024_051);
  not1 I070_530(w_070_530, w_063_085);
  nand2 I070_551(w_070_551, w_044_181, w_053_492);
  not1 I070_552(w_070_552, w_033_257);
  and2 I070_595(w_070_595, w_049_587, w_044_055);
  or2  I070_629(w_070_629, w_035_121, w_052_031);
  nand2 I070_647(w_070_647, w_046_673, w_008_435);
  and2 I070_659(w_070_659, w_025_281, w_039_333);
  or2  I070_699(w_070_699, w_069_081, w_023_656);
  or2  I070_702(w_070_702, w_010_205, w_024_093);
  not1 I070_712(w_070_712, w_064_832);
  nand2 I070_730(w_070_730, w_060_189, w_041_009);
  not1 I070_748(w_070_748, w_031_035);
  nand2 I070_752(w_070_752, w_028_167, w_064_021);
  or2  I070_784(w_070_784, w_027_414, w_005_037);
  not1 I070_792(w_070_792, w_027_548);
  nand2 I070_823(w_070_823, w_043_022, w_049_069);
  nand2 I070_829(w_070_829, w_006_299, w_040_095);
  and2 I070_847(w_070_847, w_047_404, w_015_089);
  nand2 I070_864(w_070_864, w_048_679, w_035_041);
  or2  I070_888(w_070_888, w_036_105, w_017_006);
  not1 I070_915(w_070_915, w_044_036);
  and2 I070_926(w_070_926, w_000_617, w_028_092);
  not1 I070_935(w_070_935, w_041_089);
  nand2 I071_003(w_071_003, w_024_381, w_035_323);
  or2  I071_007(w_071_007, w_056_003, w_014_078);
  nand2 I071_011(w_071_011, w_002_224, w_022_453);
  or2  I071_016(w_071_016, w_054_147, w_006_287);
  and2 I071_040(w_071_040, w_007_338, w_016_297);
  and2 I071_041(w_071_041, w_061_235, w_020_022);
  and2 I071_046(w_071_046, w_067_866, w_039_340);
  not1 I071_057(w_071_057, w_029_011);
  and2 I071_058(w_071_058, w_022_400, w_011_295);
  not1 I071_060(w_071_060, w_045_123);
  nand2 I071_071(w_071_071, w_015_323, w_018_074);
  nand2 I071_076(w_071_076, w_056_196, w_059_282);
  and2 I071_079(w_071_079, w_016_345, w_042_024);
  or2  I071_095(w_071_095, w_022_524, w_011_233);
  nand2 I071_112(w_071_112, w_025_625, w_058_317);
  nand2 I071_115(w_071_115, w_026_014, w_064_537);
  not1 I071_116(w_071_116, w_027_757);
  not1 I071_125(w_071_125, w_066_051);
  or2  I071_129(w_071_129, w_052_071, w_047_006);
  or2  I071_134(w_071_134, w_044_043, w_042_031);
  not1 I071_137(w_071_137, w_069_145);
  not1 I071_147(w_071_147, w_006_017);
  not1 I071_151(w_071_151, w_037_140);
  and2 I071_158(w_071_158, w_051_165, w_025_473);
  or2  I071_166(w_071_166, w_070_234, w_054_134);
  and2 I071_174(w_071_174, w_030_473, w_051_118);
  and2 I071_206(w_071_206, w_060_012, w_014_179);
  nand2 I071_207(w_071_207, w_026_078, w_044_048);
  not1 I071_225(w_071_225, w_014_098);
  not1 I071_230(w_071_230, w_005_396);
  or2  I071_233(w_071_233, w_042_016, w_017_027);
  not1 I071_239(w_071_239, w_043_057);
  and2 I071_246(w_071_246, w_063_071, w_041_089);
  and2 I071_249(w_071_249, w_009_036, w_044_012);
  or2  I071_250(w_071_250, w_054_079, w_043_032);
  and2 I071_253(w_071_253, w_017_020, w_004_030);
  not1 I071_276(w_071_276, w_018_107);
  nand2 I071_281(w_071_281, w_065_613, w_030_418);
  not1 I071_284(w_071_284, w_003_206);
  not1 I071_286(w_071_286, w_024_339);
  or2  I071_306(w_071_306, w_002_359, w_024_297);
  not1 I071_312(w_071_312, w_065_006);
  nand2 I071_329(w_071_329, w_060_263, w_070_915);
  nand2 I071_337(w_071_337, w_019_102, w_033_407);
  and2 I071_351(w_071_351, w_033_007, w_067_921);
  not1 I071_363(w_071_363, w_063_260);
  and2 I071_366(w_071_366, w_048_525, w_018_176);
  nand2 I071_400(w_071_400, w_065_697, w_017_015);
  or2  I071_428(w_071_428, w_038_173, w_052_002);
  or2  I071_431(w_071_431, w_009_053, w_045_142);
  nand2 I071_434(w_071_434, w_047_460, w_068_093);
  or2  I071_436(w_071_436, w_009_028, w_000_129);
  nand2 I071_447(w_071_447, w_055_223, w_060_185);
  not1 I072_000(w_072_000, w_066_114);
  or2  I072_002(w_072_002, w_019_154, w_041_027);
  nand2 I072_003(w_072_003, w_029_211, w_024_083);
  or2  I072_004(w_072_004, w_036_276, w_062_029);
  and2 I072_006(w_072_006, w_046_673, w_015_101);
  and2 I072_007(w_072_007, w_042_077, w_023_154);
  not1 I072_008(w_072_008, w_012_249);
  and2 I072_010(w_072_010, w_059_068, w_030_399);
  nand2 I072_011(w_072_011, w_020_061, w_006_136);
  and2 I072_013(w_072_013, w_027_324, w_053_181);
  or2  I072_014(w_072_014, w_004_028, w_027_656);
  or2  I072_015(w_072_015, w_064_606, w_037_127);
  not1 I072_016(w_072_016, w_022_326);
  or2  I072_017(w_072_017, w_068_108, w_012_304);
  nand2 I072_019(w_072_019, w_003_074, w_024_446);
  not1 I072_020(w_072_020, w_005_404);
  nand2 I072_021(w_072_021, w_025_358, w_042_017);
  nand2 I072_022(w_072_022, w_034_096, w_033_358);
  not1 I072_023(w_072_023, w_071_134);
  nand2 I072_024(w_072_024, w_067_363, w_051_307);
  not1 I072_026(w_072_026, w_069_070);
  not1 I072_029(w_072_029, w_058_176);
  and2 I072_030(w_072_030, w_002_273, w_062_386);
  and2 I072_031(w_072_031, w_003_111, w_051_167);
  not1 I072_032(w_072_032, w_006_232);
  nand2 I072_033(w_072_033, w_041_015, w_032_523);
  or2  I072_034(w_072_034, w_070_926, w_068_307);
  nand2 I072_037(w_072_037, w_003_194, w_023_255);
  or2  I072_038(w_072_038, w_002_276, w_071_400);
  or2  I072_040(w_072_040, w_013_488, w_051_060);
  and2 I072_041(w_072_041, w_040_127, w_058_221);
  or2  I072_042(w_072_042, w_031_454, w_064_340);
  nand2 I072_046(w_072_046, w_024_391, w_016_429);
  or2  I072_048(w_072_048, w_003_016, w_003_044);
  or2  I072_049(w_072_049, w_011_062, w_065_850);
  nand2 I072_052(w_072_052, w_008_237, w_010_465);
  and2 I072_054(w_072_054, w_035_370, w_059_263);
  and2 I072_055(w_072_055, w_036_093, w_018_167);
  or2  I072_057(w_072_057, w_024_556, w_043_049);
  nand2 I072_060(w_072_060, w_059_277, w_035_286);
  or2  I072_063(w_072_063, w_030_424, w_034_534);
  and2 I072_065(w_072_065, w_053_012, w_023_059);
  or2  I072_067(w_072_067, w_000_180, w_030_210);
  or2  I073_005(w_073_005, w_068_302, w_059_193);
  or2  I073_012(w_073_012, w_021_184, w_036_113);
  or2  I073_021(w_073_021, w_071_076, w_044_142);
  not1 I073_030(w_073_030, w_050_038);
  or2  I073_034(w_073_034, w_050_248, w_002_005);
  nand2 I073_059(w_073_059, w_045_203, w_027_383);
  and2 I073_073(w_073_073, w_004_038, w_027_564);
  nand2 I073_090(w_073_090, w_003_032, w_037_147);
  nand2 I073_092(w_073_092, w_072_013, w_052_160);
  and2 I073_095(w_073_095, w_058_227, w_015_434);
  or2  I073_114(w_073_114, w_031_216, w_070_346);
  nand2 I073_117(w_073_117, w_063_290, w_010_161);
  and2 I073_123(w_073_123, w_042_004, w_028_535);
  nand2 I073_156(w_073_156, w_001_218, w_037_079);
  and2 I073_160(w_073_160, w_002_161, w_032_047);
  nand2 I073_214(w_073_214, w_059_308, w_049_930);
  not1 I073_292(w_073_292, w_012_165);
  or2  I073_322(w_073_322, w_021_149, w_048_114);
  and2 I073_323(w_073_323, w_053_760, w_028_424);
  not1 I073_331(w_073_331, w_029_041);
  and2 I073_339(w_073_339, w_025_678, w_072_037);
  and2 I073_409(w_073_409, w_053_109, w_007_245);
  not1 I073_411(w_073_411, w_015_207);
  or2  I073_413(w_073_413, w_052_049, w_055_474);
  or2  I073_416(w_073_416, w_014_311, w_013_350);
  not1 I073_430(w_073_430, w_045_505);
  not1 I073_452(w_073_452, w_038_012);
  nand2 I073_479(w_073_479, w_039_096, w_049_445);
  and2 I073_490(w_073_490, w_032_477, w_036_209);
  or2  I073_506(w_073_506, w_029_029, w_065_920);
  or2  I073_540(w_073_540, w_001_591, w_008_815);
  and2 I073_550(w_073_550, w_060_260, w_039_336);
  and2 I073_643(w_073_643, w_000_196, w_023_470);
  or2  I073_645(w_073_645, w_051_384, w_029_191);
  nand2 I073_655(w_073_655, w_045_092, w_053_081);
  not1 I073_663(w_073_663, w_004_031);
  nand2 I073_704(w_073_704, w_013_140, w_061_034);
  nand2 I073_705(w_073_705, w_071_071, w_036_237);
  and2 I073_747(w_073_747, w_012_287, w_062_022);
  nand2 I073_766(w_073_766, w_055_762, w_071_206);
  or2  I073_804(w_073_804, w_008_051, w_008_565);
  or2  I073_818(w_073_818, w_003_198, w_020_034);
  nand2 I074_003(w_074_003, w_024_247, w_064_554);
  nand2 I074_048(w_074_048, w_052_062, w_068_275);
  nand2 I074_061(w_074_061, w_046_185, w_050_002);
  and2 I074_067(w_074_067, w_051_071, w_027_095);
  and2 I074_156(w_074_156, w_054_167, w_028_125);
  not1 I074_214(w_074_214, w_030_160);
  nand2 I074_254(w_074_254, w_057_443, w_034_092);
  or2  I074_258(w_074_258, w_024_263, w_023_633);
  or2  I074_261(w_074_261, w_032_014, w_064_453);
  not1 I074_273(w_074_273, w_055_022);
  nand2 I074_294(w_074_294, w_011_140, w_008_510);
  and2 I074_297(w_074_297, w_072_026, w_041_047);
  nand2 I074_316(w_074_316, w_028_577, w_023_059);
  and2 I074_328(w_074_328, w_024_182, w_018_093);
  not1 I074_342(w_074_342, w_041_052);
  not1 I074_358(w_074_358, w_038_035);
  or2  I074_366(w_074_366, w_058_191, w_044_183);
  or2  I074_378(w_074_378, w_008_034, w_047_226);
  nand2 I074_383(w_074_383, w_033_384, w_033_074);
  not1 I074_463(w_074_463, w_055_033);
  or2  I074_467(w_074_467, w_030_217, w_024_549);
  or2  I074_479(w_074_479, w_012_359, w_025_595);
  nand2 I074_488(w_074_488, w_062_121, w_054_170);
  and2 I074_531(w_074_531, w_038_560, w_040_322);
  or2  I074_532(w_074_532, w_059_149, w_011_211);
  not1 I074_588(w_074_588, w_047_339);
  not1 I074_607(w_074_607, w_002_264);
  nand2 I074_633(w_074_633, w_042_077, w_071_147);
  nand2 I074_681(w_074_681, w_006_235, w_063_081);
  not1 I074_691(w_074_691, w_064_091);
  not1 I074_692(w_074_692, w_065_732);
  not1 I074_751(w_074_751, w_012_339);
  or2  I074_754(w_074_754, w_050_353, w_038_489);
  not1 I074_787(w_074_787, w_057_145);
  not1 I074_846(w_074_846, w_033_497);
  and2 I074_847(w_074_847, w_032_593, w_007_167);
  or2  I074_909(w_074_909, w_066_146, w_041_116);
  or2  I074_915(w_074_915, w_022_277, w_010_626);
  not1 I074_931(w_074_931, w_050_469);
  or2  I074_944(w_074_944, w_052_029, w_031_293);
  not1 I074_963(w_074_963, w_008_194);
  not1 I075_008(w_075_008, w_019_060);
  and2 I075_016(w_075_016, w_045_093, w_067_029);
  and2 I075_024(w_075_024, w_015_707, w_006_316);
  or2  I075_029(w_075_029, w_019_073, w_053_391);
  nand2 I075_036(w_075_036, w_019_413, w_048_068);
  and2 I075_043(w_075_043, w_059_135, w_015_180);
  not1 I075_051(w_075_051, w_003_169);
  and2 I075_052(w_075_052, w_051_286, w_048_139);
  and2 I075_069(w_075_069, w_046_157, w_066_202);
  or2  I075_082(w_075_082, w_056_279, w_064_727);
  and2 I075_089(w_075_089, w_020_029, w_015_316);
  and2 I075_100(w_075_100, w_006_078, w_071_312);
  not1 I075_101(w_075_101, w_060_185);
  or2  I075_103(w_075_103, w_054_077, w_015_734);
  not1 I075_108(w_075_108, w_032_498);
  and2 I075_111(w_075_111, w_003_193, w_005_199);
  not1 I075_114(w_075_114, w_026_003);
  and2 I075_144(w_075_144, w_027_678, w_054_080);
  nand2 I075_179(w_075_179, w_019_321, w_006_020);
  and2 I075_180(w_075_180, w_072_031, w_025_183);
  nand2 I075_188(w_075_188, w_018_048, w_045_443);
  nand2 I075_189(w_075_189, w_043_002, w_025_373);
  nand2 I075_192(w_075_192, w_042_013, w_069_004);
  nand2 I075_199(w_075_199, w_017_016, w_020_078);
  nand2 I075_229(w_075_229, w_033_909, w_040_105);
  or2  I075_258(w_075_258, w_028_509, w_040_272);
  not1 I075_260(w_075_260, w_028_777);
  or2  I075_284(w_075_284, w_064_036, w_007_332);
  not1 I075_285(w_075_285, w_050_376);
  or2  I076_006(w_076_006, w_029_092, w_059_278);
  and2 I076_008(w_076_008, w_008_051, w_069_163);
  nand2 I076_012(w_076_012, w_063_059, w_037_073);
  or2  I076_044(w_076_044, w_023_267, w_075_229);
  or2  I076_053(w_076_053, w_065_204, w_042_066);
  and2 I076_056(w_076_056, w_043_045, w_075_029);
  and2 I076_102(w_076_102, w_061_216, w_048_542);
  or2  I076_107(w_076_107, w_003_141, w_053_729);
  not1 I076_136(w_076_136, w_071_060);
  or2  I076_142(w_076_142, w_013_416, w_002_110);
  not1 I076_166(w_076_166, w_070_261);
  not1 I076_175(w_076_175, w_048_734);
  or2  I076_192(w_076_192, w_074_067, w_039_188);
  nand2 I076_220(w_076_220, w_069_108, w_053_300);
  not1 I076_227(w_076_227, w_028_404);
  nand2 I076_236(w_076_236, w_029_096, w_003_071);
  not1 I076_245(w_076_245, w_065_951);
  or2  I076_269(w_076_269, w_006_225, w_045_253);
  or2  I076_273(w_076_273, w_037_012, w_025_572);
  not1 I076_310(w_076_310, w_038_432);
  or2  I076_324(w_076_324, w_006_193, w_039_235);
  nand2 I076_330(w_076_330, w_048_368, w_012_134);
  nand2 I076_336(w_076_336, w_036_153, w_031_087);
  or2  I076_342(w_076_342, w_039_129, w_041_076);
  nand2 I076_352(w_076_352, w_006_002, w_066_107);
  and2 I076_356(w_076_356, w_021_024, w_061_168);
  not1 I076_360(w_076_360, w_032_064);
  nand2 I076_363(w_076_363, w_006_154, w_069_058);
  or2  I076_388(w_076_388, w_057_252, w_056_010);
  nand2 I076_393(w_076_393, w_057_041, w_037_148);
  not1 I076_417(w_076_417, w_056_275);
  or2  I076_422(w_076_422, w_068_258, w_014_324);
  or2  I076_433(w_076_433, w_009_050, w_040_083);
  and2 I076_437(w_076_437, w_065_951, w_065_950);
  or2  I076_449(w_076_449, w_017_003, w_006_036);
  and2 I076_582(w_076_582, w_064_503, w_052_117);
  not1 I076_591(w_076_591, w_056_170);
  or2  I076_616(w_076_616, w_040_102, w_037_114);
  and2 I076_617(w_076_617, w_035_612, w_008_061);
  not1 I077_012(w_077_012, w_040_252);
  nand2 I077_016(w_077_016, w_061_414, w_015_190);
  and2 I077_018(w_077_018, w_019_008, w_060_105);
  nand2 I077_028(w_077_028, w_066_359, w_012_361);
  and2 I077_041(w_077_041, w_065_711, w_023_228);
  and2 I077_047(w_077_047, w_036_199, w_044_261);
  or2  I077_069(w_077_069, w_002_289, w_044_063);
  or2  I077_074(w_077_074, w_060_297, w_073_092);
  not1 I077_083(w_077_083, w_025_177);
  and2 I077_098(w_077_098, w_001_731, w_063_027);
  and2 I077_100(w_077_100, w_022_259, w_010_531);
  not1 I077_101(w_077_101, w_027_141);
  nand2 I077_104(w_077_104, w_076_324, w_076_582);
  or2  I077_107(w_077_107, w_002_172, w_028_693);
  not1 I077_108(w_077_108, w_055_017);
  or2  I077_112(w_077_112, w_054_160, w_017_022);
  not1 I077_121(w_077_121, w_065_585);
  or2  I077_191(w_077_191, w_000_501, w_007_046);
  not1 I077_193(w_077_193, w_036_069);
  nand2 I077_194(w_077_194, w_039_461, w_048_189);
  and2 I077_197(w_077_197, w_062_037, w_046_067);
  nand2 I077_219(w_077_219, w_072_038, w_052_128);
  nand2 I077_240(w_077_240, w_070_488, w_074_003);
  nand2 I077_266(w_077_266, w_056_280, w_038_637);
  not1 I077_281(w_077_281, w_033_037);
  and2 I077_301(w_077_301, w_052_144, w_021_320);
  or2  I077_317(w_077_317, w_018_031, w_039_204);
  or2  I077_321(w_077_321, w_059_146, w_042_052);
  nand2 I077_323(w_077_323, w_038_303, w_059_235);
  nand2 I077_347(w_077_347, w_007_078, w_025_032);
  and2 I077_381(w_077_381, w_058_281, w_031_374);
  and2 I077_385(w_077_385, w_044_276, w_072_024);
  and2 I077_400(w_077_400, w_041_020, w_044_128);
  not1 I077_410(w_077_410, w_009_034);
  nand2 I077_419(w_077_419, w_046_627, w_024_556);
  not1 I077_430(w_077_430, w_036_105);
  not1 I077_443(w_077_443, w_026_023);
  and2 I077_449(w_077_449, w_051_392, w_064_574);
  or2  I077_472(w_077_472, w_026_055, w_017_007);
  nand2 I077_491(w_077_491, w_057_043, w_065_094);
  not1 I078_007(w_078_007, w_057_050);
  not1 I078_009(w_078_009, w_014_220);
  nand2 I078_017(w_078_017, w_069_108, w_060_178);
  or2  I078_020(w_078_020, w_066_017, w_005_137);
  not1 I078_028(w_078_028, w_022_169);
  or2  I078_034(w_078_034, w_013_171, w_035_307);
  nand2 I078_042(w_078_042, w_055_071, w_005_124);
  and2 I078_044(w_078_044, w_043_004, w_032_238);
  not1 I078_049(w_078_049, w_058_010);
  not1 I078_051(w_078_051, w_057_198);
  or2  I078_053(w_078_053, w_022_479, w_039_010);
  nand2 I078_055(w_078_055, w_062_253, w_068_069);
  not1 I078_073(w_078_073, w_033_739);
  not1 I078_077(w_078_077, w_040_003);
  and2 I078_087(w_078_087, w_003_084, w_050_323);
  not1 I078_090(w_078_090, w_039_395);
  not1 I078_102(w_078_102, w_005_375);
  or2  I078_121(w_078_121, w_049_341, w_009_000);
  or2  I078_132(w_078_132, w_004_016, w_020_050);
  not1 I078_151(w_078_151, w_035_588);
  and2 I078_161(w_078_161, w_008_252, w_025_145);
  nand2 I078_189(w_078_189, w_064_679, w_035_535);
  and2 I078_199(w_078_199, w_067_880, w_003_206);
  not1 I078_201(w_078_201, w_010_670);
  or2  I078_203(w_078_203, w_062_479, w_071_225);
  and2 I078_209(w_078_209, w_027_311, w_029_131);
  or2  I078_211(w_078_211, w_070_792, w_001_528);
  or2  I078_212(w_078_212, w_055_529, w_061_071);
  and2 I078_221(w_078_221, w_032_307, w_015_339);
  and2 I078_228(w_078_228, w_050_365, w_026_257);
  nand2 I078_233(w_078_233, w_029_151, w_040_110);
  nand2 I078_240(w_078_240, w_026_379, w_003_180);
  and2 I078_251(w_078_251, w_053_070, w_074_366);
  not1 I078_265(w_078_265, w_045_021);
  and2 I078_271(w_078_271, w_051_290, w_023_134);
  not1 I078_287(w_078_287, w_027_320);
  not1 I078_288(w_078_288, w_027_144);
  and2 I078_292(w_078_292, w_058_108, w_061_174);
  not1 I078_297(w_078_297, w_053_145);
  not1 I078_302(w_078_302, w_049_786);
  or2  I079_000(w_079_000, w_066_476, w_054_060);
  and2 I079_004(w_079_004, w_036_031, w_047_364);
  nand2 I079_015(w_079_015, w_023_427, w_015_324);
  nand2 I079_021(w_079_021, w_058_086, w_004_003);
  not1 I079_046(w_079_046, w_005_359);
  or2  I079_051(w_079_051, w_050_247, w_016_178);
  not1 I079_068(w_079_068, w_013_127);
  or2  I079_074(w_079_074, w_070_464, w_049_343);
  and2 I079_078(w_079_078, w_013_357, w_067_785);
  or2  I079_084(w_079_084, w_027_198, w_059_333);
  nand2 I079_086(w_079_086, w_051_342, w_014_584);
  nand2 I079_112(w_079_112, w_021_320, w_052_031);
  nand2 I079_114(w_079_114, w_058_199, w_013_479);
  and2 I079_121(w_079_121, w_065_251, w_069_005);
  not1 I079_129(w_079_129, w_062_373);
  not1 I079_130(w_079_130, w_070_864);
  and2 I079_136(w_079_136, w_003_152, w_001_340);
  not1 I079_146(w_079_146, w_021_244);
  and2 I079_150(w_079_150, w_065_051, w_074_328);
  and2 I079_162(w_079_162, w_056_188, w_060_301);
  nand2 I079_163(w_079_163, w_007_158, w_043_006);
  and2 I079_172(w_079_172, w_046_062, w_062_174);
  nand2 I079_182(w_079_182, w_053_364, w_039_047);
  nand2 I079_199(w_079_199, w_060_316, w_038_413);
  and2 I079_218(w_079_218, w_059_076, w_077_018);
  or2  I079_219(w_079_219, w_063_303, w_026_232);
  or2  I079_228(w_079_228, w_043_040, w_008_646);
  and2 I079_231(w_079_231, w_036_040, w_036_123);
  and2 I079_234(w_079_234, w_003_204, w_068_150);
  or2  I079_244(w_079_244, w_014_282, w_003_029);
  and2 I079_247(w_079_247, w_032_416, w_050_231);
  nand2 I080_008(w_080_008, w_036_009, w_010_109);
  or2  I080_009(w_080_009, w_004_014, w_038_186);
  nand2 I080_010(w_080_010, w_003_204, w_024_331);
  and2 I080_011(w_080_011, w_032_455, w_016_251);
  nand2 I080_016(w_080_016, w_050_186, w_073_506);
  not1 I080_022(w_080_022, w_014_323);
  nand2 I080_026(w_080_026, w_073_322, w_003_034);
  not1 I080_028(w_080_028, w_073_095);
  or2  I080_030(w_080_030, w_032_765, w_002_235);
  and2 I080_031(w_080_031, w_061_403, w_020_081);
  or2  I080_032(w_080_032, w_003_039, w_044_360);
  nand2 I080_038(w_080_038, w_007_039, w_044_047);
  or2  I080_043(w_080_043, w_072_049, w_052_132);
  and2 I080_046(w_080_046, w_031_243, w_010_304);
  nand2 I080_056(w_080_056, w_002_296, w_011_356);
  or2  I080_058(w_080_058, w_036_233, w_030_071);
  nand2 I080_059(w_080_059, w_023_528, w_001_268);
  not1 I080_061(w_080_061, w_045_151);
  not1 I080_063(w_080_063, w_076_449);
  or2  I080_064(w_080_064, w_064_741, w_048_198);
  nand2 I080_071(w_080_071, w_072_065, w_074_531);
  or2  I080_075(w_080_075, w_057_167, w_024_249);
  not1 I080_080(w_080_080, w_077_381);
  or2  I080_086(w_080_086, w_021_266, w_052_126);
  nand2 I080_092(w_080_092, w_020_036, w_025_552);
  nand2 I080_093(w_080_093, w_078_228, w_071_041);
  nand2 I080_099(w_080_099, w_023_143, w_058_196);
  or2  I080_102(w_080_102, w_001_522, w_074_931);
  and2 I080_103(w_080_103, w_023_161, w_002_454);
  not1 I080_104(w_080_104, w_070_629);
  and2 I080_107(w_080_107, w_041_050, w_074_358);
  and2 I080_108(w_080_108, w_052_051, w_071_249);
  nand2 I080_112(w_080_112, w_037_095, w_053_425);
  or2  I080_114(w_080_114, w_068_178, w_068_219);
  nand2 I081_016(w_081_016, w_064_692, w_045_323);
  not1 I081_017(w_081_017, w_036_205);
  or2  I081_026(w_081_026, w_014_545, w_061_298);
  and2 I081_041(w_081_041, w_048_068, w_070_356);
  not1 I081_060(w_081_060, w_056_219);
  or2  I081_083(w_081_083, w_078_233, w_010_760);
  or2  I081_084(w_081_084, w_022_225, w_053_292);
  or2  I081_090(w_081_090, w_048_606, w_038_117);
  not1 I081_119(w_081_119, w_063_130);
  and2 I081_122(w_081_122, w_027_671, w_036_019);
  and2 I081_134(w_081_134, w_013_450, w_015_128);
  and2 I081_139(w_081_139, w_034_414, w_018_191);
  or2  I081_170(w_081_170, w_004_020, w_046_148);
  not1 I081_212(w_081_212, w_025_163);
  not1 I081_237(w_081_237, w_058_151);
  not1 I081_240(w_081_240, w_069_029);
  nand2 I081_252(w_081_252, w_047_450, w_041_033);
  or2  I081_270(w_081_270, w_041_026, w_015_722);
  or2  I081_294(w_081_294, w_006_154, w_000_144);
  or2  I081_360(w_081_360, w_010_157, w_040_248);
  and2 I081_374(w_081_374, w_005_106, w_031_082);
  or2  I081_383(w_081_383, w_048_111, w_026_253);
  or2  I081_384(w_081_384, w_049_633, w_001_266);
  nand2 I081_458(w_081_458, w_041_112, w_034_210);
  and2 I081_478(w_081_478, w_007_314, w_063_322);
  or2  I081_527(w_081_527, w_007_221, w_043_036);
  not1 I081_538(w_081_538, w_009_030);
  not1 I081_563(w_081_563, w_004_035);
  or2  I081_567(w_081_567, w_041_084, w_051_002);
  and2 I081_582(w_081_582, w_053_002, w_009_001);
  not1 I081_590(w_081_590, w_053_058);
  and2 I082_004(w_082_004, w_020_054, w_021_107);
  nand2 I082_013(w_082_013, w_011_014, w_048_308);
  nand2 I082_015(w_082_015, w_014_071, w_030_038);
  not1 I082_027(w_082_027, w_080_108);
  and2 I082_028(w_082_028, w_054_196, w_054_185);
  nand2 I082_029(w_082_029, w_015_166, w_016_211);
  and2 I082_033(w_082_033, w_049_943, w_077_098);
  or2  I082_061(w_082_061, w_017_022, w_017_019);
  or2  I082_063(w_082_063, w_026_219, w_040_361);
  or2  I082_097(w_082_097, w_061_379, w_052_135);
  or2  I082_146(w_082_146, w_039_197, w_075_089);
  not1 I082_158(w_082_158, w_044_093);
  not1 I082_163(w_082_163, w_029_134);
  not1 I082_194(w_082_194, w_027_419);
  not1 I082_197(w_082_197, w_008_446);
  and2 I082_206(w_082_206, w_004_027, w_029_148);
  nand2 I082_212(w_082_212, w_072_063, w_040_272);
  and2 I082_217(w_082_217, w_061_286, w_051_255);
  nand2 I082_218(w_082_218, w_073_123, w_012_151);
  or2  I082_222(w_082_222, w_024_084, w_078_201);
  nand2 I082_228(w_082_228, w_024_511, w_053_346);
  or2  I082_231(w_082_231, w_081_119, w_010_771);
  nand2 I082_232(w_082_232, w_077_121, w_016_221);
  nand2 I082_240(w_082_240, w_063_231, w_003_090);
  nand2 I082_248(w_082_248, w_000_414, w_013_290);
  nand2 I082_253(w_082_253, w_032_308, w_039_187);
  or2  I082_257(w_082_257, w_066_187, w_059_123);
  or2  I082_258(w_082_258, w_011_272, w_048_620);
  not1 I082_266(w_082_266, w_068_171);
  nand2 I082_285(w_082_285, w_028_664, w_045_001);
  nand2 I082_301(w_082_301, w_020_100, w_076_393);
  nand2 I082_321(w_082_321, w_004_000, w_026_038);
  not1 I082_323(w_082_323, w_080_107);
  not1 I082_330(w_082_330, w_072_021);
  nand2 I082_334(w_082_334, w_068_256, w_031_045);
  or2  I082_342(w_082_342, w_051_381, w_064_131);
  or2  I082_344(w_082_344, w_041_019, w_072_052);
  and2 I083_000(w_083_000, w_049_936, w_035_258);
  or2  I083_021(w_083_021, w_028_630, w_059_145);
  not1 I083_022(w_083_022, w_057_202);
  and2 I083_023(w_083_023, w_014_270, w_028_109);
  and2 I083_030(w_083_030, w_061_377, w_009_022);
  nand2 I083_068(w_083_068, w_056_022, w_064_142);
  not1 I083_079(w_083_079, w_060_323);
  or2  I083_087(w_083_087, w_075_036, w_037_074);
  not1 I083_095(w_083_095, w_056_235);
  nand2 I083_109(w_083_109, w_074_532, w_009_065);
  and2 I083_111(w_083_111, w_064_515, w_050_407);
  not1 I083_137(w_083_137, w_014_451);
  or2  I083_138(w_083_138, w_070_552, w_055_163);
  and2 I083_147(w_083_147, w_026_075, w_024_037);
  not1 I083_153(w_083_153, w_079_004);
  nand2 I083_158(w_083_158, w_010_751, w_044_033);
  not1 I083_164(w_083_164, w_038_028);
  and2 I083_173(w_083_173, w_019_129, w_054_253);
  and2 I083_220(w_083_220, w_021_290, w_032_636);
  and2 I083_224(w_083_224, w_007_406, w_079_112);
  or2  I083_238(w_083_238, w_021_194, w_069_149);
  or2  I083_240(w_083_240, w_042_046, w_009_062);
  or2  I083_242(w_083_242, w_052_080, w_012_425);
  nand2 I083_249(w_083_249, w_029_136, w_082_218);
  or2  I083_253(w_083_253, w_048_575, w_065_883);
  not1 I083_259(w_083_259, w_067_263);
  and2 I083_266(w_083_266, w_041_078, w_011_246);
  and2 I083_274(w_083_274, w_053_515, w_079_146);
  nand2 I083_291(w_083_291, w_071_230, w_041_045);
  nand2 I083_302(w_083_302, w_059_142, w_065_914);
  or2  I083_310(w_083_310, w_010_034, w_027_522);
  and2 I083_435(w_083_435, w_072_007, w_051_066);
  not1 I083_439(w_083_439, w_050_386);
  nand2 I083_441(w_083_441, w_022_031, w_005_129);
  not1 I083_453(w_083_453, w_074_294);
  or2  I083_596(w_083_596, w_021_330, w_034_242);
  not1 I083_597(w_083_597, w_058_238);
  or2  I083_618(w_083_618, w_043_042, w_035_607);
  or2  I083_619(w_083_619, w_049_192, w_066_014);
  not1 I083_649(w_083_649, w_080_008);
  nand2 I083_651(w_083_651, w_013_035, w_025_281);
  or2  I083_653(w_083_653, w_000_743, w_010_008);
  or2  I084_012(w_084_012, w_012_030, w_016_057);
  and2 I084_029(w_084_029, w_009_063, w_063_103);
  and2 I084_033(w_084_033, w_014_634, w_031_135);
  and2 I084_035(w_084_035, w_060_101, w_034_266);
  or2  I084_039(w_084_039, w_047_183, w_065_433);
  and2 I084_050(w_084_050, w_067_444, w_037_090);
  not1 I084_062(w_084_062, w_021_024);
  nand2 I084_074(w_084_074, w_015_713, w_033_549);
  not1 I084_114(w_084_114, w_038_701);
  not1 I084_122(w_084_122, w_006_150);
  and2 I084_125(w_084_125, w_080_093, w_044_040);
  nand2 I084_128(w_084_128, w_079_199, w_082_158);
  or2  I084_131(w_084_131, w_010_088, w_057_253);
  nand2 I084_148(w_084_148, w_037_055, w_021_171);
  nand2 I084_169(w_084_169, w_072_037, w_069_107);
  nand2 I084_190(w_084_190, w_010_436, w_014_161);
  or2  I084_208(w_084_208, w_040_167, w_000_537);
  not1 I084_231(w_084_231, w_050_395);
  nand2 I084_234(w_084_234, w_030_184, w_070_403);
  and2 I084_240(w_084_240, w_043_044, w_047_472);
  or2  I084_257(w_084_257, w_045_214, w_077_100);
  or2  I084_268(w_084_268, w_021_337, w_062_031);
  not1 I084_294(w_084_294, w_034_154);
  or2  I084_299(w_084_299, w_002_482, w_046_501);
  not1 I084_329(w_084_329, w_075_069);
  or2  I084_428(w_084_428, w_043_051, w_054_089);
  nand2 I084_494(w_084_494, w_008_461, w_002_494);
  nand2 I084_526(w_084_526, w_058_064, w_047_107);
  and2 I084_535(w_084_535, w_044_304, w_021_313);
  nand2 I084_567(w_084_567, w_009_045, w_017_007);
  or2  I084_610(w_084_610, w_044_386, w_008_142);
  and2 I085_000(w_085_000, w_048_203, w_039_444);
  and2 I085_003(w_085_003, w_067_148, w_001_579);
  nand2 I085_004(w_085_004, w_048_748, w_070_026);
  and2 I085_006(w_085_006, w_048_458, w_081_237);
  and2 I085_008(w_085_008, w_052_041, w_083_173);
  nand2 I085_010(w_085_010, w_049_259, w_060_035);
  or2  I085_011(w_085_011, w_018_086, w_023_041);
  and2 I085_013(w_085_013, w_022_343, w_065_537);
  or2  I085_016(w_085_016, w_006_099, w_061_461);
  nand2 I085_017(w_085_017, w_061_502, w_073_416);
  or2  I085_019(w_085_019, w_031_031, w_055_001);
  nand2 I085_020(w_085_020, w_059_138, w_035_150);
  nand2 I085_021(w_085_021, w_029_157, w_012_126);
  nand2 I085_022(w_085_022, w_046_504, w_064_690);
  not1 I085_023(w_085_023, w_034_043);
  and2 I085_024(w_085_024, w_022_268, w_015_600);
  not1 I085_026(w_085_026, w_032_146);
  not1 I085_027(w_085_027, w_006_304);
  not1 I085_037(w_085_037, w_049_245);
  or2  I085_039(w_085_039, w_010_323, w_046_184);
  nand2 I085_041(w_085_041, w_048_412, w_081_294);
  not1 I085_043(w_085_043, w_031_017);
  not1 I085_044(w_085_044, w_036_283);
  not1 I085_050(w_085_050, w_048_118);
  and2 I085_051(w_085_051, w_041_019, w_070_752);
  not1 I085_054(w_085_054, w_078_090);
  and2 I085_055(w_085_055, w_064_749, w_030_133);
  and2 I085_056(w_085_056, w_027_624, w_056_007);
  and2 I085_057(w_085_057, w_025_100, w_042_056);
  and2 I085_058(w_085_058, w_083_224, w_049_913);
  and2 I085_059(w_085_059, w_035_191, w_024_394);
  or2  I085_060(w_085_060, w_073_430, w_050_038);
  not1 I085_070(w_085_070, w_077_101);
  not1 I085_071(w_085_071, w_057_031);
  or2  I086_001(w_086_001, w_073_704, w_005_118);
  or2  I086_006(w_086_006, w_082_231, w_016_206);
  or2  I086_012(w_086_012, w_056_012, w_062_228);
  or2  I086_017(w_086_017, w_082_063, w_022_276);
  not1 I086_026(w_086_026, w_034_579);
  nand2 I086_059(w_086_059, w_059_151, w_000_217);
  nand2 I086_060(w_086_060, w_003_206, w_019_363);
  and2 I086_077(w_086_077, w_041_085, w_020_017);
  not1 I086_090(w_086_090, w_009_042);
  and2 I086_099(w_086_099, w_067_786, w_073_021);
  nand2 I086_106(w_086_106, w_046_479, w_084_567);
  and2 I086_116(w_086_116, w_025_126, w_057_305);
  and2 I086_143(w_086_143, w_033_011, w_008_077);
  nand2 I086_167(w_086_167, w_001_867, w_023_108);
  and2 I086_182(w_086_182, w_013_274, w_023_326);
  and2 I086_202(w_086_202, w_041_000, w_046_181);
  nand2 I086_215(w_086_215, w_064_637, w_021_264);
  nand2 I086_222(w_086_222, w_055_723, w_018_062);
  not1 I086_242(w_086_242, w_057_323);
  nand2 I086_358(w_086_358, w_009_034, w_036_005);
  or2  I086_364(w_086_364, w_064_338, w_061_298);
  nand2 I086_395(w_086_395, w_052_153, w_076_220);
  not1 I086_408(w_086_408, w_006_259);
  and2 I086_415(w_086_415, w_063_119, w_032_107);
  nand2 I086_427(w_086_427, w_076_342, w_072_023);
  or2  I086_428(w_086_428, w_073_804, w_042_110);
  or2  I086_482(w_086_482, w_060_305, w_045_227);
  nand2 I086_577(w_086_577, w_030_281, w_050_059);
  nand2 I086_590(w_086_590, w_082_146, w_062_251);
  and2 I086_596(w_086_596, w_065_423, w_019_342);
  nand2 I086_642(w_086_642, w_043_031, w_002_087);
  or2  I086_652(w_086_652, w_002_273, w_034_554);
  nand2 I086_659(w_086_659, w_013_333, w_051_204);
  and2 I086_666(w_086_666, w_058_302, w_045_013);
  or2  I086_668(w_086_668, w_065_861, w_083_240);
  or2  I086_701(w_086_701, w_034_063, w_020_007);
  and2 I086_705(w_086_705, w_058_002, w_085_023);
  not1 I086_709(w_086_709, w_028_067);
  and2 I086_720(w_086_720, w_054_054, w_022_020);
  not1 I086_721(w_086_721, w_041_114);
  not1 I086_725(w_086_725, w_045_549);
  nand2 I086_745(w_086_745, w_052_036, w_050_401);
  nand2 I086_750(w_086_750, w_041_052, w_052_009);
  or2  I086_776(w_086_776, w_010_236, w_022_482);
  nand2 I087_024(w_087_024, w_019_300, w_036_278);
  not1 I087_039(w_087_039, w_002_158);
  or2  I087_040(w_087_040, w_076_053, w_001_770);
  or2  I087_044(w_087_044, w_037_112, w_020_024);
  and2 I087_049(w_087_049, w_061_033, w_031_016);
  or2  I087_052(w_087_052, w_044_007, w_062_314);
  or2  I087_053(w_087_053, w_042_033, w_058_154);
  nand2 I087_059(w_087_059, w_028_368, w_073_160);
  or2  I087_069(w_087_069, w_030_483, w_048_694);
  and2 I087_080(w_087_080, w_067_218, w_085_059);
  not1 I087_109(w_087_109, w_086_077);
  and2 I087_135(w_087_135, w_007_001, w_018_068);
  or2  I087_144(w_087_144, w_017_019, w_049_690);
  or2  I087_145(w_087_145, w_078_251, w_086_415);
  or2  I087_147(w_087_147, w_035_265, w_057_002);
  and2 I087_177(w_087_177, w_045_474, w_069_014);
  and2 I087_195(w_087_195, w_063_217, w_061_560);
  and2 I087_220(w_087_220, w_029_111, w_065_017);
  not1 I087_226(w_087_226, w_050_152);
  and2 I087_256(w_087_256, w_038_123, w_008_387);
  or2  I087_263(w_087_263, w_035_527, w_053_592);
  and2 I087_304(w_087_304, w_013_297, w_064_806);
  or2  I087_313(w_087_313, w_045_153, w_051_134);
  or2  I087_329(w_087_329, w_066_485, w_085_013);
  or2  I087_348(w_087_348, w_050_282, w_016_181);
  or2  I088_030(w_088_030, w_063_242, w_039_103);
  nand2 I088_037(w_088_037, w_087_256, w_070_712);
  nand2 I088_063(w_088_063, w_080_059, w_019_128);
  or2  I088_077(w_088_077, w_009_049, w_073_012);
  or2  I088_098(w_088_098, w_067_905, w_072_000);
  not1 I088_108(w_088_108, w_073_030);
  and2 I088_151(w_088_151, w_000_886, w_073_766);
  or2  I088_163(w_088_163, w_013_328, w_086_721);
  or2  I088_179(w_088_179, w_065_972, w_043_035);
  or2  I088_189(w_088_189, w_010_269, w_016_146);
  not1 I088_193(w_088_193, w_065_312);
  not1 I088_207(w_088_207, w_008_211);
  not1 I088_214(w_088_214, w_086_143);
  nand2 I088_230(w_088_230, w_012_063, w_015_348);
  or2  I088_285(w_088_285, w_053_019, w_017_003);
  nand2 I088_379(w_088_379, w_086_720, w_053_437);
  not1 I088_404(w_088_404, w_001_380);
  not1 I088_458(w_088_458, w_044_223);
  and2 I088_500(w_088_500, w_025_014, w_024_014);
  nand2 I088_533(w_088_533, w_006_095, w_019_402);
  nand2 I088_534(w_088_534, w_011_162, w_034_681);
  and2 I088_618(w_088_618, w_086_659, w_016_036);
  or2  I088_619(w_088_619, w_005_159, w_054_141);
  or2  I088_655(w_088_655, w_013_251, w_002_069);
  or2  I088_695(w_088_695, w_067_508, w_001_047);
  and2 I089_006(w_089_006, w_084_074, w_021_093);
  not1 I089_009(w_089_009, w_022_414);
  not1 I089_015(w_089_015, w_029_113);
  and2 I089_018(w_089_018, w_021_219, w_057_325);
  not1 I089_019(w_089_019, w_052_129);
  and2 I089_022(w_089_022, w_016_172, w_081_139);
  nand2 I089_024(w_089_024, w_011_247, w_012_419);
  not1 I089_031(w_089_031, w_041_054);
  not1 I089_056(w_089_056, w_049_194);
  and2 I089_068(w_089_068, w_044_194, w_027_307);
  or2  I089_074(w_089_074, w_051_517, w_044_155);
  nand2 I089_078(w_089_078, w_075_051, w_074_846);
  not1 I089_079(w_089_079, w_034_567);
  not1 I089_082(w_089_082, w_083_597);
  not1 I089_088(w_089_088, w_061_055);
  and2 I089_090(w_089_090, w_007_266, w_057_425);
  and2 I089_091(w_089_091, w_074_633, w_001_101);
  or2  I089_095(w_089_095, w_044_184, w_081_567);
  or2  I089_098(w_089_098, w_059_213, w_023_403);
  and2 I089_107(w_089_107, w_021_230, w_038_057);
  and2 I089_113(w_089_113, w_087_059, w_065_223);
  nand2 I089_127(w_089_127, w_056_010, w_003_215);
  and2 I089_135(w_089_135, w_081_252, w_032_237);
  or2  I090_003(w_090_003, w_046_467, w_014_325);
  and2 I090_019(w_090_019, w_039_036, w_036_046);
  or2  I090_026(w_090_026, w_089_015, w_036_271);
  and2 I090_038(w_090_038, w_038_047, w_084_148);
  nand2 I090_048(w_090_048, w_042_067, w_014_524);
  not1 I090_066(w_090_066, w_039_005);
  not1 I090_079(w_090_079, w_002_022);
  or2  I090_086(w_090_086, w_081_060, w_000_212);
  not1 I090_121(w_090_121, w_056_236);
  not1 I090_127(w_090_127, w_084_128);
  not1 I090_139(w_090_139, w_039_228);
  nand2 I090_160(w_090_160, w_050_396, w_033_692);
  nand2 I090_200(w_090_200, w_085_037, w_002_489);
  or2  I090_205(w_090_205, w_012_106, w_031_171);
  nand2 I090_209(w_090_209, w_029_207, w_035_135);
  and2 I090_212(w_090_212, w_087_348, w_086_143);
  not1 I090_220(w_090_220, w_075_179);
  not1 I090_224(w_090_224, w_071_046);
  and2 I090_238(w_090_238, w_043_047, w_069_114);
  not1 I090_244(w_090_244, w_045_053);
  or2  I090_250(w_090_250, w_066_493, w_081_122);
  not1 I090_252(w_090_252, w_031_246);
  and2 I090_268(w_090_268, w_077_400, w_080_092);
  or2  I090_270(w_090_270, w_012_275, w_018_074);
  nand2 I090_271(w_090_271, w_088_655, w_002_471);
  and2 I090_281(w_090_281, w_012_138, w_013_126);
  not1 I090_283(w_090_283, w_022_353);
  or2  I090_295(w_090_295, w_024_557, w_049_321);
  or2  I090_297(w_090_297, w_025_060, w_024_079);
  and2 I090_328(w_090_328, w_026_028, w_019_077);
  and2 I090_332(w_090_332, w_026_089, w_063_037);
  nand2 I090_335(w_090_335, w_081_084, w_084_125);
  or2  I090_336(w_090_336, w_027_067, w_058_320);
  not1 I090_337(w_090_337, w_084_039);
  nand2 I090_384(w_090_384, w_085_008, w_061_222);
  not1 I090_393(w_090_393, w_033_437);
  nand2 I091_000(w_091_000, w_065_895, w_035_563);
  not1 I091_002(w_091_002, w_049_521);
  not1 I091_031(w_091_031, w_032_603);
  nand2 I091_036(w_091_036, w_080_043, w_014_248);
  or2  I091_048(w_091_048, w_075_260, w_059_214);
  not1 I091_068(w_091_068, w_018_177);
  and2 I091_082(w_091_082, w_013_478, w_052_016);
  and2 I091_125(w_091_125, w_053_341, w_030_177);
  or2  I091_127(w_091_127, w_017_023, w_017_003);
  and2 I091_145(w_091_145, w_007_168, w_064_002);
  and2 I091_150(w_091_150, w_024_357, w_078_265);
  nand2 I091_170(w_091_170, w_016_371, w_024_072);
  and2 I091_173(w_091_173, w_070_935, w_074_061);
  nand2 I091_179(w_091_179, w_046_689, w_043_011);
  nand2 I091_182(w_091_182, w_058_197, w_019_243);
  or2  I091_186(w_091_186, w_072_004, w_058_065);
  and2 I091_190(w_091_190, w_039_175, w_048_313);
  nand2 I091_206(w_091_206, w_064_311, w_081_527);
  nand2 I091_214(w_091_214, w_061_147, w_078_292);
  and2 I091_232(w_091_232, w_042_004, w_070_595);
  or2  I091_233(w_091_233, w_030_012, w_078_007);
  and2 I091_279(w_091_279, w_010_208, w_023_240);
  or2  I091_316(w_091_316, w_047_226, w_056_212);
  and2 I091_347(w_091_347, w_014_058, w_088_533);
  or2  I091_403(w_091_403, w_063_293, w_039_268);
  and2 I091_408(w_091_408, w_017_016, w_000_416);
  nand2 I091_507(w_091_507, w_062_474, w_028_739);
  nand2 I091_552(w_091_552, w_088_193, w_050_035);
  or2  I091_555(w_091_555, w_047_464, w_085_019);
  not1 I092_011(w_092_011, w_006_287);
  nand2 I092_033(w_092_033, w_040_140, w_024_008);
  or2  I092_034(w_092_034, w_001_696, w_032_383);
  not1 I092_037(w_092_037, w_021_328);
  and2 I092_038(w_092_038, w_003_041, w_004_011);
  nand2 I092_043(w_092_043, w_043_064, w_014_345);
  nand2 I092_083(w_092_083, w_049_886, w_031_324);
  or2  I092_092(w_092_092, w_018_056, w_040_340);
  not1 I092_122(w_092_122, w_043_011);
  nand2 I092_129(w_092_129, w_023_058, w_056_166);
  or2  I092_130(w_092_130, w_021_198, w_002_488);
  not1 I092_138(w_092_138, w_090_384);
  or2  I092_210(w_092_210, w_073_818, w_015_019);
  or2  I092_239(w_092_239, w_065_333, w_002_047);
  nand2 I092_282(w_092_282, w_021_083, w_066_317);
  or2  I092_461(w_092_461, w_065_652, w_028_890);
  or2  I092_503(w_092_503, w_042_074, w_086_668);
  or2  I092_524(w_092_524, w_073_073, w_050_003);
  or2  I092_546(w_092_546, w_024_094, w_085_004);
  and2 I092_644(w_092_644, w_066_376, w_049_334);
  not1 I092_680(w_092_680, w_052_034);
  or2  I092_706(w_092_706, w_050_039, w_048_158);
  and2 I092_747(w_092_747, w_041_010, w_049_307);
  and2 I093_015(w_093_015, w_033_254, w_029_094);
  nand2 I093_107(w_093_107, w_091_031, w_063_138);
  and2 I093_111(w_093_111, w_011_009, w_040_156);
  or2  I093_130(w_093_130, w_057_262, w_086_167);
  not1 I093_137(w_093_137, w_056_231);
  nand2 I093_169(w_093_169, w_032_095, w_001_418);
  or2  I093_200(w_093_200, w_036_166, w_068_138);
  nand2 I093_203(w_093_203, w_072_008, w_059_147);
  or2  I093_227(w_093_227, w_032_100, w_069_033);
  or2  I093_241(w_093_241, w_020_074, w_001_491);
  not1 I093_258(w_093_258, w_046_185);
  not1 I093_279(w_093_279, w_079_074);
  nand2 I093_320(w_093_320, w_057_017, w_050_229);
  nand2 I093_346(w_093_346, w_062_140, w_089_098);
  not1 I093_353(w_093_353, w_034_103);
  and2 I093_374(w_093_374, w_010_147, w_033_045);
  or2  I093_423(w_093_423, w_041_119, w_065_279);
  and2 I093_484(w_093_484, w_013_389, w_053_824);
  nand2 I093_600(w_093_600, w_086_182, w_026_390);
  and2 I093_720(w_093_720, w_090_335, w_085_021);
  or2  I093_734(w_093_734, w_031_314, w_076_107);
  not1 I093_769(w_093_769, w_012_446);
  or2  I093_791(w_093_791, w_067_816, w_023_604);
  not1 I093_825(w_093_825, w_024_200);
  nand2 I093_858(w_093_858, w_058_070, w_058_155);
  not1 I093_878(w_093_878, w_006_315);
  or2  I093_911(w_093_911, w_028_625, w_073_117);
  not1 I093_915(w_093_915, w_044_199);
  and2 I093_919(w_093_919, w_082_266, w_027_040);
  nand2 I094_011(w_094_011, w_088_037, w_056_177);
  not1 I094_028(w_094_028, w_047_492);
  or2  I094_055(w_094_055, w_072_041, w_033_053);
  not1 I094_078(w_094_078, w_006_292);
  or2  I094_113(w_094_113, w_026_217, w_053_151);
  or2  I094_115(w_094_115, w_023_012, w_082_212);
  nand2 I094_124(w_094_124, w_029_031, w_025_576);
  nand2 I094_134(w_094_134, w_023_522, w_033_467);
  and2 I094_150(w_094_150, w_043_018, w_068_203);
  nand2 I094_169(w_094_169, w_054_016, w_012_138);
  nand2 I094_208(w_094_208, w_003_120, w_093_346);
  and2 I094_217(w_094_217, w_002_406, w_087_220);
  and2 I094_292(w_094_292, w_068_194, w_025_171);
  nand2 I094_313(w_094_313, w_071_166, w_004_020);
  not1 I094_415(w_094_415, w_063_274);
  or2  I094_506(w_094_506, w_021_172, w_022_391);
  or2  I094_671(w_094_671, w_060_249, w_081_458);
  not1 I094_710(w_094_710, w_086_026);
  and2 I094_726(w_094_726, w_058_058, w_093_203);
  nand2 I094_763(w_094_763, w_085_020, w_082_013);
  nand2 I094_781(w_094_781, w_042_043, w_008_002);
  not1 I094_794(w_094_794, w_063_210);
  and2 I094_817(w_094_817, w_008_485, w_011_407);
  nand2 I094_869(w_094_869, w_061_255, w_039_089);
  and2 I094_884(w_094_884, w_037_130, w_086_745);
  and2 I095_000(w_095_000, w_003_161, w_039_049);
  or2  I095_002(w_095_002, w_012_242, w_069_151);
  nand2 I095_008(w_095_008, w_027_400, w_063_099);
  not1 I095_009(w_095_009, w_034_250);
  or2  I095_017(w_095_017, w_069_024, w_078_240);
  or2  I095_019(w_095_019, w_024_051, w_094_124);
  nand2 I095_022(w_095_022, w_028_216, w_077_194);
  nand2 I095_028(w_095_028, w_013_099, w_039_443);
  nand2 I095_030(w_095_030, w_043_039, w_042_084);
  not1 I095_040(w_095_040, w_038_573);
  and2 I095_054(w_095_054, w_050_166, w_065_373);
  nand2 I095_074(w_095_074, w_016_215, w_004_028);
  nand2 I095_081(w_095_081, w_034_089, w_002_249);
  nand2 I095_094(w_095_094, w_071_151, w_055_611);
  and2 I095_101(w_095_101, w_048_090, w_084_190);
  or2  I095_108(w_095_108, w_042_074, w_040_186);
  and2 I095_112(w_095_112, w_046_674, w_075_108);
  and2 I095_115(w_095_115, w_033_454, w_032_732);
  not1 I095_128(w_095_128, w_013_355);
  not1 I095_131(w_095_131, w_009_049);
  and2 I095_149(w_095_149, w_084_169, w_036_193);
  or2  I095_150(w_095_150, w_044_140, w_090_297);
  not1 I095_153(w_095_153, w_051_047);
  or2  I095_163(w_095_163, w_019_242, w_010_391);
  nand2 I095_164(w_095_164, w_065_422, w_078_199);
  not1 I095_165(w_095_165, w_065_978);
  nand2 I095_181(w_095_181, w_006_305, w_040_308);
  and2 I095_182(w_095_182, w_079_228, w_016_099);
  nand2 I096_028(w_096_028, w_058_080, w_044_343);
  or2  I096_075(w_096_075, w_094_313, w_052_082);
  not1 I096_086(w_096_086, w_078_020);
  or2  I096_097(w_096_097, w_000_786, w_074_909);
  not1 I096_100(w_096_100, w_068_275);
  not1 I096_108(w_096_108, w_017_015);
  not1 I096_114(w_096_114, w_091_068);
  and2 I096_118(w_096_118, w_054_195, w_079_150);
  and2 I096_120(w_096_120, w_049_742, w_089_082);
  nand2 I096_124(w_096_124, w_013_086, w_046_660);
  not1 I096_130(w_096_130, w_081_083);
  or2  I096_131(w_096_131, w_031_095, w_016_320);
  not1 I096_139(w_096_139, w_010_623);
  nand2 I096_160(w_096_160, w_034_573, w_076_582);
  not1 I096_168(w_096_168, w_093_769);
  nand2 I096_185(w_096_185, w_030_216, w_033_610);
  or2  I096_218(w_096_218, w_057_113, w_021_088);
  and2 I096_229(w_096_229, w_039_008, w_040_298);
  or2  I096_248(w_096_248, w_015_445, w_094_869);
  nand2 I096_254(w_096_254, w_063_146, w_068_187);
  nand2 I096_255(w_096_255, w_041_114, w_093_015);
  and2 I096_293(w_096_293, w_075_008, w_028_729);
  or2  I096_299(w_096_299, w_080_112, w_014_091);
  nand2 I096_346(w_096_346, w_011_041, w_050_200);
  not1 I096_348(w_096_348, w_053_616);
  not1 I096_380(w_096_380, w_094_169);
  nand2 I096_381(w_096_381, w_066_399, w_044_231);
  not1 I096_419(w_096_419, w_019_314);
  or2  I096_475(w_096_475, w_045_662, w_076_336);
  or2  I096_566(w_096_566, w_066_115, w_033_675);
  nand2 I096_581(w_096_581, w_016_112, w_044_391);
  nand2 I096_627(w_096_629, w_010_492, w_096_628);
  and2 I096_628(w_096_630, w_096_629, w_003_107);
  and2 I096_629(w_096_631, w_096_630, w_096_653);
  nand2 I096_630(w_096_632, w_096_631, w_014_474);
  and2 I096_631(w_096_633, w_043_028, w_096_632);
  nand2 I096_632(w_096_634, w_093_600, w_096_633);
  or2  I096_633(w_096_635, w_096_634, w_051_123);
  and2 I096_634(w_096_636, w_082_323, w_096_635);
  nand2 I096_635(w_096_637, w_086_060, w_096_636);
  not1 I096_636(w_096_638, w_096_637);
  and2 I096_637(w_096_628, w_096_638, w_025_532);
  or2  I096_638(w_096_643, w_096_642, w_005_259);
  not1 I096_639(w_096_644, w_096_643);
  and2 I096_640(w_096_645, w_017_011, w_096_644);
  or2  I096_641(w_096_646, w_020_013, w_096_645);
  not1 I096_642(w_096_647, w_096_646);
  nand2 I096_643(w_096_648, w_096_647, w_075_189);
  nand2 I096_644(w_096_649, w_096_648, w_026_309);
  not1 I096_645(w_096_650, w_096_649);
  nand2 I096_646(w_096_651, w_046_539, w_096_650);
  not1 I096_647(w_096_642, w_096_631);
  and2 I096_648(w_096_653, w_084_131, w_096_651);
  not1 I097_001(w_097_001, w_045_348);
  not1 I097_030(w_097_030, w_091_048);
  or2  I097_038(w_097_038, w_062_069, w_096_419);
  not1 I097_041(w_097_041, w_031_002);
  not1 I097_045(w_097_045, w_071_281);
  nand2 I097_054(w_097_054, w_088_230, w_089_018);
  and2 I097_057(w_097_057, w_037_141, w_034_206);
  or2  I097_058(w_097_058, w_064_169, w_034_344);
  not1 I097_069(w_097_069, w_096_108);
  nand2 I097_073(w_097_073, w_018_126, w_059_032);
  nand2 I097_077(w_097_077, w_068_198, w_081_478);
  nand2 I097_141(w_097_141, w_015_135, w_006_123);
  nand2 I097_171(w_097_171, w_055_603, w_064_526);
  or2  I097_183(w_097_183, w_034_088, w_063_193);
  nand2 I097_192(w_097_192, w_079_084, w_073_655);
  not1 I097_228(w_097_228, w_044_036);
  nand2 I097_231(w_097_231, w_090_281, w_010_501);
  or2  I097_260(w_097_260, w_002_322, w_078_049);
  or2  I097_329(w_097_329, w_071_246, w_018_150);
  not1 I097_441(w_097_441, w_034_034);
  or2  I097_495(w_097_495, w_001_072, w_027_324);
  not1 I097_501(w_097_501, w_019_215);
  nand2 I097_502(w_097_502, w_046_540, w_055_731);
  nand2 I097_513(w_097_513, w_000_572, w_088_379);
  or2  I097_583(w_097_583, w_082_027, w_003_169);
  not1 I097_595(w_097_595, w_086_001);
  or2  I097_602(w_097_602, w_056_081, w_000_783);
  and2 I097_634(w_097_634, w_010_033, w_063_038);
  nand2 I097_636(w_097_636, w_056_227, w_026_174);
  not1 I098_025(w_098_025, w_072_023);
  or2  I098_035(w_098_035, w_025_348, w_002_015);
  nand2 I098_036(w_098_036, w_093_111, w_054_160);
  not1 I098_048(w_098_048, w_060_247);
  nand2 I098_079(w_098_079, w_014_307, w_018_091);
  or2  I098_095(w_098_095, w_000_916, w_013_079);
  not1 I098_189(w_098_189, w_049_397);
  nand2 I098_222(w_098_222, w_003_047, w_053_310);
  nand2 I098_231(w_098_231, w_036_132, w_004_022);
  or2  I098_257(w_098_257, w_072_048, w_069_114);
  and2 I098_278(w_098_278, w_089_056, w_047_396);
  and2 I098_310(w_098_310, w_050_371, w_048_591);
  nand2 I098_315(w_098_315, w_025_158, w_086_364);
  not1 I098_329(w_098_329, w_083_079);
  and2 I098_341(w_098_341, w_037_152, w_008_187);
  not1 I098_410(w_098_410, w_039_417);
  not1 I098_422(w_098_422, w_070_530);
  and2 I098_450(w_098_450, w_028_289, w_063_135);
  and2 I098_451(w_098_451, w_054_112, w_020_012);
  not1 I098_465(w_098_465, w_020_100);
  or2  I099_006(w_099_006, w_071_079, w_069_022);
  and2 I099_020(w_099_020, w_004_015, w_025_208);
  and2 I099_035(w_099_035, w_021_037, w_027_619);
  and2 I099_036(w_099_036, w_070_528, w_073_479);
  and2 I099_038(w_099_038, w_050_198, w_020_063);
  not1 I099_059(w_099_059, w_060_331);
  not1 I099_070(w_099_070, w_041_075);
  nand2 I099_077(w_099_077, w_097_054, w_010_531);
  or2  I099_082(w_099_082, w_060_307, w_041_073);
  not1 I099_085(w_099_085, w_018_026);
  not1 I099_102(w_099_102, w_015_047);
  or2  I099_105(w_099_105, w_052_143, w_071_040);
  not1 I099_114(w_099_114, w_084_231);
  not1 I099_120(w_099_120, w_049_925);
  or2  I099_128(w_099_128, w_006_232, w_081_563);
  nand2 I099_130(w_099_130, w_095_108, w_057_023);
  and2 I099_157(w_099_157, w_040_071, w_077_104);
  nand2 I099_158(w_099_158, w_023_040, w_016_474);
  not1 I099_171(w_099_171, w_051_114);
  not1 I099_181(w_099_181, w_096_124);
  nand2 I099_182(w_099_182, w_019_357, w_095_022);
  or2  I099_183(w_099_183, w_039_170, w_004_004);
  and2 I099_187(w_099_187, w_048_427, w_081_582);
  nand2 I099_194(w_099_194, w_034_138, w_041_048);
  and2 I099_196(w_099_196, w_052_115, w_080_061);
  or2  I099_205(w_099_205, w_006_064, w_004_005);
  not1 I099_210(w_099_210, w_042_014);
  nand2 I099_230(w_099_230, w_070_147, w_039_183);
  nand2 I099_231(w_099_231, w_045_111, w_042_045);
  or2  I099_234(w_099_234, w_031_367, w_064_277);
  or2  I100_045(w_100_045, w_062_280, w_085_059);
  not1 I100_104(w_100_104, w_073_452);
  not1 I100_160(w_100_160, w_089_068);
  or2  I100_171(w_100_171, w_029_166, w_048_732);
  or2  I100_172(w_100_172, w_049_071, w_073_411);
  or2  I100_174(w_100_174, w_029_080, w_017_004);
  nand2 I100_201(w_100_201, w_091_082, w_000_775);
  not1 I100_202(w_100_202, w_099_194);
  or2  I100_225(w_100_225, w_046_328, w_003_186);
  and2 I100_257(w_100_257, w_029_138, w_041_120);
  or2  I100_283(w_100_283, w_067_939, w_047_475);
  and2 I100_305(w_100_305, w_070_847, w_059_152);
  or2  I100_313(w_100_313, w_037_052, w_094_763);
  not1 I100_335(w_100_335, w_084_033);
  not1 I100_368(w_100_368, w_051_540);
  not1 I100_392(w_100_392, w_086_482);
  nand2 I100_414(w_100_414, w_077_321, w_097_058);
  nand2 I100_429(w_100_429, w_007_216, w_024_057);
  or2  I100_533(w_100_533, w_058_040, w_084_257);
  or2  I100_556(w_100_556, w_050_322, w_080_032);
  not1 I100_565(w_100_565, w_058_220);
  nand2 I100_608(w_100_608, w_072_055, w_021_064);
  and2 I100_626(w_100_626, w_035_025, w_029_093);
  nand2 I100_642(w_100_642, w_060_241, w_091_170);
  and2 I100_657(w_100_657, w_076_591, w_033_015);
  nand2 I100_754(w_100_754, w_020_132, w_017_007);
  and2 I100_756(w_100_756, w_056_088, w_069_018);
  or2  I100_819(w_100_819, w_023_432, w_004_009);
  nand2 I100_847(w_100_847, w_091_233, w_025_606);
  and2 I100_914(w_100_914, w_064_375, w_042_014);
  nand2 I100_926(w_100_926, w_093_915, w_063_133);
  not1 I101_002(w_101_002, w_037_106);
  nand2 I101_012(w_101_012, w_019_294, w_013_407);
  and2 I101_016(w_101_016, w_097_057, w_100_847);
  nand2 I101_043(w_101_043, w_022_395, w_018_039);
  and2 I101_047(w_101_047, w_035_622, w_048_380);
  and2 I101_055(w_101_055, w_020_012, w_041_058);
  and2 I101_066(w_101_066, w_009_034, w_045_102);
  and2 I101_081(w_101_081, w_047_105, w_093_734);
  not1 I101_083(w_101_083, w_097_513);
  nand2 I101_094(w_101_094, w_057_385, w_099_157);
  or2  I101_106(w_101_106, w_035_313, w_049_651);
  nand2 I101_120(w_101_120, w_026_103, w_044_347);
  not1 I101_122(w_101_122, w_052_143);
  nand2 I101_128(w_101_128, w_078_251, w_072_067);
  and2 I101_130(w_101_130, w_097_441, w_070_647);
  nand2 I101_133(w_101_133, w_034_527, w_019_077);
  not1 I101_141(w_101_141, w_007_169);
  nand2 I101_143(w_101_143, w_049_075, w_006_235);
  or2  I101_144(w_101_144, w_062_037, w_095_019);
  or2  I101_148(w_101_148, w_089_006, w_037_131);
  or2  I101_152(w_101_152, w_037_163, w_004_011);
  or2  I101_153(w_101_153, w_037_040, w_085_006);
  nand2 I101_159(w_101_159, w_010_627, w_009_051);
  not1 I101_176(w_101_176, w_015_012);
  or2  I101_185(w_101_185, w_032_033, w_072_049);
  not1 I102_004(w_102_004, w_075_192);
  not1 I102_031(w_102_031, w_016_380);
  or2  I102_070(w_102_070, w_035_127, w_094_028);
  nand2 I102_094(w_102_094, w_046_194, w_043_038);
  not1 I102_124(w_102_124, w_040_201);
  nand2 I102_155(w_102_155, w_036_103, w_037_122);
  not1 I102_159(w_102_159, w_016_190);
  or2  I102_160(w_102_160, w_022_310, w_067_121);
  or2  I102_162(w_102_162, w_009_065, w_071_276);
  and2 I102_195(w_102_195, w_082_334, w_082_248);
  not1 I102_215(w_102_215, w_063_212);
  not1 I102_233(w_102_233, w_065_095);
  nand2 I102_298(w_102_298, w_031_204, w_040_217);
  nand2 I102_381(w_102_381, w_042_024, w_052_067);
  nand2 I102_400(w_102_400, w_066_345, w_081_374);
  not1 I102_450(w_102_450, w_067_075);
  and2 I102_563(w_102_563, w_038_224, w_015_255);
  nand2 I102_571(w_102_571, w_068_315, w_040_210);
  and2 I102_610(w_102_610, w_066_037, w_030_105);
  or2  I102_611(w_102_611, w_034_060, w_038_696);
  and2 I102_676(w_102_676, w_072_022, w_036_125);
  not1 I102_678(w_102_678, w_075_199);
  and2 I102_721(w_102_721, w_010_280, w_091_347);
  nand2 I102_750(w_102_750, w_077_347, w_036_068);
  and2 I102_754(w_102_754, w_008_820, w_081_360);
  and2 I102_779(w_102_779, w_101_159, w_062_165);
  not1 I103_011(w_103_011, w_083_618);
  or2  I103_040(w_103_040, w_052_121, w_080_046);
  and2 I103_049(w_103_049, w_083_147, w_021_007);
  nand2 I103_057(w_103_057, w_071_351, w_064_804);
  nand2 I103_063(w_103_063, w_101_153, w_095_008);
  and2 I103_160(w_103_160, w_011_485, w_044_188);
  nand2 I103_236(w_103_236, w_077_016, w_070_699);
  not1 I103_246(w_103_246, w_009_028);
  or2  I103_271(w_103_271, w_010_190, w_087_040);
  nand2 I103_302(w_103_302, w_063_181, w_008_015);
  not1 I103_306(w_103_306, w_041_039);
  and2 I103_361(w_103_361, w_023_291, w_047_436);
  and2 I103_444(w_103_444, w_021_089, w_057_021);
  or2  I103_447(w_103_447, w_067_085, w_058_341);
  not1 I103_498(w_103_498, w_019_116);
  or2  I103_582(w_103_582, w_015_142, w_059_193);
  or2  I103_640(w_103_640, w_092_038, w_085_010);
  and2 I103_649(w_103_649, w_076_433, w_030_294);
  and2 I103_658(w_103_658, w_074_273, w_061_238);
  nand2 I103_663(w_103_663, w_071_434, w_025_154);
  or2  I103_765(w_103_765, w_078_288, w_043_045);
  and2 I103_791(w_103_791, w_080_028, w_073_416);
  or2  I103_812(w_103_812, w_029_008, w_099_234);
  or2  I103_825(w_103_825, w_006_307, w_015_041);
  or2  I103_843(w_103_843, w_067_168, w_005_400);
  and2 I103_848(w_103_848, w_012_155, w_077_083);
  nand2 I103_894(w_103_894, w_062_029, w_026_307);
  or2  I104_012(w_104_012, w_061_333, w_008_355);
  or2  I104_013(w_104_013, w_031_303, w_079_218);
  or2  I104_019(w_104_019, w_091_507, w_070_730);
  and2 I104_024(w_104_024, w_032_753, w_092_282);
  or2  I104_035(w_104_035, w_015_595, w_026_349);
  or2  I104_036(w_104_036, w_020_075, w_090_271);
  or2  I104_038(w_104_038, w_095_150, w_101_122);
  and2 I104_042(w_104_042, w_072_014, w_085_022);
  nand2 I104_062(w_104_062, w_074_787, w_099_128);
  not1 I104_091(w_104_091, w_082_258);
  or2  I104_108(w_104_108, w_022_392, w_015_522);
  nand2 I104_116(w_104_116, w_030_149, w_007_097);
  nand2 I104_122(w_104_122, w_083_138, w_080_010);
  nand2 I104_140(w_104_140, w_090_026, w_092_011);
  nand2 I104_159(w_104_159, w_029_063, w_039_002);
  or2  I104_169(w_104_169, w_091_000, w_029_192);
  or2  I104_176(w_104_176, w_059_028, w_032_378);
  or2  I104_180(w_104_180, w_101_144, w_044_263);
  and2 I104_225(w_104_225, w_047_288, w_077_443);
  not1 I104_233(w_104_233, w_067_216);
  and2 I104_246(w_104_246, w_006_220, w_018_073);
  nand2 I104_250(w_104_250, w_026_424, w_010_494);
  nand2 I105_017(w_105_017, w_099_006, w_068_141);
  or2  I105_029(w_105_029, w_083_030, w_002_017);
  or2  I105_038(w_105_038, w_019_094, w_006_084);
  nand2 I105_044(w_105_044, w_052_148, w_036_061);
  and2 I105_117(w_105_117, w_026_438, w_059_058);
  and2 I105_189(w_105_189, w_102_124, w_008_631);
  nand2 I105_190(w_105_190, w_074_751, w_075_082);
  or2  I105_198(w_105_198, w_090_337, w_100_819);
  not1 I105_219(w_105_219, w_021_108);
  and2 I105_249(w_105_249, w_085_027, w_050_111);
  or2  I105_255(w_105_255, w_021_079, w_030_189);
  or2  I105_342(w_105_342, w_019_067, w_008_768);
  or2  I105_346(w_105_346, w_008_437, w_051_046);
  not1 I105_380(w_105_380, w_066_400);
  not1 I105_397(w_105_397, w_077_112);
  and2 I105_467(w_105_467, w_082_321, w_002_052);
  not1 I105_486(w_105_486, w_054_077);
  nand2 I105_498(w_105_498, w_037_000, w_018_086);
  nand2 I105_533(w_105_533, w_073_645, w_100_392);
  nand2 I105_626(w_105_626, w_012_533, w_051_240);
  nand2 I105_701(w_105_701, w_045_018, w_057_210);
  or2  I105_718(w_105_718, w_027_440, w_052_068);
  or2  I105_787(w_105_787, w_073_430, w_103_791);
  and2 I105_827(w_105_827, w_092_546, w_032_178);
  and2 I105_852(w_105_852, w_090_393, w_037_162);
  not1 I105_855(w_105_855, w_103_649);
  or2  I105_891(w_105_891, w_058_292, w_066_082);
  and2 I106_008(w_106_008, w_103_894, w_034_012);
  and2 I106_016(w_106_016, w_085_054, w_091_173);
  nand2 I106_018(w_106_018, w_036_146, w_009_035);
  and2 I106_049(w_106_049, w_002_108, w_009_066);
  not1 I106_103(w_106_103, w_016_029);
  not1 I106_115(w_106_115, w_004_019);
  not1 I106_137(w_106_137, w_061_069);
  or2  I106_141(w_106_141, w_040_168, w_054_251);
  not1 I106_167(w_106_167, w_077_069);
  not1 I106_205(w_106_205, w_097_231);
  not1 I106_224(w_106_224, w_029_072);
  not1 I106_237(w_106_237, w_086_012);
  nand2 I106_253(w_106_253, w_071_016, w_101_012);
  and2 I106_291(w_106_291, w_060_173, w_014_453);
  not1 I106_299(w_106_299, w_061_380);
  not1 I106_302(w_106_302, w_043_025);
  and2 I106_334(w_106_334, w_035_598, w_079_114);
  or2  I106_418(w_106_418, w_084_240, w_054_217);
  or2  I106_438(w_106_438, w_076_310, w_024_174);
  and2 I106_512(w_106_512, w_081_170, w_033_326);
  not1 I106_622(w_106_622, w_058_177);
  and2 I106_642(w_106_642, w_102_610, w_050_147);
  and2 I107_013(w_107_013, w_079_086, w_081_384);
  nand2 I107_014(w_107_014, w_098_036, w_020_020);
  nand2 I107_016(w_107_016, w_040_176, w_014_465);
  nand2 I107_018(w_107_018, w_006_158, w_026_436);
  or2  I107_019(w_107_019, w_056_284, w_062_021);
  or2  I107_021(w_107_021, w_067_728, w_071_158);
  or2  I107_022(w_107_022, w_023_493, w_104_038);
  nand2 I107_025(w_107_025, w_012_350, w_027_440);
  nand2 I107_027(w_107_027, w_059_279, w_086_006);
  and2 I107_030(w_107_030, w_013_096, w_007_048);
  or2  I107_038(w_107_038, w_079_136, w_051_306);
  and2 I107_046(w_107_046, w_064_482, w_101_143);
  and2 I107_050(w_107_050, w_053_654, w_084_428);
  or2  I107_072(w_107_072, w_094_292, w_104_012);
  or2  I107_077(w_107_077, w_079_051, w_105_249);
  and2 I107_082(w_107_082, w_102_070, w_039_381);
  and2 I107_088(w_107_088, w_097_030, w_028_427);
  nand2 I107_100(w_107_100, w_008_857, w_045_633);
  or2  I107_110(w_107_110, w_068_049, w_093_374);
  and2 I107_115(w_107_115, w_085_016, w_016_345);
  not1 I107_126(w_107_126, w_024_270);
  nand2 I107_127(w_107_127, w_074_258, w_008_708);
  nand2 I107_128(w_107_128, w_058_172, w_057_169);
  not1 I107_141(w_107_141, w_080_026);
  or2  I107_145(w_107_145, w_088_207, w_055_596);
  and2 I107_147(w_107_147, w_098_341, w_027_063);
  and2 I107_165(w_107_165, w_093_858, w_053_112);
  and2 I107_169(w_107_169, w_025_539, w_022_508);
  nand2 I107_180(w_107_180, w_073_331, w_038_713);
  or2  I107_181(w_107_181, w_019_277, w_044_110);
  and2 I107_182(w_107_182, w_041_044, w_103_361);
  nand2 I107_190(w_107_190, w_012_099, w_022_314);
  not1 I107_197(w_107_197, w_092_037);
  nand2 I107_203(w_107_203, w_065_551, w_053_193);
  not1 I107_206(w_107_206, w_018_196);
  and2 I108_000(w_108_000, w_017_005, w_027_055);
  not1 I108_001(w_108_001, w_088_063);
  not1 I108_002(w_108_002, w_075_024);
  not1 I108_003(w_108_003, w_086_242);
  and2 I108_005(w_108_005, w_076_352, w_091_190);
  and2 I108_006(w_108_006, w_060_240, w_024_397);
  nand2 I108_007(w_108_007, w_083_023, w_012_325);
  and2 I108_008(w_108_008, w_017_003, w_052_053);
  or2  I108_009(w_108_009, w_020_108, w_003_038);
  not1 I108_011(w_108_011, w_002_359);
  not1 I109_005(w_109_005, w_005_054);
  not1 I109_019(w_109_019, w_103_765);
  not1 I109_040(w_109_040, w_103_444);
  and2 I109_048(w_109_048, w_043_046, w_089_079);
  and2 I109_049(w_109_049, w_086_106, w_071_207);
  nand2 I109_058(w_109_058, w_106_512, w_011_203);
  or2  I109_068(w_109_068, w_084_610, w_012_178);
  nand2 I109_083(w_109_083, w_003_170, w_023_472);
  or2  I109_130(w_109_130, w_023_112, w_039_456);
  nand2 I109_133(w_109_133, w_083_291, w_067_226);
  or2  I109_142(w_109_142, w_062_478, w_058_250);
  and2 I109_145(w_109_145, w_105_342, w_075_284);
  or2  I109_147(w_109_147, w_049_363, w_071_125);
  and2 I109_150(w_109_150, w_055_129, w_033_547);
  or2  I109_153(w_109_153, w_063_104, w_063_083);
  nand2 I109_167(w_109_167, w_002_430, w_069_081);
  nand2 I109_169(w_109_169, w_093_169, w_090_328);
  or2  I109_178(w_109_178, w_045_548, w_072_010);
  not1 I109_232(w_109_232, w_097_602);
  nand2 I109_257(w_109_257, w_010_272, w_003_099);
  and2 I109_259(w_109_259, w_022_321, w_007_182);
  not1 I109_268(w_109_268, w_077_472);
  nand2 I109_275(w_109_275, w_011_649, w_087_313);
  and2 I109_283(w_109_283, w_029_178, w_081_563);
  not1 I110_005(w_110_005, w_048_490);
  and2 I110_010(w_110_010, w_023_477, w_055_010);
  and2 I110_041(w_110_041, w_066_213, w_018_133);
  nand2 I110_051(w_110_051, w_107_115, w_011_243);
  and2 I110_053(w_110_053, w_092_129, w_050_361);
  not1 I110_090(w_110_090, w_016_364);
  not1 I110_095(w_110_095, w_048_605);
  not1 I110_123(w_110_123, w_103_302);
  nand2 I110_143(w_110_143, w_030_001, w_099_020);
  nand2 I110_179(w_110_179, w_020_088, w_066_058);
  nand2 I110_195(w_110_195, w_057_337, w_107_077);
  or2  I110_232(w_110_232, w_033_645, w_052_137);
  nand2 I110_303(w_110_303, w_091_127, w_043_005);
  nand2 I110_347(w_110_347, w_076_236, w_092_092);
  and2 I110_350(w_110_350, w_108_006, w_095_131);
  not1 I110_404(w_110_404, w_047_272);
  and2 I110_414(w_110_414, w_009_033, w_095_101);
  not1 I110_455(w_110_455, w_033_311);
  nand2 I110_486(w_110_486, w_019_005, w_109_275);
  and2 I110_581(w_110_581, w_026_273, w_030_412);
  or2  I110_647(w_110_647, w_041_052, w_041_096);
  and2 I110_663(w_110_663, w_023_065, w_027_460);
  nand2 I110_664(w_110_664, w_073_550, w_080_080);
  and2 I111_018(w_111_018, w_051_313, w_024_291);
  or2  I111_028(w_111_028, w_008_914, w_109_048);
  or2  I111_031(w_111_031, w_000_064, w_024_131);
  or2  I111_044(w_111_044, w_096_381, w_053_835);
  or2  I111_048(w_111_048, w_071_431, w_057_322);
  nand2 I111_062(w_111_062, w_098_231, w_099_230);
  not1 I111_071(w_111_071, w_012_105);
  not1 I111_082(w_111_082, w_053_069);
  and2 I111_092(w_111_092, w_056_045, w_098_329);
  and2 I111_101(w_111_101, w_019_147, w_045_667);
  or2  I111_140(w_111_140, w_043_065, w_069_139);
  or2  I111_146(w_111_146, w_009_009, w_033_726);
  and2 I111_162(w_111_162, w_011_359, w_031_270);
  not1 I111_183(w_111_183, w_002_114);
  nand2 I111_196(w_111_196, w_007_367, w_110_041);
  or2  I111_202(w_111_202, w_028_079, w_015_424);
  not1 I111_206(w_111_206, w_035_400);
  or2  I111_238(w_111_238, w_011_112, w_021_185);
  and2 I111_291(w_111_291, w_021_052, w_044_139);
  and2 I111_312(w_111_312, w_013_238, w_060_071);
  and2 I111_339(w_111_339, w_087_304, w_100_414);
  not1 I112_013(w_112_013, w_041_077);
  not1 I112_029(w_112_029, w_014_289);
  not1 I112_048(w_112_048, w_036_013);
  nand2 I112_049(w_112_049, w_072_054, w_004_003);
  or2  I112_060(w_112_060, w_106_334, w_029_027);
  or2  I112_063(w_112_063, w_042_021, w_046_143);
  and2 I112_067(w_112_067, w_099_181, w_046_000);
  not1 I112_071(w_112_071, w_075_016);
  not1 I112_082(w_112_082, w_092_461);
  and2 I112_086(w_112_086, w_097_073, w_079_130);
  not1 I112_087(w_112_087, w_027_413);
  nand2 I112_088(w_112_088, w_065_944, w_068_056);
  nand2 I112_089(w_112_089, w_048_517, w_094_671);
  not1 I112_092(w_112_092, w_020_009);
  not1 I112_095(w_112_095, w_096_131);
  not1 I113_019(w_113_019, w_101_130);
  and2 I113_041(w_113_041, w_000_898, w_014_070);
  nand2 I113_070(w_113_070, w_096_075, w_019_406);
  nand2 I113_080(w_113_080, w_068_313, w_022_205);
  or2  I113_155(w_113_155, w_013_152, w_003_017);
  or2  I113_167(w_113_167, w_107_030, w_009_065);
  or2  I113_185(w_113_185, w_092_210, w_105_380);
  not1 I113_210(w_113_210, w_111_028);
  not1 I113_220(w_113_220, w_053_707);
  not1 I113_223(w_113_223, w_056_086);
  nand2 I113_239(w_113_239, w_100_756, w_005_346);
  not1 I113_248(w_113_248, w_016_278);
  not1 I113_299(w_113_299, w_078_051);
  not1 I113_304(w_113_304, w_090_252);
  and2 I113_305(w_113_305, w_051_392, w_065_556);
  and2 I113_322(w_113_322, w_052_035, w_008_405);
  not1 I113_331(w_113_331, w_022_270);
  or2  I113_351(w_113_351, w_082_257, w_082_194);
  and2 I113_372(w_113_372, w_043_062, w_082_004);
  not1 I113_423(w_113_423, w_020_126);
  not1 I113_428(w_113_428, w_079_162);
  nand2 I113_453(w_113_453, w_045_076, w_030_174);
  and2 I113_455(w_113_455, w_086_652, w_100_174);
  or2  I113_515(w_113_515, w_059_179, w_112_089);
  not1 I113_524(w_113_524, w_044_014);
  not1 I113_548(w_113_548, w_005_449);
  or2  I113_629(w_113_629, w_044_392, w_006_296);
  not1 I114_006(w_114_006, w_045_324);
  and2 I114_010(w_114_010, w_080_093, w_098_310);
  or2  I114_024(w_114_024, w_090_066, w_063_215);
  not1 I114_025(w_114_025, w_105_626);
  not1 I114_048(w_114_048, w_056_228);
  and2 I114_058(w_114_058, w_026_023, w_086_395);
  and2 I114_059(w_114_059, w_035_156, w_013_452);
  or2  I114_113(w_114_113, w_113_304, w_064_146);
  and2 I114_132(w_114_132, w_103_049, w_010_253);
  not1 I114_136(w_114_136, w_083_158);
  nand2 I114_187(w_114_187, w_050_413, w_099_205);
  nand2 I114_190(w_114_190, w_084_299, w_058_247);
  not1 I114_231(w_114_231, w_006_110);
  nand2 I114_283(w_114_283, w_031_232, w_083_220);
  not1 I114_286(w_114_286, w_093_911);
  nand2 I114_295(w_114_295, w_018_052, w_085_071);
  nand2 I114_302(w_114_302, w_077_281, w_081_212);
  nand2 I114_303(w_114_303, w_099_171, w_110_414);
  and2 I114_318(w_114_318, w_001_858, w_113_372);
  not1 I114_356(w_114_356, w_029_190);
  nand2 I114_366(w_114_366, w_097_634, w_084_035);
  or2  I115_003(w_115_003, w_032_151, w_017_012);
  and2 I115_019(w_115_019, w_109_133, w_016_156);
  and2 I115_021(w_115_021, w_103_843, w_094_055);
  and2 I115_025(w_115_025, w_008_917, w_076_360);
  or2  I115_030(w_115_030, w_047_386, w_020_126);
  nand2 I115_031(w_115_031, w_106_141, w_090_127);
  nand2 I115_034(w_115_034, w_004_007, w_039_332);
  nand2 I115_036(w_115_036, w_109_150, w_093_919);
  and2 I115_037(w_115_037, w_106_302, w_028_886);
  not1 I115_045(w_115_045, w_030_247);
  or2  I115_046(w_115_046, w_022_072, w_100_045);
  not1 I115_057(w_115_057, w_097_192);
  and2 I115_062(w_115_062, w_022_304, w_025_025);
  or2  I115_069(w_115_069, w_073_323, w_088_458);
  nand2 I115_071(w_115_071, w_096_120, w_014_101);
  or2  I115_073(w_115_073, w_056_048, w_108_007);
  nand2 I115_075(w_115_075, w_001_726, w_041_014);
  nand2 I115_079(w_115_079, w_060_341, w_092_644);
  and2 I115_084(w_115_084, w_108_006, w_089_078);
  nand2 I115_086(w_115_086, w_007_295, w_027_111);
  and2 I115_089(w_115_089, w_061_490, w_069_144);
  not1 I116_007(w_116_007, w_015_444);
  not1 I116_011(w_116_011, w_086_090);
  nand2 I116_013(w_116_013, w_067_242, w_046_182);
  or2  I116_014(w_116_014, w_037_079, w_040_219);
  or2  I116_018(w_116_018, w_011_409, w_067_920);
  nand2 I116_023(w_116_023, w_064_070, w_114_059);
  nand2 I116_027(w_116_027, w_054_085, w_024_507);
  not1 I116_032(w_116_032, w_043_013);
  nand2 I116_034(w_116_034, w_085_070, w_024_228);
  nand2 I116_035(w_116_035, w_068_068, w_010_697);
  and2 I116_037(w_116_037, w_080_108, w_111_044);
  not1 I116_038(w_116_038, w_007_302);
  and2 I116_040(w_116_040, w_038_548, w_008_616);
  and2 I116_041(w_116_041, w_024_196, w_099_120);
  nand2 I117_015(w_117_015, w_038_122, w_019_275);
  and2 I117_080(w_117_080, w_110_486, w_037_085);
  and2 I117_081(w_117_081, w_037_017, w_107_027);
  nand2 I117_082(w_117_082, w_040_116, w_043_060);
  or2  I117_087(w_117_087, w_083_111, w_082_028);
  or2  I117_100(w_117_100, w_037_105, w_075_108);
  or2  I117_105(w_117_105, w_106_167, w_087_069);
  and2 I117_112(w_117_112, w_111_238, w_008_033);
  not1 I117_135(w_117_135, w_074_463);
  nand2 I117_148(w_117_148, w_080_043, w_065_160);
  not1 I117_156(w_117_156, w_089_009);
  not1 I117_184(w_117_184, w_072_023);
  not1 I117_185(w_117_185, w_021_237);
  or2  I117_193(w_117_193, w_087_039, w_096_254);
  not1 I117_196(w_117_196, w_033_050);
  not1 I117_240(w_117_240, w_048_097);
  or2  I117_247(w_117_247, w_095_115, w_083_000);
  and2 I117_263(w_117_263, w_059_230, w_025_156);
  and2 I117_283(w_117_283, w_045_079, w_025_294);
  or2  I117_287(w_117_287, w_053_735, w_045_226);
  nand2 I117_290(w_117_290, w_094_115, w_040_142);
  nand2 I117_313(w_117_313, w_011_577, w_015_695);
  or2  I117_315(w_117_315, w_093_878, w_087_109);
  nand2 I117_324(w_117_324, w_063_357, w_098_278);
  or2  I118_035(w_118_035, w_008_494, w_107_013);
  not1 I118_085(w_118_085, w_015_000);
  or2  I118_091(w_118_091, w_091_403, w_016_247);
  nand2 I118_102(w_118_102, w_020_092, w_096_581);
  and2 I118_112(w_118_112, w_107_019, w_027_344);
  or2  I118_142(w_118_142, w_049_541, w_054_240);
  or2  I118_160(w_118_160, w_103_011, w_104_019);
  nand2 I118_180(w_118_180, w_014_329, w_086_428);
  not1 I118_181(w_118_181, w_061_063);
  not1 I118_184(w_118_184, w_117_240);
  or2  I118_190(w_118_190, w_094_113, w_040_132);
  and2 I118_192(w_118_192, w_078_028, w_060_155);
  nand2 I118_211(w_118_211, w_055_574, w_095_000);
  nand2 I118_217(w_118_217, w_022_511, w_072_055);
  or2  I118_234(w_118_234, w_040_325, w_071_057);
  nand2 I118_245(w_118_245, w_043_055, w_072_026);
  and2 I118_258(w_118_258, w_107_141, w_107_169);
  and2 I118_288(w_118_288, w_061_257, w_031_298);
  and2 I118_291(w_118_291, w_102_750, w_098_095);
  not1 I118_295(w_118_295, w_090_003);
  not1 I118_325(w_118_325, w_011_460);
  and2 I118_347(w_118_347, w_113_455, w_061_045);
  nand2 I118_350(w_118_350, w_069_017, w_031_161);
  nand2 I118_360(w_118_360, w_112_063, w_067_245);
  nand2 I118_384(w_118_384, w_008_314, w_091_279);
  nand2 I118_447(w_118_447, w_054_086, w_059_097);
  or2  I118_580(w_118_580, w_016_170, w_108_001);
  not1 I119_046(w_119_046, w_013_207);
  and2 I119_051(w_119_051, w_063_353, w_107_126);
  nand2 I119_080(w_119_080, w_064_665, w_114_318);
  and2 I119_117(w_119_117, w_008_566, w_003_039);
  and2 I119_119(w_119_119, w_026_051, w_080_032);
  not1 I119_121(w_119_121, w_077_047);
  or2  I119_140(w_119_140, w_008_574, w_014_024);
  or2  I119_148(w_119_148, w_040_314, w_093_423);
  nand2 I119_189(w_119_189, w_002_013, w_085_004);
  or2  I119_190(w_119_190, w_009_014, w_023_660);
  or2  I119_202(w_119_202, w_022_370, w_084_268);
  and2 I119_221(w_119_221, w_089_135, w_096_130);
  or2  I119_238(w_119_238, w_025_317, w_022_206);
  nand2 I119_285(w_119_285, w_072_046, w_094_150);
  nand2 I119_297(w_119_297, w_071_447, w_006_089);
  nand2 I119_299(w_119_299, w_095_017, w_064_076);
  nand2 I119_361(w_119_361, w_006_195, w_066_285);
  or2  I119_363(w_119_363, w_080_086, w_015_457);
  or2  I119_368(w_119_368, w_063_193, w_101_016);
  not1 I119_406(w_119_406, w_036_016);
  or2  I119_408(w_119_408, w_100_914, w_072_055);
  not1 I119_419(w_119_419, w_049_797);
  not1 I119_517(w_119_517, w_069_067);
  nand2 I119_561(w_119_561, w_100_754, w_009_027);
  or2  I119_575(w_119_575, w_045_111, w_019_374);
  or2  I120_005(w_120_005, w_064_247, w_034_033);
  and2 I120_013(w_120_013, w_005_141, w_009_053);
  and2 I120_016(w_120_016, w_119_238, w_057_275);
  and2 I120_018(w_120_018, w_000_979, w_056_190);
  or2  I120_021(w_120_021, w_000_232, w_083_087);
  or2  I120_032(w_120_032, w_033_546, w_116_018);
  nand2 I120_035(w_120_035, w_085_026, w_004_011);
  and2 I120_045(w_120_045, w_048_418, w_009_058);
  not1 I120_055(w_120_055, w_007_235);
  not1 I120_066(w_120_066, w_067_711);
  or2  I120_068(w_120_068, w_074_156, w_066_141);
  or2  I120_078(w_120_078, w_040_170, w_009_039);
  or2  I120_087(w_120_087, w_098_450, w_023_306);
  not1 I120_097(w_120_097, w_063_162);
  not1 I120_102(w_120_102, w_066_039);
  or2  I120_110(w_120_110, w_076_245, w_118_288);
  not1 I120_111(w_120_111, w_028_302);
  or2  I121_003(w_121_003, w_090_238, w_017_010);
  nand2 I121_077(w_121_077, w_119_368, w_116_027);
  or2  I121_081(w_121_081, w_011_281, w_114_366);
  or2  I121_124(w_121_124, w_096_086, w_002_020);
  nand2 I121_174(w_121_174, w_111_062, w_033_718);
  nand2 I121_175(w_121_175, w_002_274, w_036_122);
  not1 I121_178(w_121_178, w_056_077);
  or2  I121_182(w_121_182, w_011_059, w_065_363);
  and2 I121_260(w_121_260, w_049_944, w_045_223);
  or2  I121_301(w_121_301, w_041_035, w_095_028);
  and2 I121_331(w_121_331, w_118_447, w_070_551);
  not1 I121_354(w_121_354, w_111_048);
  nand2 I121_384(w_121_384, w_071_129, w_071_095);
  and2 I121_470(w_121_470, w_092_747, w_038_709);
  or2  I121_484(w_121_484, w_019_214, w_004_022);
  and2 I121_485(w_121_485, w_095_040, w_096_293);
  not1 I121_557(w_121_557, w_030_341);
  not1 I121_590(w_121_590, w_005_047);
  not1 I121_610(w_121_610, w_017_004);
  and2 I121_637(w_121_637, w_083_453, w_056_125);
  and2 I122_066(w_122_066, w_092_130, w_012_307);
  nand2 I122_069(w_122_069, w_101_128, w_087_049);
  or2  I122_088(w_122_088, w_001_751, w_088_098);
  not1 I122_135(w_122_135, w_082_344);
  and2 I122_137(w_122_137, w_079_247, w_067_294);
  or2  I122_208(w_122_208, w_041_060, w_100_335);
  nand2 I122_256(w_122_256, w_066_355, w_004_009);
  or2  I122_268(w_122_268, w_072_032, w_054_203);
  not1 I122_270(w_122_270, w_105_198);
  and2 I122_278(w_122_278, w_121_331, w_080_099);
  and2 I122_281(w_122_281, w_057_397, w_045_296);
  or2  I122_302(w_122_302, w_114_318, w_086_215);
  or2  I122_309(w_122_309, w_083_274, w_001_809);
  not1 I122_348(w_122_348, w_110_347);
  not1 I122_366(w_122_366, w_036_277);
  nand2 I122_385(w_122_385, w_031_010, w_030_408);
  nand2 I122_399(w_122_399, w_009_049, w_072_034);
  or2  I122_436(w_122_436, w_001_354, w_094_217);
  nand2 I122_447(w_122_447, w_066_392, w_114_113);
  not1 I122_458(w_122_458, w_073_030);
  and2 I122_472(w_122_472, w_048_738, w_090_121);
  not1 I123_011(w_123_011, w_039_190);
  and2 I123_025(w_123_025, w_082_061, w_117_185);
  and2 I123_027(w_123_027, w_106_115, w_101_002);
  and2 I123_048(w_123_048, w_026_037, w_103_658);
  not1 I123_062(w_123_062, w_080_016);
  not1 I123_066(w_123_066, w_083_435);
  nand2 I123_073(w_123_073, w_111_291, w_047_278);
  not1 I123_080(w_123_080, w_120_087);
  not1 I123_090(w_123_090, w_005_113);
  not1 I123_129(w_123_129, w_090_295);
  not1 I123_160(w_123_160, w_004_015);
  and2 I123_168(w_123_168, w_039_427, w_120_021);
  or2  I123_191(w_123_191, w_096_139, w_008_936);
  and2 I124_071(w_124_071, w_061_478, w_033_221);
  nand2 I124_091(w_124_091, w_032_705, w_118_295);
  and2 I124_128(w_124_128, w_041_122, w_052_026);
  or2  I124_134(w_124_134, w_099_158, w_004_038);
  not1 I124_142(w_124_142, w_100_608);
  or2  I124_157(w_124_157, w_096_168, w_085_024);
  not1 I124_235(w_124_235, w_068_081);
  or2  I124_283(w_124_283, w_026_032, w_104_035);
  and2 I124_305(w_124_305, w_048_078, w_019_116);
  nand2 I124_470(w_124_470, w_095_081, w_122_458);
  not1 I124_649(w_124_649, w_072_040);
  and2 I124_697(w_124_697, w_078_203, w_041_106);
  or2  I124_701(w_124_701, w_068_091, w_067_200);
  nand2 I125_007(w_125_007, w_112_067, w_079_163);
  nand2 I125_019(w_125_019, w_076_417, w_078_151);
  or2  I125_022(w_125_022, w_086_358, w_088_695);
  and2 I125_032(w_125_032, w_105_827, w_105_486);
  not1 I125_054(w_125_054, w_074_691);
  or2  I125_089(w_125_089, w_088_285, w_122_268);
  not1 I125_092(w_125_092, w_121_301);
  nand2 I125_101(w_125_101, w_082_206, w_085_037);
  and2 I125_124(w_125_124, w_117_193, w_114_187);
  not1 I125_129(w_125_129, w_054_227);
  nand2 I125_181(w_125_181, w_072_016, w_114_048);
  not1 I125_186(w_125_186, w_096_566);
  not1 I125_190(w_125_190, w_075_103);
  nand2 I125_199(w_125_199, w_013_176, w_114_006);
  not1 I125_207(w_125_207, w_068_306);
  not1 I125_213(w_125_213, w_014_099);
  or2  I126_034(w_126_034, w_020_134, w_106_642);
  and2 I126_053(w_126_053, w_113_548, w_019_074);
  or2  I126_112(w_126_112, w_009_065, w_069_107);
  and2 I126_118(w_126_118, w_118_350, w_002_094);
  nand2 I126_141(w_126_141, w_053_587, w_084_329);
  or2  I126_166(w_126_166, w_112_082, w_117_324);
  or2  I126_241(w_126_241, w_120_097, w_048_801);
  not1 I126_251(w_126_251, w_031_016);
  or2  I126_280(w_126_280, w_118_184, w_009_066);
  or2  I126_304(w_126_304, w_079_074, w_057_403);
  and2 I126_385(w_126_385, w_052_120, w_106_253);
  not1 I126_398(w_126_398, w_103_663);
  and2 I126_461(w_126_461, w_102_678, w_068_309);
  and2 I126_484(w_126_484, w_086_642, w_035_261);
  and2 I126_517(w_126_517, w_049_607, w_080_063);
  nand2 I127_023(w_127_023, w_073_409, w_026_325);
  or2  I127_029(w_127_029, w_103_640, w_025_531);
  and2 I127_065(w_127_065, w_019_279, w_003_053);
  or2  I127_068(w_127_068, w_047_401, w_118_112);
  or2  I127_071(w_127_071, w_113_331, w_086_701);
  or2  I127_076(w_127_076, w_029_089, w_099_196);
  or2  I127_077(w_127_077, w_012_143, w_078_161);
  and2 I127_085(w_127_085, w_090_283, w_037_189);
  or2  I127_095(w_127_095, w_106_049, w_029_099);
  and2 I127_109(w_127_109, w_099_130, w_034_044);
  nand2 I127_116(w_127_116, w_066_414, w_012_115);
  or2  I127_130(w_127_130, w_119_117, w_022_498);
  nand2 I127_141(w_127_141, w_047_124, w_079_219);
  or2  I128_003(w_128_003, w_083_242, w_002_019);
  not1 I128_004(w_128_004, w_017_015);
  not1 I128_005(w_128_005, w_101_055);
  nand2 I128_024(w_128_024, w_119_561, w_098_079);
  and2 I128_027(w_128_027, w_103_848, w_006_127);
  not1 I128_075(w_128_075, w_066_124);
  or2  I128_081(w_128_081, w_090_220, w_045_353);
  nand2 I128_094(w_128_094, w_005_422, w_123_073);
  nand2 I128_103(w_128_103, w_078_240, w_062_240);
  and2 I128_116(w_128_116, w_115_057, w_022_318);
  or2  I128_125(w_128_125, w_084_208, w_089_091);
  not1 I128_133(w_128_133, w_109_019);
  or2  I128_146(w_128_146, w_076_437, w_102_004);
  not1 I128_149(w_128_149, w_035_102);
  and2 I128_162(w_128_162, w_071_337, w_072_067);
  not1 I128_179(w_128_179, w_057_311);
  nand2 I128_199(w_128_199, w_073_034, w_012_474);
  and2 I128_201(w_128_201, w_081_016, w_006_009);
  nand2 I128_202(w_128_202, w_021_256, w_001_725);
  nand2 I128_203(w_128_203, w_042_026, w_034_184);
  nand2 I128_208(w_128_208, w_118_181, w_110_195);
  or2  I128_216(w_128_216, w_030_445, w_045_243);
  not1 I128_217(w_128_217, w_070_829);
  nand2 I128_220(w_128_220, w_036_013, w_006_015);
  not1 I128_239(w_128_239, w_100_283);
  nand2 I128_240(w_128_240, w_003_140, w_016_188);
  or2  I128_243(w_128_243, w_024_353, w_063_286);
  nand2 I129_000(w_129_000, w_034_122, w_073_214);
  and2 I129_001(w_129_001, w_085_006, w_022_479);
  and2 I129_004(w_129_004, w_082_097, w_112_060);
  nand2 I129_006(w_129_006, w_005_017, w_127_095);
  nand2 I129_008(w_129_008, w_115_071, w_090_250);
  nand2 I129_011(w_129_011, w_016_326, w_036_153);
  nand2 I129_016(w_129_016, w_090_336, w_010_652);
  and2 I129_022(w_129_022, w_122_069, w_106_018);
  and2 I129_024(w_129_024, w_036_056, w_113_629);
  or2  I130_002(w_130_002, w_113_423, w_073_643);
  not1 I130_104(w_130_104, w_091_173);
  and2 I130_213(w_130_213, w_062_166, w_027_614);
  nand2 I130_262(w_130_262, w_054_009, w_045_004);
  nand2 I130_269(w_130_269, w_056_099, w_063_360);
  not1 I130_271(w_130_271, w_104_250);
  or2  I130_291(w_130_291, w_056_256, w_070_289);
  and2 I130_340(w_130_340, w_032_790, w_128_125);
  not1 I130_422(w_130_422, w_099_231);
  and2 I130_545(w_130_545, w_093_227, w_009_007);
  not1 I130_620(w_130_620, w_128_199);
  and2 I130_661(w_130_661, w_062_312, w_125_213);
  not1 I130_726(w_130_726, w_118_245);
  not1 I130_747(w_130_747, w_017_003);
  not1 I130_767(w_130_767, w_057_024);
  or2  I130_860(w_130_860, w_040_245, w_118_325);
  and2 I130_866(w_130_866, w_047_443, w_017_021);
  not1 I130_882(w_130_882, w_044_193);
  not1 I130_917(w_130_917, w_017_021);
  nand2 I130_922(w_130_922, w_108_005, w_053_036);
  and2 I130_925(w_130_925, w_017_002, w_050_147);
  or2  I131_028(w_131_028, w_050_369, w_021_020);
  nand2 I131_070(w_131_070, w_076_006, w_083_259);
  and2 I131_081(w_131_081, w_059_169, w_083_653);
  nand2 I131_082(w_131_082, w_081_240, w_107_181);
  nand2 I131_094(w_131_094, w_093_825, w_077_041);
  or2  I131_100(w_131_100, w_058_225, w_033_771);
  and2 I131_116(w_131_116, w_106_299, w_002_102);
  not1 I131_120(w_131_120, w_069_022);
  or2  I131_121(w_131_121, w_048_029, w_074_754);
  and2 I131_181(w_131_181, w_130_422, w_100_202);
  and2 I131_185(w_131_185, w_030_089, w_078_287);
  not1 I131_578(w_131_578, w_111_202);
  or2  I131_617(w_131_617, w_078_017, w_055_192);
  and2 I131_632(w_131_632, w_085_039, w_089_079);
  not1 I131_634(w_131_634, w_102_215);
  or2  I131_682(w_131_682, w_043_001, w_130_545);
  not1 I131_685(w_131_685, w_027_285);
  or2  I132_033(w_132_033, w_015_703, w_125_124);
  nand2 I132_145(w_132_145, w_104_062, w_020_047);
  not1 I132_160(w_132_160, w_077_317);
  not1 I132_166(w_132_166, w_090_038);
  not1 I132_192(w_132_192, w_105_718);
  not1 I132_288(w_132_288, w_064_003);
  not1 I132_300(w_132_300, w_063_258);
  nand2 I132_338(w_132_338, w_114_286, w_078_077);
  not1 I132_353(w_132_353, w_034_806);
  nand2 I132_367(w_132_367, w_130_291, w_008_097);
  nand2 I132_383(w_132_383, w_055_159, w_125_186);
  nand2 I132_529(w_132_529, w_001_486, w_025_339);
  nand2 I133_010(w_133_010, w_127_068, w_081_134);
  or2  I133_016(w_133_016, w_119_148, w_022_375);
  and2 I133_024(w_133_024, w_096_097, w_004_013);
  and2 I133_057(w_133_057, w_128_027, w_093_200);
  and2 I133_086(w_133_086, w_070_446, w_037_066);
  and2 I133_097(w_133_097, w_066_282, w_091_125);
  or2  I133_158(w_133_158, w_085_051, w_117_184);
  or2  I133_177(w_133_177, w_126_241, w_074_681);
  or2  I133_236(w_133_236, w_039_074, w_054_218);
  and2 I133_252(w_133_252, w_022_271, w_046_067);
  not1 I133_266(w_133_266, w_040_274);
  and2 I133_298(w_133_298, w_050_255, w_060_095);
  nand2 I133_327(w_133_327, w_077_430, w_044_216);
  and2 I133_374(w_133_374, w_000_453, w_063_287);
  nand2 I133_416(w_133_416, w_096_114, w_072_011);
  not1 I133_430(w_133_430, w_059_044);
  not1 I133_516(w_133_516, w_001_320);
  or2  I133_521(w_133_521, w_124_283, w_131_028);
  nand2 I133_559(w_133_559, w_032_807, w_027_573);
  nand2 I133_790(w_133_790, w_030_371, w_023_064);
  nand2 I134_003(w_134_003, w_048_276, w_001_326);
  nand2 I134_010(w_134_010, w_032_233, w_126_141);
  and2 I134_097(w_134_097, w_117_135, w_085_003);
  or2  I134_127(w_134_127, w_073_090, w_026_392);
  nand2 I134_203(w_134_203, w_099_187, w_128_024);
  not1 I134_205(w_134_205, w_054_017);
  or2  I134_252(w_134_252, w_064_630, w_106_205);
  not1 I134_267(w_134_267, w_099_105);
  and2 I134_285(w_134_285, w_067_224, w_130_860);
  or2  I134_291(w_134_291, w_031_280, w_084_122);
  not1 I134_326(w_134_326, w_080_028);
  or2  I135_006(w_135_006, w_040_122, w_034_137);
  or2  I135_009(w_135_009, w_081_360, w_007_168);
  not1 I135_020(w_135_020, w_026_396);
  and2 I135_047(w_135_047, w_117_247, w_026_301);
  not1 I135_054(w_135_054, w_023_311);
  or2  I135_064(w_135_064, w_097_038, w_105_787);
  not1 I135_072(w_135_072, w_082_285);
  nand2 I135_074(w_135_074, w_122_436, w_032_570);
  nand2 I135_083(w_135_083, w_021_027, w_091_555);
  or2  I135_105(w_135_105, w_114_295, w_090_139);
  or2  I135_123(w_135_123, w_076_102, w_114_136);
  and2 I135_139(w_135_139, w_041_086, w_050_409);
  nand2 I135_203(w_135_203, w_076_356, w_022_294);
  or2  I135_204(w_135_204, w_127_029, w_128_203);
  or2  I135_207(w_135_207, w_101_185, w_019_011);
  not1 I135_219(w_135_219, w_125_129);
  and2 I135_221(w_135_221, w_132_160, w_008_912);
  not1 I135_226(w_135_226, w_021_152);
  not1 I136_012(w_136_012, w_081_017);
  nand2 I136_037(w_136_037, w_104_013, w_080_030);
  not1 I136_049(w_136_049, w_072_002);
  and2 I136_050(w_136_050, w_100_160, w_073_540);
  and2 I136_052(w_136_052, w_115_003, w_131_094);
  and2 I136_093(w_136_093, w_051_339, w_002_375);
  or2  I136_133(w_136_133, w_019_378, w_049_044);
  not1 I136_307(w_136_307, w_102_195);
  nand2 I136_319(w_136_319, w_086_725, w_031_324);
  or2  I136_504(w_136_504, w_043_046, w_103_271);
  or2  I136_588(w_136_588, w_004_008, w_103_246);
  and2 I136_694(w_136_694, w_124_697, w_029_007);
  and2 I136_920(w_136_920, w_025_015, w_021_266);
  nand2 I137_009(w_137_009, w_003_005, w_136_588);
  or2  I137_019(w_137_019, w_040_194, w_063_204);
  and2 I137_044(w_137_044, w_032_738, w_113_351);
  or2  I137_068(w_137_068, w_080_008, w_067_754);
  not1 I137_119(w_137_119, w_024_200);
  and2 I137_150(w_137_150, w_099_114, w_100_926);
  or2  I137_165(w_137_165, w_077_028, w_119_517);
  not1 I137_199(w_137_199, w_115_062);
  not1 I137_202(w_137_202, w_002_104);
  and2 I137_249(w_137_249, w_082_197, w_086_427);
  or2  I137_265(w_137_265, w_127_065, w_121_354);
  or2  I137_297(w_137_297, w_049_619, w_048_121);
  and2 I137_383(w_137_383, w_005_113, w_127_116);
  nand2 I137_394(w_137_394, w_058_324, w_134_285);
  not1 I137_424(w_137_424, w_108_002);
  nand2 I137_478(w_137_478, w_115_031, w_109_147);
  not1 I137_554(w_137_554, w_061_017);
  or2  I137_579(w_137_579, w_091_179, w_074_214);
  and2 I137_594(w_137_594, w_060_311, w_009_029);
  not1 I137_613(w_137_613, w_104_122);
  and2 I137_643(w_137_643, w_037_077, w_036_273);
  or2  I138_021(w_138_021, w_061_300, w_114_025);
  not1 I138_023(w_138_023, w_007_190);
  or2  I138_061(w_138_061, w_113_305, w_100_313);
  not1 I138_065(w_138_065, w_079_021);
  nand2 I138_084(w_138_084, w_017_007, w_026_049);
  or2  I138_127(w_138_127, w_114_024, w_087_177);
  and2 I138_145(w_138_145, w_074_383, w_039_128);
  and2 I138_147(w_138_147, w_033_314, w_049_270);
  not1 I138_183(w_138_183, w_110_143);
  nand2 I138_187(w_138_187, w_008_442, w_060_257);
  and2 I138_191(w_138_191, w_137_199, w_008_021);
  not1 I138_192(w_138_192, w_094_794);
  or2  I138_261(w_138_261, w_103_306, w_069_159);
  not1 I138_269(w_138_269, w_023_248);
  not1 I138_416(w_138_416, w_079_244);
  not1 I138_465(w_138_465, w_040_194);
  and2 I138_569(w_138_569, w_137_019, w_098_189);
  and2 I138_674(w_138_674, w_020_008, w_051_142);
  and2 I138_690(w_138_690, w_078_055, w_027_164);
  not1 I138_693(w_138_693, w_122_281);
  nand2 I138_726(w_138_726, w_123_129, w_073_747);
  and2 I138_738(w_138_738, w_131_116, w_030_202);
  and2 I139_001(w_139_001, w_065_941, w_032_267);
  not1 I139_002(w_139_002, w_134_127);
  and2 I139_003(w_139_003, w_039_149, w_119_406);
  not1 I139_005(w_139_005, w_070_748);
  or2  I139_006(w_139_006, w_121_182, w_101_016);
  and2 I139_007(w_139_007, w_138_192, w_047_357);
  not1 I139_009(w_139_009, w_115_037);
  nand2 I139_012(w_139_012, w_001_278, w_108_007);
  or2  I139_013(w_139_013, w_070_659, w_038_227);
  not1 I140_051(w_140_051, w_059_142);
  nand2 I140_101(w_140_101, w_007_282, w_065_750);
  or2  I140_150(w_140_150, w_026_351, w_102_450);
  or2  I140_219(w_140_219, w_066_465, w_044_174);
  or2  I140_273(w_140_273, w_014_104, w_053_055);
  nand2 I140_280(w_140_280, w_014_095, w_002_440);
  or2  I140_284(w_140_284, w_115_079, w_125_186);
  nand2 I140_289(w_140_289, w_105_038, w_063_315);
  or2  I140_308(w_140_308, w_114_190, w_116_023);
  or2  I140_319(w_140_319, w_011_072, w_117_082);
  or2  I140_333(w_140_333, w_042_094, w_091_214);
  and2 I140_630(w_140_630, w_138_269, w_130_269);
  or2  I141_052(w_141_052, w_078_042, w_111_018);
  or2  I141_061(w_141_061, w_045_076, w_138_023);
  nand2 I141_078(w_141_078, w_027_257, w_117_081);
  or2  I141_088(w_141_088, w_006_116, w_090_019);
  and2 I141_342(w_141_342, w_117_315, w_081_383);
  nand2 I141_358(w_141_358, w_032_421, w_026_341);
  and2 I141_409(w_141_409, w_048_218, w_124_701);
  nand2 I141_465(w_141_465, w_109_268, w_022_517);
  or2  I141_610(w_141_610, w_003_038, w_128_243);
  not1 I141_673(w_141_673, w_068_013);
  not1 I141_706(w_141_706, w_016_494);
  and2 I141_707(w_141_707, w_087_024, w_072_057);
  not1 I141_726(w_141_726, w_116_034);
  nand2 I141_823(w_141_823, w_109_153, w_012_212);
  not1 I142_011(w_142_011, w_021_076);
  or2  I142_062(w_142_062, w_034_435, w_035_277);
  nand2 I142_087(w_142_087, w_046_178, w_006_009);
  or2  I142_130(w_142_130, w_137_249, w_122_256);
  or2  I142_158(w_142_158, w_031_277, w_054_058);
  not1 I142_208(w_142_208, w_000_067);
  not1 I142_340(w_142_340, w_134_003);
  not1 I142_493(w_142_493, w_008_750);
  not1 I142_567(w_142_567, w_138_726);
  not1 I142_598(w_142_598, w_010_596);
  or2  I143_002(w_143_002, w_067_334, w_016_198);
  and2 I143_055(w_143_055, w_029_051, w_107_128);
  and2 I143_115(w_143_115, w_118_234, w_097_171);
  nand2 I143_129(w_143_129, w_028_767, w_098_451);
  and2 I143_159(w_143_159, w_130_661, w_137_297);
  not1 I143_241(w_143_241, w_021_163);
  not1 I143_253(w_143_253, w_082_240);
  and2 I143_256(w_143_256, w_002_255, w_123_168);
  not1 I143_279(w_143_279, w_122_135);
  not1 I143_311(w_143_311, w_100_104);
  or2  I143_328(w_143_328, w_090_212, w_118_347);
  or2  I143_356(w_143_356, w_013_300, w_112_029);
  and2 I143_402(w_143_402, w_026_017, w_126_484);
  not1 I143_418(w_143_418, w_021_046);
  and2 I143_510(w_143_510, w_135_054, w_124_071);
  and2 I143_549(w_143_549, w_015_440, w_113_210);
  not1 I143_575(w_143_577, w_143_576);
  not1 I143_576(w_143_578, w_143_577);
  or2  I143_577(w_143_576, w_031_011, w_143_578);
  and2 I144_022(w_144_022, w_073_490, w_052_046);
  nand2 I144_097(w_144_097, w_139_005, w_107_038);
  and2 I144_128(w_144_128, w_036_082, w_020_057);
  or2  I144_131(w_144_131, w_061_254, w_004_008);
  nand2 I144_158(w_144_158, w_026_116, w_009_046);
  or2  I144_234(w_144_234, w_093_241, w_117_112);
  not1 I144_282(w_144_282, w_035_460);
  and2 I144_289(w_144_289, w_060_171, w_051_360);
  nand2 I144_299(w_144_299, w_082_330, w_034_032);
  not1 I144_323(w_144_323, w_034_211);
  or2  I144_347(w_144_347, w_040_155, w_059_279);
  nand2 I144_394(w_144_394, w_045_029, w_026_142);
  nand2 I144_412(w_144_412, w_024_068, w_047_171);
  or2  I144_417(w_144_417, w_002_141, w_002_138);
  and2 I145_008(w_145_008, w_049_750, w_015_103);
  and2 I145_017(w_145_017, w_110_414, w_051_409);
  and2 I145_023(w_145_023, w_090_200, w_078_189);
  or2  I145_029(w_145_029, w_077_419, w_047_056);
  or2  I145_030(w_145_030, w_125_181, w_138_569);
  not1 I145_046(w_145_046, w_074_944);
  nand2 I145_047(w_145_047, w_006_021, w_000_155);
  or2  I145_050(w_145_050, w_005_303, w_067_615);
  and2 I145_052(w_145_052, w_118_180, w_011_457);
  nand2 I145_054(w_145_054, w_049_334, w_101_043);
  not1 I145_059(w_145_059, w_107_082);
  or2  I145_062(w_145_062, w_078_209, w_003_195);
  and2 I145_091(w_145_091, w_066_295, w_030_011);
  nand2 I145_097(w_145_097, w_040_117, w_051_336);
  or2  I146_012(w_146_012, w_077_191, w_076_273);
  and2 I146_065(w_146_065, w_006_259, w_012_343);
  or2  I146_073(w_146_073, w_128_103, w_012_543);
  not1 I146_106(w_146_106, w_119_297);
  and2 I146_122(w_146_122, w_006_140, w_041_062);
  and2 I146_124(w_146_124, w_109_068, w_034_042);
  not1 I146_129(w_146_129, w_082_228);
  not1 I146_170(w_146_170, w_090_160);
  nand2 I146_196(w_146_196, w_062_272, w_141_358);
  not1 I146_222(w_146_222, w_133_016);
  or2  I146_224(w_146_224, w_126_461, w_000_452);
  nand2 I146_231(w_146_231, w_041_012, w_053_238);
  nand2 I146_264(w_146_264, w_130_340, w_098_422);
  nand2 I146_274(w_146_274, w_024_129, w_021_277);
  and2 I146_296(w_146_296, w_071_003, w_129_000);
  or2  I146_314(w_146_314, w_017_024, w_000_671);
  not1 I146_328(w_146_328, w_010_530);
  and2 I147_047(w_147_047, w_096_118, w_013_315);
  nand2 I147_085(w_147_085, w_142_062, w_044_105);
  and2 I147_125(w_147_125, w_105_219, w_074_316);
  and2 I147_140(w_147_140, w_133_516, w_006_181);
  or2  I147_152(w_147_152, w_048_673, w_123_191);
  nand2 I147_189(w_147_189, w_002_372, w_011_272);
  and2 I147_213(w_147_213, w_085_017, w_059_180);
  not1 I147_263(w_147_263, w_057_467);
  nand2 I147_269(w_147_269, w_070_484, w_125_207);
  not1 I147_338(w_147_338, w_077_410);
  nand2 I147_491(w_147_491, w_020_057, w_106_137);
  not1 I147_520(w_147_520, w_071_116);
  nand2 I148_028(w_148_028, w_045_016, w_078_073);
  or2  I148_102(w_148_102, w_115_036, w_074_048);
  and2 I148_111(w_148_111, w_091_150, w_099_085);
  and2 I148_280(w_148_280, w_070_204, w_105_467);
  and2 I148_311(w_148_311, w_006_266, w_021_151);
  nand2 I148_327(w_148_327, w_012_062, w_021_130);
  nand2 I148_364(w_148_364, w_045_074, w_005_238);
  not1 I148_371(w_148_371, w_013_044);
  or2  I148_379(w_148_379, w_070_702, w_130_922);
  or2  I148_417(w_148_417, w_121_610, w_121_175);
  and2 I148_429(w_148_429, w_109_040, w_006_286);
  and2 I148_441(w_148_441, w_030_240, w_125_019);
  nand2 I148_444(w_148_444, w_068_175, w_107_022);
  and2 I148_460(w_148_460, w_080_071, w_001_323);
  or2  I148_495(w_148_495, w_043_048, w_097_069);
  not1 I149_065(w_149_065, w_041_121);
  nand2 I149_069(w_149_069, w_128_075, w_027_069);
  or2  I149_145(w_149_145, w_122_137, w_124_235);
  nand2 I149_161(w_149_161, w_051_382, w_049_657);
  or2  I149_232(w_149_232, w_137_594, w_018_074);
  or2  I149_239(w_149_239, w_079_182, w_001_044);
  and2 I149_266(w_149_266, w_000_649, w_034_451);
  nand2 I149_315(w_149_315, w_148_441, w_107_147);
  or2  I149_353(w_149_353, w_061_331, w_028_066);
  and2 I149_355(w_149_355, w_079_129, w_011_059);
  or2  I149_392(w_149_392, w_097_141, w_006_184);
  nand2 I149_449(w_149_449, w_091_206, w_010_539);
  nand2 I149_546(w_149_546, w_049_078, w_087_263);
  and2 I149_559(w_149_559, w_057_209, w_029_171);
  not1 I149_707(w_149_707, w_016_204);
  not1 I150_043(w_150_043, w_060_288);
  or2  I150_122(w_150_122, w_057_316, w_135_009);
  nand2 I150_140(w_150_140, w_017_012, w_100_171);
  not1 I150_154(w_150_154, w_024_158);
  or2  I150_160(w_150_160, w_036_171, w_117_015);
  not1 I150_194(w_150_194, w_036_282);
  and2 I151_000(w_151_000, w_059_237, w_113_223);
  or2  I151_003(w_151_003, w_125_092, w_002_215);
  or2  I151_034(w_151_034, w_087_329, w_094_217);
  or2  I151_109(w_151_109, w_098_315, w_017_022);
  or2  I151_196(w_151_196, w_100_565, w_128_003);
  not1 I151_210(w_151_210, w_143_402);
  not1 I151_223(w_151_223, w_054_020);
  not1 I151_226(w_151_226, w_093_258);
  nand2 I151_246(w_151_246, w_034_798, w_131_121);
  not1 I151_249(w_151_249, w_006_119);
  nand2 I151_255(w_151_255, w_122_088, w_040_033);
  nand2 I151_282(w_151_282, w_008_252, w_014_281);
  nand2 I151_283(w_151_283, w_072_029, w_066_119);
  or2  I151_288(w_151_288, w_048_296, w_034_729);
  and2 I151_298(w_151_298, w_128_220, w_000_871);
  not1 I151_307(w_151_307, w_133_010);
  nand2 I152_042(w_152_042, w_082_029, w_059_179);
  nand2 I152_059(w_152_059, w_076_269, w_114_302);
  nand2 I152_087(w_152_087, w_078_302, w_077_301);
  or2  I152_116(w_152_116, w_097_045, w_097_502);
  or2  I152_130(w_152_130, w_085_019, w_097_041);
  nand2 I152_278(w_152_278, w_133_252, w_136_920);
  or2  I152_395(w_152_395, w_085_059, w_025_614);
  or2  I152_422(w_152_422, w_023_531, w_148_327);
  not1 I152_460(w_152_460, w_018_180);
  nand2 I152_476(w_152_476, w_047_098, w_000_063);
  not1 I152_479(w_152_479, w_060_024);
  and2 I152_505(w_152_505, w_119_121, w_067_804);
  nand2 I152_611(w_152_611, w_001_641, w_137_044);
  nand2 I152_621(w_152_621, w_130_882, w_002_291);
  or2  I152_632(w_152_632, w_135_139, w_074_378);
  or2  I152_696(w_152_696, w_009_038, w_140_051);
  not1 I152_769(w_152_771, w_152_770);
  and2 I152_770(w_152_772, w_152_771, w_136_037);
  and2 I152_771(w_152_773, w_152_772, w_062_124);
  or2  I152_772(w_152_774, w_024_298, w_152_773);
  or2  I152_773(w_152_775, w_021_128, w_152_774);
  nand2 I152_774(w_152_770, w_152_786, w_152_775);
  nand2 I152_775(w_152_780, w_152_779, w_080_064);
  or2  I152_776(w_152_781, w_115_046, w_152_780);
  and2 I152_777(w_152_782, w_152_781, w_009_001);
  nand2 I152_778(w_152_783, w_152_782, w_110_404);
  or2  I152_779(w_152_784, w_124_142, w_152_783);
  not1 I152_780(w_152_779, w_152_770);
  and2 I152_781(w_152_786, w_080_075, w_152_784);
  or2  I153_056(w_153_056, w_017_000, w_084_234);
  and2 I153_072(w_153_072, w_021_126, w_012_327);
  and2 I153_114(w_153_114, w_095_128, w_060_155);
  nand2 I153_152(w_153_152, w_092_524, w_071_250);
  or2  I153_177(w_153_177, w_005_036, w_130_271);
  nand2 I153_210(w_153_210, w_057_067, w_131_634);
  or2  I153_385(w_153_385, w_111_140, w_145_017);
  not1 I153_415(w_153_415, w_138_147);
  or2  I153_457(w_153_457, w_102_571, w_010_253);
  nand2 I153_471(w_153_471, w_103_498, w_122_302);
  or2  I154_004(w_154_004, w_086_590, w_102_160);
  nand2 I154_083(w_154_083, w_145_030, w_019_130);
  not1 I154_113(w_154_113, w_078_009);
  not1 I154_137(w_154_137, w_087_144);
  nand2 I154_148(w_154_148, w_133_430, w_057_200);
  and2 I154_154(w_154_154, w_141_823, w_054_058);
  nand2 I154_243(w_154_243, w_115_084, w_007_275);
  nand2 I154_297(w_154_297, w_032_259, w_089_022);
  and2 I154_555(w_154_555, w_128_081, w_053_733);
  and2 I154_563(w_154_563, w_052_004, w_012_387);
  not1 I154_586(w_154_586, w_138_693);
  not1 I154_799(w_154_799, w_022_084);
  not1 I155_011(w_155_011, w_028_073);
  and2 I155_013(w_155_013, w_064_493, w_077_074);
  or2  I155_027(w_155_027, w_057_043, w_101_152);
  and2 I155_054(w_155_054, w_029_008, w_084_526);
  and2 I155_061(w_155_061, w_061_355, w_144_412);
  nand2 I155_079(w_155_079, w_149_546, w_079_172);
  not1 I155_108(w_155_108, w_096_248);
  or2  I155_109(w_155_109, w_110_053, w_119_408);
  not1 I155_124(w_155_124, w_067_945);
  not1 I156_092(w_156_092, w_035_292);
  and2 I156_302(w_156_302, w_060_269, w_148_371);
  nand2 I156_315(w_156_315, w_128_162, w_006_232);
  and2 I156_422(w_156_422, w_002_497, w_138_061);
  and2 I156_456(w_156_456, w_036_112, w_081_090);
  not1 I156_622(w_156_622, w_102_159);
  and2 I156_661(w_156_661, w_125_054, w_140_308);
  not1 I156_707(w_156_709, w_156_708);
  or2  I156_708(w_156_710, w_156_709, w_071_284);
  not1 I156_709(w_156_711, w_156_710);
  or2  I156_710(w_156_712, w_038_157, w_156_711);
  nand2 I156_711(w_156_713, w_101_141, w_156_712);
  nand2 I156_712(w_156_708, w_058_002, w_156_713);
  nand2 I157_016(w_157_016, w_055_105, w_105_498);
  not1 I157_038(w_157_038, w_119_190);
  and2 I157_105(w_157_105, w_084_029, w_032_012);
  nand2 I157_180(w_157_180, w_086_666, w_071_137);
  and2 I157_528(w_157_528, w_008_848, w_138_674);
  nand2 I157_539(w_157_539, w_110_090, w_038_689);
  or2  I157_557(w_157_557, w_100_626, w_131_185);
  nand2 I157_739(w_157_739, w_121_637, w_061_247);
  and2 I157_754(w_157_754, w_103_040, w_116_035);
  nand2 I157_814(w_157_814, w_014_159, w_136_049);
  nand2 I158_009(w_158_009, w_010_086, w_112_089);
  and2 I158_069(w_158_069, w_136_050, w_113_019);
  not1 I158_076(w_158_076, w_060_307);
  not1 I158_079(w_158_079, w_122_066);
  and2 I158_082(w_158_082, w_118_192, w_008_306);
  or2  I158_145(w_158_145, w_071_239, w_049_459);
  or2  I158_198(w_158_198, w_105_117, w_059_121);
  not1 I158_213(w_158_213, w_118_291);
  not1 I158_225(w_158_225, w_104_091);
  not1 I158_356(w_158_356, w_113_322);
  and2 I158_392(w_158_392, w_105_701, w_086_099);
  and2 I158_546(w_158_546, w_020_126, w_058_050);
  or2  I158_633(w_158_633, w_091_036, w_138_187);
  and2 I158_643(w_158_643, w_032_003, w_016_317);
  not1 I158_841(w_158_841, w_154_154);
  not1 I158_847(w_158_847, w_073_059);
  or2  I159_004(w_159_004, w_088_404, w_056_092);
  and2 I159_062(w_159_062, w_153_471, w_051_031);
  nand2 I159_064(w_159_064, w_044_083, w_029_024);
  not1 I159_074(w_159_074, w_062_353);
  or2  I159_102(w_159_102, w_000_670, w_148_311);
  or2  I159_149(w_159_149, w_016_210, w_013_143);
  or2  I159_169(w_159_169, w_156_092, w_002_225);
  not1 I159_192(w_159_192, w_016_213);
  not1 I159_221(w_159_221, w_118_142);
  and2 I159_227(w_159_227, w_069_125, w_103_812);
  or2  I159_245(w_159_245, w_015_704, w_001_452);
  or2  I159_253(w_159_253, w_129_001, w_141_061);
  and2 I159_260(w_159_260, w_040_017, w_076_056);
  nand2 I159_264(w_159_264, w_071_306, w_088_179);
  not1 I159_285(w_159_285, w_095_182);
  nand2 I160_072(w_160_072, w_016_217, w_035_554);
  and2 I160_073(w_160_073, w_122_399, w_035_074);
  nand2 I160_081(w_160_081, w_102_676, w_005_548);
  not1 I160_088(w_160_088, w_151_246);
  nand2 I160_155(w_160_155, w_066_054, w_136_133);
  or2  I160_181(w_160_181, w_017_012, w_138_261);
  nand2 I160_320(w_160_320, w_137_265, w_159_227);
  not1 I160_359(w_160_359, w_078_034);
  and2 I160_431(w_160_431, w_068_234, w_128_240);
  not1 I160_599(w_160_599, w_136_319);
  nand2 I160_638(w_160_638, w_082_033, w_085_050);
  or2  I161_081(w_161_081, w_133_024, w_072_019);
  nand2 I161_104(w_161_104, w_112_086, w_034_100);
  nand2 I161_124(w_161_124, w_135_203, w_152_422);
  and2 I161_221(w_161_221, w_063_200, w_033_420);
  nand2 I162_051(w_162_051, w_064_264, w_010_259);
  and2 I162_133(w_162_133, w_150_194, w_020_037);
  or2  I162_139(w_162_139, w_093_107, w_095_181);
  or2  I162_146(w_162_146, w_014_222, w_083_095);
  not1 I162_154(w_162_154, w_089_090);
  not1 I162_173(w_162_173, w_096_299);
  or2  I162_181(w_162_181, w_033_499, w_130_767);
  or2  I162_210(w_162_210, w_007_405, w_125_199);
  or2  I162_244(w_162_244, w_090_268, w_017_024);
  nand2 I162_249(w_162_249, w_022_290, w_145_008);
  not1 I162_298(w_162_298, w_037_020);
  nand2 I162_321(w_162_321, w_023_088, w_147_263);
  and2 I162_326(w_162_326, w_026_355, w_095_054);
  not1 I162_359(w_162_359, w_092_239);
  and2 I162_396(w_162_396, w_047_208, w_078_297);
  not1 I162_427(w_162_427, w_155_054);
  not1 I162_466(w_162_466, w_021_058);
  nand2 I163_002(w_163_002, w_158_633, w_133_236);
  and2 I163_047(w_163_047, w_015_013, w_154_243);
  nand2 I163_068(w_163_068, w_086_202, w_139_005);
  nand2 I163_095(w_163_095, w_148_379, w_061_360);
  nand2 I163_120(w_163_120, w_138_065, w_045_563);
  not1 I163_176(w_163_176, w_023_271);
  nand2 I163_181(w_163_181, w_059_116, w_022_464);
  not1 I163_215(w_163_215, w_010_264);
  or2  I163_235(w_163_235, w_025_556, w_107_197);
  or2  I163_237(w_163_237, w_077_385, w_118_085);
  and2 I163_341(w_163_341, w_131_100, w_159_004);
  not1 I163_536(w_163_536, w_090_332);
  or2  I163_642(w_163_642, w_118_160, w_047_244);
  nand2 I164_035(w_164_035, w_148_111, w_033_598);
  or2  I164_037(w_164_037, w_028_025, w_031_454);
  or2  I164_042(w_164_042, w_089_127, w_046_572);
  nand2 I164_069(w_164_069, w_113_524, w_111_312);
  or2  I164_109(w_164_109, w_000_396, w_148_102);
  and2 I164_129(w_164_129, w_037_011, w_010_703);
  not1 I164_131(w_164_131, w_145_047);
  or2  I164_155(w_164_155, w_107_110, w_040_043);
  and2 I164_183(w_164_183, w_077_197, w_061_433);
  and2 I164_186(w_164_186, w_153_072, w_096_346);
  or2  I164_193(w_164_193, w_066_209, w_162_139);
  not1 I164_314(w_164_314, w_021_105);
  and2 I164_326(w_164_326, w_027_568, w_004_033);
  not1 I164_375(w_164_375, w_043_017);
  or2  I165_098(w_165_098, w_136_093, w_004_012);
  nand2 I165_120(w_165_120, w_080_038, w_153_457);
  not1 I165_140(w_165_140, w_010_798);
  and2 I165_187(w_165_187, w_136_012, w_107_014);
  and2 I165_203(w_165_203, w_110_455, w_148_417);
  nand2 I165_277(w_165_277, w_105_189, w_136_694);
  and2 I165_362(w_165_362, w_148_444, w_028_506);
  or2  I165_550(w_165_550, w_025_478, w_043_058);
  or2  I166_015(w_166_015, w_111_339, w_151_307);
  not1 I166_020(w_166_020, w_128_149);
  and2 I166_041(w_166_041, w_083_441, w_015_676);
  not1 I166_047(w_166_047, w_160_359);
  or2  I166_120(w_166_120, w_023_503, w_158_841);
  nand2 I166_219(w_166_219, w_070_117, w_109_167);
  nand2 I166_269(w_166_269, w_025_428, w_068_128);
  not1 I166_294(w_166_294, w_135_204);
  and2 I166_327(w_166_327, w_071_112, w_135_072);
  not1 I166_331(w_166_331, w_029_034);
  or2  I166_360(w_166_360, w_037_006, w_058_182);
  nand2 I166_531(w_166_531, w_139_003, w_120_018);
  and2 I167_031(w_167_031, w_057_008, w_079_078);
  and2 I167_042(w_167_042, w_106_291, w_159_074);
  not1 I167_069(w_167_069, w_026_209);
  or2  I167_234(w_167_234, w_084_535, w_054_246);
  or2  I167_265(w_167_265, w_148_495, w_133_158);
  not1 I167_275(w_167_275, w_147_491);
  nand2 I167_280(w_167_280, w_163_536, w_154_083);
  nand2 I167_290(w_167_290, w_068_005, w_076_008);
  and2 I167_406(w_167_406, w_067_265, w_002_272);
  or2  I167_416(w_167_416, w_121_590, w_138_021);
  not1 I167_458(w_167_458, w_123_066);
  nand2 I167_495(w_167_495, w_130_620, w_155_011);
  and2 I167_557(w_167_557, w_013_350, w_064_041);
  or2  I167_656(w_167_656, w_158_009, w_039_362);
  and2 I168_104(w_168_104, w_006_295, w_028_024);
  nand2 I168_128(w_168_128, w_128_162, w_019_073);
  and2 I168_133(w_168_133, w_003_047, w_104_225);
  nand2 I168_361(w_168_361, w_107_182, w_018_015);
  not1 I168_387(w_168_387, w_167_557);
  not1 I168_412(w_168_412, w_050_294);
  and2 I168_541(w_168_541, w_106_103, w_048_101);
  or2  I168_767(w_168_767, w_144_097, w_137_119);
  or2  I169_017(w_169_017, w_005_237, w_062_032);
  nand2 I169_021(w_169_021, w_018_079, w_130_747);
  and2 I169_022(w_169_022, w_141_052, w_084_294);
  nand2 I169_034(w_169_034, w_103_582, w_003_121);
  not1 I169_036(w_169_036, w_166_120);
  or2  I169_042(w_169_042, w_039_284, w_097_583);
  or2  I169_050(w_169_050, w_045_170, w_168_128);
  and2 I169_068(w_169_068, w_154_148, w_168_133);
  not1 I170_032(w_170_032, w_013_375);
  or2  I170_045(w_170_045, w_067_178, w_072_042);
  nand2 I170_166(w_170_166, w_011_041, w_005_325);
  or2  I170_171(w_170_171, w_021_075, w_054_240);
  or2  I170_199(w_170_199, w_042_077, w_090_209);
  not1 I170_220(w_170_220, w_064_347);
  not1 I170_275(w_170_275, w_115_069);
  not1 I170_289(w_170_289, w_062_292);
  not1 I170_407(w_170_407, w_160_081);
  or2  I171_042(w_171_042, w_154_555, w_144_131);
  nand2 I171_188(w_171_188, w_085_041, w_152_087);
  nand2 I171_189(w_171_189, w_160_181, w_141_409);
  nand2 I171_215(w_171_215, w_013_317, w_099_035);
  nand2 I171_242(w_171_242, w_160_638, w_138_465);
  or2  I171_264(w_171_264, w_153_210, w_023_175);
  and2 I171_280(w_171_280, w_001_603, w_055_105);
  nand2 I171_296(w_171_296, w_099_210, w_110_663);
  or2  I171_326(w_171_326, w_041_036, w_157_739);
  or2  I171_333(w_171_333, w_042_011, w_065_742);
  and2 I171_359(w_171_359, w_127_085, w_016_010);
  nand2 I171_369(w_171_369, w_031_171, w_040_095);
  or2  I171_391(w_171_391, w_030_358, w_126_034);
  not1 I171_472(w_171_472, w_157_016);
  and2 I172_030(w_172_030, w_052_150, w_080_038);
  and2 I172_060(w_172_060, w_158_213, w_060_320);
  and2 I172_109(w_172_109, w_028_369, w_100_225);
  nand2 I172_299(w_172_299, w_052_078, w_122_447);
  and2 I172_315(w_172_315, w_049_338, w_054_234);
  or2  I172_357(w_172_357, w_170_032, w_140_273);
  and2 I172_365(w_172_365, w_153_385, w_157_557);
  or2  I172_388(w_172_388, w_137_613, w_078_102);
  and2 I172_405(w_172_405, w_149_449, w_013_119);
  not1 I173_043(w_173_043, w_054_203);
  and2 I173_069(w_173_069, w_019_138, w_025_657);
  nand2 I173_110(w_173_110, w_107_165, w_143_510);
  and2 I173_120(w_173_120, w_064_032, w_161_104);
  or2  I173_158(w_173_158, w_159_221, w_068_191);
  not1 I173_432(w_173_432, w_110_095);
  or2  I174_149(w_174_149, w_151_226, w_173_120);
  and2 I174_189(w_174_189, w_111_031, w_034_220);
  not1 I174_269(w_174_269, w_118_580);
  or2  I174_453(w_174_453, w_101_106, w_035_092);
  not1 I174_516(w_174_516, w_069_084);
  nand2 I174_538(w_174_538, w_115_034, w_078_271);
  and2 I174_762(w_174_762, w_030_166, w_050_192);
  and2 I174_857(w_174_857, w_146_222, w_036_234);
  nand2 I175_182(w_175_182, w_096_229, w_152_505);
  nand2 I175_456(w_175_456, w_010_315, w_167_290);
  or2  I175_551(w_175_551, w_094_710, w_162_146);
  nand2 I175_828(w_175_828, w_137_068, w_089_074);
  or2  I176_067(w_176_067, w_026_325, w_003_110);
  nand2 I176_154(w_176_154, w_148_429, w_047_146);
  or2  I176_180(w_176_180, w_035_492, w_006_237);
  or2  I176_201(w_176_201, w_148_460, w_063_195);
  or2  I176_270(w_176_270, w_081_270, w_162_298);
  nand2 I176_361(w_176_361, w_084_125, w_113_428);
  not1 I176_380(w_176_380, w_160_320);
  not1 I176_479(w_176_479, w_125_101);
  nand2 I177_030(w_177_030, w_083_266, w_108_008);
  and2 I177_072(w_177_072, w_072_003, w_132_383);
  and2 I177_095(w_177_095, w_059_258, w_147_189);
  nand2 I177_278(w_177_278, w_131_685, w_172_109);
  not1 I177_347(w_177_347, w_052_164);
  not1 I177_395(w_177_395, w_028_033);
  not1 I177_524(w_177_524, w_094_781);
  not1 I177_549(w_177_549, w_107_203);
  nand2 I177_639(w_177_639, w_031_198, w_066_368);
  nand2 I177_701(w_177_701, w_018_153, w_043_041);
  not1 I177_790(w_177_790, w_170_289);
  nand2 I177_863(w_177_863, w_148_028, w_054_221);
  and2 I177_912(w_177_912, w_031_251, w_076_192);
  or2  I178_014(w_178_014, w_093_279, w_160_088);
  or2  I178_016(w_178_016, w_133_521, w_087_053);
  or2  I178_351(w_178_351, w_100_533, w_072_026);
  or2  I178_504(w_178_504, w_113_453, w_003_163);
  nand2 I178_590(w_178_590, w_029_190, w_015_201);
  and2 I178_600(w_178_600, w_128_202, w_152_042);
  and2 I178_883(w_178_883, w_078_212, w_086_116);
  nand2 I178_943(w_178_943, w_022_339, w_147_085);
  and2 I179_022(w_179_022, w_137_383, w_167_495);
  nand2 I179_218(w_179_218, w_043_013, w_089_024);
  nand2 I179_549(w_179_549, w_045_629, w_176_479);
  nand2 I179_713(w_179_713, w_026_194, w_094_134);
  or2  I179_724(w_179_724, w_022_406, w_076_330);
  not1 I179_888(w_179_888, w_154_799);
  and2 I180_005(w_180_005, w_168_387, w_047_348);
  or2  I180_050(w_180_050, w_117_080, w_122_278);
  not1 I180_075(w_180_075, w_062_032);
  nand2 I180_160(w_180_160, w_063_053, w_152_460);
  not1 I180_172(w_180_172, w_060_153);
  or2  I180_210(w_180_210, w_177_701, w_063_205);
  nand2 I180_269(w_180_269, w_071_007, w_071_253);
  nand2 I180_305(w_180_305, w_158_392, w_164_193);
  or2  I180_333(w_180_333, w_158_079, w_085_011);
  or2  I181_103(w_181_103, w_169_021, w_084_012);
  and2 I181_162(w_181_162, w_010_653, w_085_016);
  or2  I181_211(w_181_211, w_140_284, w_114_231);
  and2 I181_234(w_181_234, w_151_249, w_120_045);
  and2 I181_388(w_181_388, w_141_465, w_104_036);
  nand2 I181_495(w_181_495, w_053_102, w_088_108);
  or2  I181_516(w_181_516, w_076_227, w_133_097);
  and2 I181_790(w_181_790, w_109_259, w_022_033);
  and2 I181_802(w_181_802, w_050_058, w_005_017);
  nand2 I182_038(w_182_038, w_021_133, w_089_031);
  nand2 I182_039(w_182_039, w_076_012, w_028_855);
  or2  I182_073(w_182_073, w_138_416, w_159_260);
  not1 I182_091(w_182_091, w_143_055);
  nand2 I182_115(w_182_115, w_100_429, w_175_182);
  or2  I182_120(w_182_120, w_108_009, w_040_254);
  nand2 I182_122(w_182_122, w_080_011, w_115_021);
  not1 I182_159(w_182_159, w_019_168);
  or2  I182_188(w_182_188, w_038_156, w_164_109);
  nand2 I182_193(w_182_193, w_092_706, w_153_152);
  or2  I182_210(w_182_210, w_002_357, w_034_588);
  and2 I182_223(w_182_223, w_131_082, w_047_067);
  or2  I182_227(w_182_227, w_071_115, w_093_353);
  not1 I182_228(w_182_228, w_168_361);
  and2 I182_274(w_182_274, w_124_134, w_007_265);
  nand2 I183_035(w_183_035, w_120_016, w_142_493);
  not1 I183_041(w_183_041, w_172_357);
  not1 I183_053(w_183_053, w_051_527);
  or2  I183_067(w_183_067, w_140_280, w_107_088);
  or2  I183_070(w_183_070, w_101_047, w_061_095);
  nand2 I183_110(w_183_110, w_001_042, w_126_053);
  not1 I183_224(w_183_224, w_182_227);
  nand2 I184_008(w_184_008, w_149_707, w_042_070);
  or2  I184_039(w_184_039, w_105_852, w_009_068);
  and2 I184_049(w_184_049, w_082_253, w_038_119);
  or2  I184_085(w_184_085, w_093_720, w_079_046);
  not1 I184_157(w_184_157, w_109_142);
  not1 I184_173(w_184_173, w_142_158);
  nand2 I184_191(w_184_191, w_004_003, w_143_129);
  nand2 I184_243(w_184_243, w_062_436, w_012_288);
  and2 I185_031(w_185_031, w_072_057, w_073_705);
  not1 I185_061(w_185_061, w_006_268);
  or2  I185_078(w_185_078, w_124_157, w_031_003);
  nand2 I185_100(w_185_100, w_182_159, w_169_036);
  not1 I185_103(w_185_103, w_041_050);
  not1 I185_118(w_185_118, w_083_022);
  or2  I185_149(w_185_149, w_029_026, w_092_680);
  not1 I185_202(w_185_202, w_072_060);
  nand2 I185_277(w_185_277, w_077_107, w_132_145);
  and2 I186_001(w_186_001, w_083_238, w_107_050);
  and2 I186_007(w_186_007, w_119_575, w_070_784);
  or2  I186_042(w_186_042, w_107_100, w_119_221);
  not1 I186_070(w_186_070, w_061_009);
  not1 I186_198(w_186_198, w_132_033);
  not1 I186_304(w_186_304, w_021_184);
  or2  I186_442(w_186_442, w_054_128, w_025_155);
  or2  I186_479(w_186_479, w_080_056, w_077_449);
  not1 I186_544(w_186_544, w_145_059);
  or2  I186_609(w_186_609, w_066_072, w_105_029);
  or2  I186_618(w_186_618, w_181_802, w_119_140);
  and2 I186_642(w_186_642, w_135_020, w_122_309);
  not1 I187_011(w_187_011, w_126_304);
  not1 I187_022(w_187_022, w_027_742);
  nand2 I187_024(w_187_024, w_118_091, w_003_216);
  or2  I187_096(w_187_096, w_134_252, w_108_008);
  or2  I187_099(w_187_099, w_110_664, w_114_010);
  and2 I187_131(w_187_131, w_128_133, w_100_657);
  and2 I187_148(w_187_148, w_082_013, w_031_103);
  nand2 I187_153(w_187_153, w_134_205, w_151_288);
  not1 I187_161(w_187_161, w_100_257);
  and2 I187_175(w_187_175, w_010_473, w_025_067);
  not1 I187_183(w_187_183, w_053_030);
  nand2 I187_203(w_187_203, w_103_063, w_146_122);
  not1 I188_073(w_188_073, w_087_226);
  or2  I188_087(w_188_087, w_149_355, w_128_208);
  or2  I188_123(w_188_123, w_030_005, w_045_160);
  not1 I188_161(w_188_161, w_119_361);
  or2  I188_427(w_188_427, w_114_132, w_074_915);
  or2  I188_430(w_188_430, w_030_312, w_147_125);
  nand2 I188_491(w_188_491, w_181_211, w_070_027);
  nand2 I188_534(w_188_536, w_188_535, w_072_033);
  or2  I188_535(w_188_537, w_029_056, w_188_536);
  nand2 I188_536(w_188_538, w_117_313, w_188_537);
  and2 I188_537(w_188_539, w_188_538, w_110_350);
  or2  I188_538(w_188_535, w_188_550, w_188_539);
  and2 I188_539(w_188_544, w_188_543, w_085_055);
  nand2 I188_540(w_188_545, w_188_544, w_133_374);
  not1 I188_541(w_188_546, w_188_545);
  and2 I188_542(w_188_547, w_031_219, w_188_546);
  not1 I188_543(w_188_548, w_188_547);
  not1 I188_544(w_188_543, w_188_535);
  and2 I188_545(w_188_550, w_140_289, w_188_548);
  nand2 I189_071(w_189_071, w_073_339, w_184_008);
  nand2 I189_115(w_189_115, w_063_054, w_116_013);
  or2  I189_117(w_189_117, w_052_008, w_022_307);
  and2 I189_298(w_189_298, w_014_363, w_014_415);
  not1 I189_346(w_189_346, w_070_381);
  nand2 I189_525(w_189_525, w_158_847, w_080_058);
  not1 I189_974(w_189_974, w_121_178);
  nand2 I190_000(w_190_000, w_162_051, w_052_012);
  not1 I190_068(w_190_068, w_025_020);
  nand2 I190_168(w_190_168, w_160_431, w_167_234);
  or2  I190_222(w_190_222, w_000_865, w_162_249);
  not1 I190_237(w_190_237, w_189_974);
  not1 I190_261(w_190_261, w_000_665);
  not1 I190_289(w_190_289, w_177_790);
  nand2 I190_348(w_190_348, w_126_517, w_041_037);
  nand2 I190_394(w_190_394, w_054_163, w_070_493);
  or2  I191_036(w_191_036, w_155_079, w_090_038);
  or2  I191_037(w_191_037, w_063_084, w_074_488);
  not1 I191_083(w_191_083, w_097_636);
  nand2 I191_118(w_191_118, w_083_109, w_065_686);
  and2 I191_135(w_191_135, w_181_162, w_032_057);
  and2 I191_142(w_191_142, w_097_001, w_155_124);
  nand2 I191_174(w_191_174, w_052_073, w_101_176);
  or2  I191_211(w_191_211, w_162_173, w_003_103);
  and2 I191_278(w_191_278, w_129_024, w_119_189);
  and2 I191_294(w_191_294, w_190_068, w_066_115);
  or2  I191_316(w_191_316, w_040_173, w_015_504);
  and2 I191_325(w_191_325, w_104_233, w_054_179);
  and2 I191_385(w_191_385, w_036_177, w_105_891);
  and2 I191_392(w_191_392, w_096_028, w_126_280);
  or2  I192_000(w_192_000, w_129_016, w_121_470);
  nand2 I192_001(w_192_001, w_165_362, w_152_476);
  or2  I192_002(w_192_002, w_063_266, w_077_323);
  nand2 I193_003(w_193_003, w_130_866, w_171_326);
  nand2 I193_042(w_193_042, w_073_663, w_177_278);
  or2  I193_197(w_193_197, w_157_754, w_158_069);
  and2 I193_252(w_193_252, w_059_134, w_068_010);
  or2  I193_290(w_193_290, w_158_225, w_068_025);
  or2  I193_291(w_193_291, w_058_080, w_090_079);
  not1 I193_314(w_193_314, w_096_348);
  nand2 I193_340(w_193_340, w_074_467, w_135_207);
  nand2 I193_416(w_193_416, w_111_196, w_034_217);
  or2  I193_418(w_193_418, w_047_230, w_179_888);
  not1 I193_454(w_193_454, w_021_129);
  not1 I193_669(w_193_669, w_080_009);
  nand2 I194_011(w_194_011, w_049_414, w_140_150);
  nand2 I194_077(w_194_077, w_045_255, w_051_178);
  or2  I194_089(w_194_089, w_174_189, w_087_044);
  or2  I194_211(w_194_211, w_035_532, w_026_353);
  not1 I194_219(w_194_219, w_012_139);
  not1 I194_268(w_194_268, w_100_368);
  and2 I194_283(w_194_283, w_013_261, w_171_242);
  and2 I194_433(w_194_433, w_014_289, w_187_099);
  nand2 I194_453(w_194_453, w_111_071, w_043_059);
  nand2 I194_471(w_194_471, w_167_656, w_018_122);
  and2 I194_495(w_194_495, w_018_163, w_104_140);
  nand2 I194_593(w_194_593, w_072_030, w_035_024);
  not1 I194_699(w_194_699, w_021_008);
  not1 I194_909(w_194_909, w_032_060);
  and2 I195_029(w_195_029, w_105_533, w_079_218);
  or2  I195_070(w_195_070, w_174_149, w_112_095);
  or2  I195_082(w_195_082, w_058_360, w_169_017);
  not1 I195_181(w_195_181, w_065_380);
  nand2 I195_256(w_195_256, w_077_193, w_099_102);
  or2  I195_335(w_195_335, w_097_077, w_095_164);
  nand2 I195_348(w_195_348, w_176_067, w_083_439);
  not1 I195_487(w_195_487, w_061_123);
  not1 I195_517(w_195_517, w_109_147);
  or2  I196_045(w_196_045, w_067_724, w_148_364);
  and2 I196_274(w_196_274, w_119_285, w_016_354);
  or2  I196_306(w_196_306, w_145_052, w_086_596);
  and2 I196_453(w_196_453, w_128_179, w_132_288);
  not1 I196_712(w_196_712, w_047_203);
  not1 I196_728(w_196_728, w_060_313);
  not1 I196_808(w_196_808, w_053_005);
  not1 I197_140(w_197_140, w_099_182);
  nand2 I197_143(w_197_143, w_172_365, w_076_388);
  and2 I197_189(w_197_189, w_081_590, w_169_068);
  and2 I197_237(w_197_237, w_098_048, w_115_045);
  nand2 I197_352(w_197_352, w_186_642, w_083_310);
  or2  I197_422(w_197_422, w_131_617, w_155_109);
  not1 I197_541(w_197_541, w_023_628);
  nand2 I197_674(w_197_674, w_109_257, w_112_092);
  nand2 I197_746(w_197_746, w_141_610, w_035_473);
  and2 I197_778(w_197_778, w_190_168, w_024_335);
  or2  I197_838(w_197_838, w_101_094, w_083_649);
  and2 I197_896(w_197_896, w_164_037, w_144_158);
  and2 I198_040(w_198_040, w_082_163, w_004_037);
  and2 I198_074(w_198_074, w_020_004, w_185_031);
  or2  I198_220(w_198_220, w_116_037, w_047_474);
  nand2 I198_315(w_198_315, w_037_036, w_089_019);
  or2  I198_322(w_198_322, w_042_056, w_151_003);
  not1 I198_330(w_198_330, w_006_094);
  or2  I198_578(w_198_578, w_018_032, w_054_201);
  or2  I198_741(w_198_741, w_194_283, w_085_058);
  and2 I199_044(w_199_044, w_148_280, w_184_173);
  nand2 I199_056(w_199_056, w_194_593, w_167_031);
  and2 I199_060(w_199_060, w_024_382, w_085_043);
  or2  I199_131(w_199_131, w_130_726, w_134_291);
  and2 I199_419(w_199_419, w_004_009, w_083_153);
  nand2 I199_751(w_199_751, w_155_013, w_129_000);
  and2 I199_795(w_199_795, w_170_171, w_091_232);
  or2  I199_829(w_199_829, w_074_692, w_166_327);
  and2 I200_029(w_200_029, w_092_083, w_135_219);
  and2 I200_166(w_200_166, w_010_440, w_005_391);
  or2  I200_262(w_200_262, w_088_619, w_114_303);
  nand2 I200_683(w_200_683, w_099_183, w_002_310);
  nand2 I201_076(w_201_076, w_076_166, w_090_270);
  nand2 I201_095(w_201_095, w_066_511, w_191_278);
  nand2 I201_276(w_201_276, w_133_086, w_120_078);
  not1 I201_514(w_201_514, w_035_268);
  not1 I201_655(w_201_655, w_107_016);
  nand2 I201_698(w_201_698, w_063_107, w_122_385);
  not1 I201_719(w_201_719, w_109_058);
  nand2 I202_003(w_202_003, w_159_227, w_150_043);
  and2 I202_009(w_202_009, w_121_557, w_015_661);
  nand2 I202_011(w_202_011, w_091_408, w_004_003);
  nand2 I202_012(w_202_012, w_057_445, w_156_661);
  not1 I202_015(w_202_015, w_015_048);
  nand2 I202_018(w_202_018, w_166_047, w_062_100);
  not1 I202_019(w_202_019, w_047_279);
  nand2 I202_020(w_202_020, w_079_234, w_146_231);
  or2  I203_061(w_203_061, w_074_607, w_018_159);
  and2 I203_082(w_203_082, w_189_525, w_022_081);
  or2  I203_098(w_203_098, w_017_024, w_177_639);
  nand2 I203_110(w_203_110, w_079_068, w_142_598);
  nand2 I203_156(w_203_156, w_001_443, w_011_376);
  or2  I203_258(w_203_258, w_149_353, w_039_119);
  and2 I203_304(w_203_304, w_117_156, w_051_417);
  or2  I203_312(w_203_312, w_101_066, w_202_020);
  nand2 I203_407(w_203_407, w_173_158, w_008_619);
  not1 I203_512(w_203_512, w_167_265);
  not1 I204_218(w_204_218, w_198_074);
  and2 I204_257(w_204_257, w_154_563, w_149_266);
  not1 I204_342(w_204_342, w_120_087);
  and2 I204_363(w_204_363, w_120_111, w_057_157);
  nand2 I205_113(w_205_113, w_202_011, w_070_488);
  and2 I205_126(w_205_126, w_057_051, w_138_127);
  nand2 I205_427(w_205_427, w_028_406, w_107_018);
  not1 I205_566(w_205_566, w_151_210);
  nand2 I206_057(w_206_057, w_141_726, w_192_001);
  or2  I206_126(w_206_126, w_112_088, w_011_395);
  or2  I206_334(w_206_334, w_158_082, w_136_052);
  and2 I207_005(w_207_005, w_189_117, w_090_224);
  nand2 I207_023(w_207_023, w_113_248, w_010_767);
  or2  I207_104(w_207_104, w_091_316, w_064_695);
  or2  I207_147(w_207_147, w_078_028, w_163_047);
  nand2 I207_226(w_207_226, w_041_111, w_024_501);
  and2 I207_236(w_207_236, w_137_478, w_125_022);
  and2 I207_244(w_207_244, w_127_023, w_030_477);
  nand2 I207_353(w_207_353, w_153_114, w_112_087);
  nand2 I208_026(w_208_026, w_098_035, w_039_062);
  not1 I208_028(w_208_028, w_031_215);
  nand2 I208_032(w_208_032, w_185_118, w_043_009);
  or2  I208_267(w_208_267, w_086_705, w_182_188);
  or2  I209_171(w_209_171, w_037_079, w_137_424);
  not1 I209_179(w_209_179, w_163_176);
  nand2 I209_180(w_209_180, w_033_218, w_088_151);
  and2 I209_203(w_209_203, w_143_256, w_161_221);
  nand2 I210_314(w_210_314, w_055_245, w_101_081);
  nand2 I210_523(w_210_523, w_171_189, w_121_484);
  nand2 I210_574(w_210_574, w_166_041, w_126_398);
  or2  I210_681(w_210_681, w_056_065, w_010_795);
  nand2 I211_029(w_211_029, w_103_447, w_167_280);
  and2 I211_040(w_211_040, w_099_036, w_025_614);
  or2  I211_050(w_211_050, w_123_080, w_110_232);
  or2  I211_052(w_211_052, w_096_100, w_024_255);
  not1 I211_133(w_211_133, w_108_003);
  or2  I211_150(w_211_150, w_184_191, w_026_265);
  and2 I211_241(w_211_241, w_132_353, w_182_073);
  or2  I211_276(w_211_276, w_159_245, w_021_139);
  not1 I211_498(w_211_498, w_193_003);
  or2  I211_528(w_211_528, w_182_120, w_086_577);
  or2  I212_013(w_212_013, w_095_030, w_069_000);
  not1 I212_084(w_212_084, w_076_363);
  or2  I212_102(w_212_102, w_196_808, w_092_038);
  and2 I212_109(w_212_109, w_109_232, w_108_002);
  or2  I213_041(w_213_041, w_017_012, w_146_124);
  not1 I213_433(w_213_433, w_157_105);
  and2 I213_538(w_213_538, w_026_279, w_041_061);
  nand2 I214_005(w_214_005, w_183_067, w_163_235);
  or2  I214_027(w_214_027, w_019_344, w_143_328);
  or2  I214_039(w_214_039, w_124_305, w_018_117);
  or2  I214_052(w_214_052, w_120_013, w_146_264);
  or2  I214_070(w_214_070, w_107_145, w_124_091);
  or2  I214_075(w_214_075, w_044_203, w_149_145);
  nand2 I214_092(w_214_092, w_164_375, w_102_031);
  not1 I214_100(w_214_100, w_041_011);
  not1 I214_107(w_214_107, w_088_163);
  nand2 I215_092(w_215_092, w_195_181, w_154_586);
  and2 I215_170(w_215_170, w_213_538, w_193_314);
  nand2 I215_267(w_215_267, w_151_223, w_200_029);
  and2 I215_322(w_215_322, w_116_014, w_163_341);
  and2 I215_422(w_215_422, w_043_047, w_161_081);
  or2  I215_428(w_215_428, w_173_432, w_125_032);
  and2 I215_565(w_215_565, w_146_196, w_028_456);
  and2 I216_050(w_216_050, w_214_100, w_016_021);
  not1 I216_102(w_216_102, w_041_068);
  not1 I216_126(w_216_126, w_137_009);
  or2  I216_129(w_216_129, w_029_056, w_158_076);
  or2  I217_209(w_217_209, w_089_095, w_129_000);
  and2 I217_279(w_217_279, w_085_026, w_214_039);
  or2  I217_372(w_217_372, w_001_842, w_066_224);
  nand2 I217_797(w_217_797, w_078_221, w_110_303);
  or2  I217_819(w_217_819, w_165_277, w_084_114);
  nand2 I218_004(w_218_004, w_007_363, w_163_068);
  not1 I218_016(w_218_016, w_110_179);
  or2  I218_141(w_218_141, w_191_392, w_168_541);
  or2  I218_204(w_218_204, w_199_044, w_041_118);
  nand2 I218_428(w_218_428, w_163_215, w_039_289);
  and2 I218_582(w_218_582, w_146_012, w_083_021);
  or2  I219_030(w_219_030, w_017_015, w_111_082);
  and2 I219_038(w_219_038, w_163_642, w_083_596);
  not1 I219_064(w_219_064, w_176_270);
  nand2 I219_069(w_219_069, w_000_602, w_123_090);
  not1 I219_146(w_219_146, w_104_108);
  nand2 I219_217(w_219_217, w_155_108, w_009_048);
  or2  I219_277(w_219_277, w_028_429, w_001_219);
  and2 I220_034(w_220_034, w_140_319, w_110_647);
  or2  I220_055(w_220_055, w_024_435, w_044_043);
  or2  I220_257(w_220_257, w_190_394, w_117_100);
  or2  I220_604(w_220_604, w_208_028, w_202_009);
  and2 I220_608(w_220_608, w_144_022, w_218_428);
  and2 I220_821(w_220_821, w_177_863, w_121_003);
  or2  I221_070(w_221_070, w_160_073, w_152_130);
  nand2 I221_136(w_221_136, w_211_241, w_180_075);
  or2  I221_396(w_221_396, w_103_236, w_118_360);
  nand2 I221_550(w_221_550, w_181_516, w_211_498);
  not1 I222_045(w_222_045, w_085_060);
  not1 I222_259(w_222_259, w_108_011);
  and2 I222_477(w_222_477, w_069_137, w_202_015);
  and2 I222_662(w_222_662, w_025_412, w_111_183);
  nand2 I223_023(w_223_023, w_117_283, w_119_363);
  or2  I223_141(w_223_141, w_047_001, w_033_325);
  nand2 I223_157(w_223_157, w_220_055, w_119_419);
  and2 I223_278(w_223_278, w_093_137, w_064_271);
  or2  I223_379(w_223_379, w_205_427, w_076_617);
  or2  I223_493(w_223_493, w_083_651, w_208_267);
  and2 I223_582(w_223_582, w_144_289, w_006_046);
  not1 I223_631(w_223_631, w_066_371);
  and2 I223_840(w_223_840, w_022_100, w_042_059);
  not1 I223_925(w_223_925, w_005_397);
  not1 I224_009(w_224_009, w_023_435);
  or2  I224_038(w_224_038, w_028_143, w_182_122);
  not1 I224_041(w_224_041, w_205_126);
  nand2 I224_042(w_224_042, w_088_030, w_100_556);
  and2 I224_052(w_224_052, w_025_553, w_002_054);
  or2  I224_058(w_224_058, w_115_086, w_049_309);
  and2 I224_075(w_224_075, w_114_058, w_183_224);
  or2  I225_002(w_225_002, w_108_011, w_030_281);
  or2  I225_022(w_225_022, w_218_204, w_156_315);
  or2  I225_026(w_225_026, w_189_346, w_153_056);
  nand2 I226_000(w_226_000, w_152_611, w_054_023);
  or2  I226_001(w_226_001, w_071_428, w_120_066);
  nand2 I226_005(w_226_005, w_057_063, w_113_185);
  not1 I226_008(w_226_008, w_167_406);
  and2 I226_010(w_226_010, w_113_155, w_187_148);
  nand2 I226_013(w_226_013, w_124_128, w_042_011);
  not1 I227_012(w_227_012, w_037_133);
  not1 I227_067(w_227_067, w_136_504);
  not1 I227_199(w_227_199, w_081_538);
  nand2 I227_260(w_227_260, w_178_883, w_191_142);
  and2 I227_408(w_227_408, w_062_432, w_075_051);
  not1 I227_416(w_227_416, w_144_417);
  and2 I227_522(w_227_522, w_076_136, w_018_176);
  and2 I227_547(w_227_547, w_207_226, w_117_087);
  nand2 I228_267(w_228_267, w_128_116, w_143_311);
  nand2 I228_288(w_228_288, w_135_105, w_071_174);
  and2 I228_329(w_228_329, w_116_040, w_090_086);
  or2  I228_637(w_228_637, w_161_124, w_165_203);
  and2 I228_745(w_228_745, w_006_096, w_164_035);
  or2  I229_076(w_229_076, w_069_126, w_157_814);
  nand2 I229_125(w_229_125, w_193_291, w_097_501);
  not1 I229_274(w_229_274, w_193_454);
  and2 I229_295(w_229_295, w_068_157, w_164_069);
  and2 I230_032(w_230_032, w_199_795, w_205_566);
  or2  I230_036(w_230_036, w_115_089, w_194_495);
  nand2 I230_048(w_230_048, w_001_079, w_067_516);
  or2  I230_082(w_230_082, w_162_359, w_054_191);
  nand2 I230_238(w_230_238, w_073_005, w_139_009);
  and2 I230_246(w_230_246, w_047_427, w_117_287);
  not1 I230_248(w_230_248, w_171_391);
  nand2 I230_251(w_230_251, w_032_777, w_014_279);
  not1 I230_252(w_230_252, w_049_965);
  and2 I230_262(w_230_262, w_043_051, w_109_005);
  or2  I230_295(w_230_295, w_002_299, w_014_088);
  and2 I231_002(w_231_002, w_230_262, w_037_049);
  and2 I231_026(w_231_026, w_000_497, w_015_003);
  and2 I231_036(w_231_036, w_133_559, w_080_043);
  not1 I231_049(w_231_049, w_130_104);
  and2 I231_057(w_231_057, w_046_333, w_147_338);
  and2 I231_083(w_231_083, w_012_253, w_119_202);
  or2  I232_008(w_232_008, w_025_238, w_065_631);
  nand2 I232_029(w_232_029, w_003_212, w_121_174);
  not1 I232_032(w_232_032, w_223_278);
  not1 I232_146(w_232_146, w_075_285);
  or2  I232_202(w_232_202, w_065_305, w_210_314);
  or2  I232_235(w_232_235, w_029_157, w_140_219);
  not1 I232_363(w_232_363, w_156_422);
  not1 I233_078(w_233_078, w_187_183);
  and2 I233_128(w_233_128, w_179_022, w_092_503);
  nand2 I233_319(w_233_319, w_203_098, w_079_231);
  nand2 I233_342(w_233_342, w_203_061, w_199_060);
  and2 I233_384(w_233_384, w_226_010, w_180_160);
  nand2 I233_391(w_233_391, w_159_102, w_159_264);
  nand2 I234_050(w_234_050, w_011_415, w_105_190);
  nand2 I234_515(w_234_515, w_057_350, w_049_525);
  not1 I234_554(w_234_554, w_046_734);
  and2 I235_019(w_235_019, w_014_549, w_120_055);
  nand2 I235_058(w_235_058, w_104_116, w_035_129);
  and2 I235_140(w_235_140, w_025_307, w_111_092);
  or2  I236_047(w_236_047, w_195_517, w_199_829);
  and2 I236_050(w_236_050, w_105_255, w_045_043);
  not1 I236_151(w_236_151, w_182_039);
  or2  I236_154(w_236_154, w_108_011, w_068_145);
  nand2 I236_162(w_236_162, w_055_210, w_086_709);
  nand2 I236_300(w_236_300, w_215_565, w_177_072);
  or2  I236_315(w_236_315, w_013_108, w_128_004);
  or2  I236_410(w_236_410, w_059_018, w_196_453);
  and2 I236_606(w_236_606, w_192_001, w_181_790);
  or2  I237_228(w_237_228, w_183_035, w_213_433);
  nand2 I237_276(w_237_276, w_102_381, w_171_188);
  and2 I237_376(w_237_376, w_164_183, w_187_024);
  nand2 I237_379(w_237_379, w_141_673, w_201_276);
  not1 I237_423(w_237_423, w_202_018);
  and2 I238_033(w_238_033, w_078_121, w_050_102);
  not1 I238_053(w_238_053, w_000_929);
  not1 I238_080(w_238_080, w_015_521);
  and2 I238_159(w_238_159, w_124_470, w_042_108);
  not1 I238_218(w_238_218, w_061_528);
  or2  I238_231(w_238_231, w_058_006, w_201_719);
  or2  I238_251(w_238_251, w_046_367, w_087_145);
  not1 I238_285(w_238_285, w_159_253);
  not1 I238_312(w_238_312, w_055_138);
  or2  I238_350(w_238_350, w_236_050, w_133_327);
  or2  I238_360(w_238_360, w_072_017, w_046_171);
  nand2 I238_389(w_238_389, w_135_047, w_040_058);
  or2  I239_054(w_239_054, w_059_318, w_181_103);
  and2 I239_174(w_239_174, w_133_298, w_152_632);
  or2  I239_183(w_239_183, w_238_350, w_118_035);
  nand2 I239_648(w_239_648, w_022_412, w_044_156);
  not1 I239_678(w_239_678, w_226_008);
  not1 I239_728(w_239_728, w_135_064);
  and2 I240_011(w_240_011, w_052_022, w_155_061);
  or2  I240_178(w_240_178, w_078_132, w_005_296);
  and2 I240_754(w_240_754, w_126_385, w_226_000);
  nand2 I240_813(w_240_815, w_240_814, w_236_047);
  nand2 I240_814(w_240_816, w_240_815, w_053_676);
  nand2 I240_815(w_240_817, w_046_120, w_240_816);
  nand2 I240_816(w_240_818, w_219_146, w_240_817);
  nand2 I240_817(w_240_819, w_129_008, w_240_818);
  nand2 I240_818(w_240_820, w_128_005, w_240_819);
  not1 I240_819(w_240_821, w_240_820);
  not1 I240_820(w_240_814, w_240_821);
  or2  I241_027(w_241_027, w_121_384, w_217_797);
  and2 I241_065(w_241_065, w_075_258, w_169_050);
  nand2 I241_142(w_241_142, w_235_019, w_121_077);
  nand2 I241_276(w_241_276, w_201_095, w_014_576);
  nand2 I241_336(w_241_336, w_082_232, w_011_138);
  not1 I241_344(w_241_344, w_029_070);
  and2 I242_106(w_242_106, w_215_170, w_166_331);
  nand2 I242_173(w_242_173, w_135_074, w_139_002);
  or2  I242_223(w_242_223, w_164_326, w_118_211);
  nand2 I243_003(w_243_003, w_005_518, w_016_362);
  and2 I243_013(w_243_013, w_064_433, w_164_186);
  or2  I243_075(w_243_075, w_043_053, w_140_219);
  or2  I243_109(w_243_109, w_080_022, w_166_294);
  or2  I243_141(w_243_141, w_186_198, w_191_037);
  and2 I243_147(w_243_147, w_137_202, w_087_147);
  or2  I243_152(w_243_152, w_018_076, w_016_125);
  nand2 I243_205(w_243_205, w_085_000, w_113_080);
  nand2 I243_223(w_243_223, w_059_209, w_082_217);
  nand2 I244_160(w_244_160, w_139_005, w_096_185);
  and2 I244_220(w_244_220, w_075_188, w_208_032);
  not1 I245_076(w_245_076, w_087_135);
  or2  I245_090(w_245_090, w_020_001, w_044_371);
  not1 I245_236(w_245_236, w_022_090);
  nand2 I245_277(w_245_277, w_201_698, w_018_079);
  or2  I245_297(w_245_297, w_082_222, w_050_037);
  and2 I246_002(w_246_002, w_236_410, w_126_251);
  and2 I246_107(w_246_107, w_227_012, w_172_405);
  not1 I246_253(w_246_253, w_011_251);
  not1 I246_274(w_246_274, w_012_174);
  and2 I246_276(w_246_276, w_031_224, w_212_109);
  nand2 I246_287(w_246_287, w_129_022, w_120_032);
  not1 I247_091(w_247_091, w_071_233);
  nand2 I247_092(w_247_092, w_174_857, w_232_032);
  not1 I247_496(w_247_496, w_229_295);
  or2  I247_498(w_247_498, w_064_534, w_165_550);
  or2  I247_610(w_247_610, w_198_578, w_010_077);
  or2  I247_611(w_247_611, w_189_115, w_191_211);
  or2  I248_014(w_248_014, w_230_032, w_086_776);
  nand2 I248_299(w_248_299, w_164_314, w_072_015);
  or2  I248_327(w_248_327, w_187_203, w_061_245);
  or2  I248_459(w_248_459, w_032_762, w_052_015);
  nand2 I248_648(w_248_648, w_029_125, w_199_751);
  and2 I249_036(w_249_036, w_047_062, w_170_220);
  nand2 I249_065(w_249_065, w_245_236, w_090_205);
  and2 I249_193(w_249_193, w_127_109, w_134_326);
  not1 I249_223(w_249_223, w_074_261);
  nand2 I249_255(w_249_255, w_088_500, w_158_643);
  or2  I250_003(w_250_003, w_204_342, w_134_010);
  nand2 I250_055(w_250_055, w_106_237, w_095_074);
  or2  I250_059(w_250_059, w_029_207, w_055_011);
  nand2 I250_068(w_250_068, w_186_442, w_095_094);
  nand2 I250_226(w_250_226, w_103_160, w_102_155);
  nand2 I250_287(w_250_287, w_197_838, w_194_089);
  nand2 I250_420(w_250_420, w_121_081, w_240_754);
  nand2 I250_445(w_250_445, w_239_174, w_055_055);
  not1 I251_026(w_251_026, w_056_299);
  not1 I251_031(w_251_031, w_036_166);
  or2  I251_208(w_251_208, w_026_383, w_085_051);
  or2  I251_229(w_251_229, w_180_005, w_013_005);
  nand2 I251_259(w_251_259, w_223_631, w_129_016);
  not1 I251_262(w_251_262, w_082_342);
  or2  I252_190(w_252_190, w_052_101, w_062_469);
  or2  I252_225(w_252_225, w_159_169, w_233_384);
  or2  I252_358(w_252_358, w_006_063, w_226_000);
  and2 I252_383(w_252_383, w_230_036, w_224_075);
  nand2 I253_000(w_253_000, w_195_256, w_118_217);
  not1 I253_003(w_253_003, w_080_104);
  and2 I253_005(w_253_005, w_106_438, w_243_013);
  or2  I253_009(w_253_009, w_223_582, w_165_140);
  or2  I253_031(w_253_031, w_163_120, w_028_854);
  and2 I253_032(w_253_032, w_184_243, w_187_096);
  nand2 I253_048(w_253_048, w_168_104, w_183_070);
  nand2 I254_057(w_254_057, w_045_018, w_075_100);
  and2 I254_184(w_254_184, w_043_040, w_105_044);
  or2  I254_269(w_254_269, w_239_054, w_033_751);
  not1 I254_306(w_254_306, w_187_131);
  not1 I255_000(w_255_000, w_230_246);
  not1 I255_003(w_255_003, w_231_083);
  not1 I255_007(w_255_007, w_058_085);
  nand2 I255_033(w_255_033, w_095_009, w_227_260);
  not1 I255_036(w_255_036, w_069_143);
  or2  I256_020(w_256_020, w_059_192, w_013_228);
  and2 I256_047(w_256_047, w_133_790, w_245_076);
  not1 I256_124(w_256_124, w_152_116);
  or2  I257_044(w_257_044, w_097_228, w_057_122);
  nand2 I257_146(w_257_146, w_181_388, w_113_299);
  and2 I257_271(w_257_271, w_194_268, w_151_283);
  or2  I257_402(w_257_402, w_152_395, w_171_369);
  or2  I257_428(w_257_428, w_046_327, w_024_180);
  not1 I257_512(w_257_512, w_104_062);
  or2  I257_562(w_257_562, w_127_071, w_033_471);
  and2 I258_122(w_258_122, w_095_112, w_045_534);
  and2 I258_236(w_258_236, w_162_154, w_067_649);
  not1 I258_754(w_258_754, w_055_615);
  not1 I259_099(w_259_099, w_044_047);
  not1 I259_167(w_259_167, w_252_190);
  and2 I259_234(w_259_234, w_058_190, w_034_032);
  not1 I259_308(w_259_308, w_180_172);
  not1 I259_372(w_259_372, w_184_085);
  or2  I259_461(w_259_461, w_102_563, w_080_031);
  and2 I259_505(w_259_505, w_075_101, w_043_029);
  nand2 I260_123(w_260_123, w_062_149, w_178_504);
  nand2 I260_154(w_260_154, w_213_041, w_243_223);
  not1 I260_373(w_260_373, w_187_153);
  and2 I260_510(w_260_510, w_236_154, w_077_108);
  not1 I260_578(w_260_578, w_186_007);
  not1 I260_616(w_260_616, w_123_027);
  not1 I260_751(w_260_751, w_163_095);
  not1 I260_812(w_260_812, w_251_031);
  nand2 I261_418(w_261_418, w_145_023, w_094_208);
  or2  I261_469(w_261_469, w_084_050, w_042_099);
  or2  I262_035(w_262_035, w_215_428, w_135_226);
  or2  I262_059(w_262_059, w_022_020, w_043_032);
  not1 I262_086(w_262_086, w_227_416);
  or2  I262_110(w_262_110, w_029_029, w_143_418);
  and2 I262_146(w_262_146, w_102_162, w_236_606);
  nand2 I263_069(w_263_069, w_230_238, w_100_642);
  nand2 I263_077(w_263_077, w_070_053, w_220_821);
  and2 I263_093(w_263_093, w_252_225, w_105_855);
  not1 I263_174(w_263_174, w_010_159);
  nand2 I263_189(w_263_189, w_257_562, w_172_060);
  or2  I263_199(w_263_199, w_092_043, w_023_170);
  and2 I264_132(w_264_132, w_211_029, w_095_002);
  or2  I264_371(w_264_371, w_020_003, w_095_149);
  or2  I264_439(w_264_439, w_128_217, w_171_333);
  nand2 I264_606(w_264_606, w_219_030, w_038_648);
  and2 I264_782(w_264_782, w_023_548, w_097_595);
  and2 I264_796(w_264_796, w_024_200, w_104_180);
  nand2 I264_900(w_264_900, w_151_282, w_010_522);
  nand2 I265_059(w_265_059, w_010_251, w_209_179);
  and2 I265_060(w_265_060, w_039_037, w_174_453);
  nand2 I265_065(w_265_065, w_160_599, w_086_408);
  not1 I265_068(w_265_068, w_171_264);
  or2  I265_075(w_265_075, w_230_251, w_185_103);
  and2 I265_202(w_265_202, w_121_260, w_068_018);
  or2  I265_414(w_265_414, w_204_257, w_088_077);
  nand2 I265_528(w_265_528, w_077_240, w_007_431);
  nand2 I266_295(w_266_295, w_177_347, w_115_025);
  nand2 I266_429(w_266_429, w_044_273, w_083_068);
  and2 I266_451(w_266_451, w_160_155, w_056_096);
  nand2 I267_076(w_267_076, w_244_220, w_083_249);
  and2 I267_088(w_267_088, w_162_133, w_105_397);
  and2 I267_111(w_267_111, w_086_017, w_000_848);
  or2  I267_141(w_267_141, w_113_167, w_008_034);
  not1 I267_225(w_267_225, w_243_152);
  nand2 I267_550(w_267_550, w_110_051, w_028_376);
  not1 I267_602(w_267_602, w_186_304);
  or2  I268_116(w_268_116, w_260_373, w_126_304);
  nand2 I268_172(w_268_172, w_087_195, w_193_252);
  or2  I268_353(w_268_353, w_047_164, w_074_479);
  and2 I268_446(w_268_446, w_083_253, w_086_750);
  not1 I269_017(w_269_017, w_084_494);
  and2 I269_031(w_269_031, w_147_520, w_214_027);
  not1 I269_035(w_269_035, w_166_269);
  not1 I270_103(w_270_103, w_137_643);
  not1 I270_166(w_270_166, w_267_602);
  nand2 I270_174(w_270_174, w_050_289, w_149_232);
  and2 I270_473(w_270_473, w_265_060, w_036_095);
  nand2 I270_681(w_270_681, w_020_010, w_074_588);
  or2  I271_002(w_271_002, w_142_340, w_238_360);
  or2  I271_038(w_271_038, w_249_223, w_118_258);
  nand2 I271_039(w_271_039, w_139_002, w_000_075);
  nand2 I271_074(w_271_074, w_267_141, w_207_104);
  nand2 I271_107(w_271_107, w_171_296, w_120_005);
  and2 I271_157(w_271_157, w_010_220, w_107_127);
  and2 I272_135(w_272_135, w_270_473, w_144_394);
  or2  I273_061(w_273_061, w_215_322, w_159_062);
  and2 I273_127(w_273_127, w_021_131, w_109_178);
  not1 I273_366(w_273_366, w_039_023);
  nand2 I274_000(w_274_000, w_193_669, w_008_892);
  and2 I274_002(w_274_002, w_022_161, w_119_051);
  not1 I275_000(w_275_000, w_057_091);
  not1 I275_002(w_275_002, w_228_267);
  not1 I275_003(w_275_003, w_174_269);
  nand2 I276_645(w_276_645, w_248_459, w_106_224);
  or2  I276_686(w_276_686, w_240_011, w_002_194);
  and2 I277_033(w_277_033, w_249_193, w_177_912);
  not1 I277_088(w_277_088, w_122_348);
  nand2 I277_106(w_277_106, w_087_080, w_154_137);
  or2  I277_109(w_277_109, w_006_012, w_113_515);
  or2  I278_065(w_278_065, w_264_900, w_150_122);
  and2 I278_216(w_278_216, w_198_330, w_268_116);
  not1 I278_224(w_278_224, w_119_080);
  or2  I278_359(w_278_359, w_256_020, w_062_440);
  or2  I278_442(w_278_442, w_091_186, w_031_027);
  or2  I279_032(w_279_032, w_026_275, w_219_038);
  nand2 I279_088(w_279_088, w_057_157, w_094_011);
  or2  I279_344(w_279_344, w_253_032, w_180_050);
  and2 I280_002(w_280_002, w_250_226, w_146_224);
  or2  I280_016(w_280_016, w_102_233, w_253_031);
  nand2 I280_018(w_280_018, w_055_503, w_217_279);
  nand2 I280_019(w_280_019, w_185_100, w_206_057);
  and2 I280_023(w_280_023, w_019_360, w_210_574);
  not1 I281_029(w_281_029, w_078_087);
  or2  I281_115(w_281_115, w_117_105, w_060_057);
  not1 I281_197(w_281_197, w_211_052);
  and2 I281_344(w_281_344, w_090_048, w_195_070);
  and2 I281_706(w_281_706, w_182_223, w_051_184);
  and2 I282_074(w_282_074, w_145_046, w_057_190);
  or2  I282_103(w_282_103, w_117_263, w_025_087);
  not1 I283_079(w_283_079, w_093_791);
  nand2 I283_250(w_283_250, w_119_299, w_074_342);
  not1 I283_283(w_283_283, w_065_363);
  nand2 I283_335(w_283_335, w_170_166, w_008_384);
  and2 I283_355(w_283_355, w_143_159, w_009_006);
  or2  I283_373(w_283_373, w_093_320, w_132_192);
  nand2 I283_498(w_283_498, w_153_177, w_012_373);
  and2 I284_079(w_284_079, w_197_896, w_278_359);
  or2  I284_092(w_284_092, w_175_828, w_203_312);
  nand2 I284_102(w_284_102, w_035_015, w_042_078);
  not1 I284_229(w_284_229, w_195_348);
  not1 I284_312(w_284_312, w_058_233);
  or2  I284_405(w_284_405, w_067_283, w_077_012);
  not1 I284_430(w_284_430, w_061_172);
  and2 I284_462(w_284_462, w_137_394, w_046_052);
  not1 I285_102(w_285_102, w_090_079);
  and2 I285_158(w_285_158, w_012_218, w_211_528);
  or2  I286_249(w_286_249, w_106_008, w_268_446);
  not1 I287_109(w_287_109, w_144_234);
  nand2 I287_110(w_287_110, w_197_674, w_082_301);
  not1 I287_395(w_287_395, w_241_142);
  nand2 I287_695(w_287_695, w_053_645, w_070_888);
  nand2 I288_135(w_288_135, w_147_269, w_092_138);
  and2 I288_203(w_288_203, w_072_006, w_114_283);
  nand2 I288_353(w_288_353, w_214_092, w_052_125);
  nand2 I288_665(w_288_665, w_151_255, w_015_406);
  not1 I289_304(w_289_304, w_003_052);
  or2  I289_480(w_289_480, w_188_491, w_049_190);
  or2  I289_855(w_289_855, w_035_397, w_180_305);
  or2  I290_052(w_290_052, w_242_173, w_074_847);
  and2 I290_115(w_290_115, w_024_171, w_009_055);
  and2 I290_183(w_290_183, w_023_089, w_250_068);
  or2  I290_260(w_290_260, w_186_001, w_055_607);
  and2 I291_035(w_291_035, w_190_222, w_118_384);
  or2  I291_052(w_291_052, w_282_074, w_015_226);
  nand2 I291_707(w_291_707, w_290_183, w_214_052);
  and2 I292_109(w_292_109, w_164_155, w_207_236);
  and2 I292_160(w_292_160, w_018_177, w_260_123);
  and2 I292_235(w_292_235, w_278_442, w_193_418);
  or2  I292_413(w_292_413, w_274_002, w_110_010);
  or2  I292_704(w_292_706, w_179_549, w_292_705);
  nand2 I292_705(w_292_707, w_080_103, w_292_706);
  not1 I292_706(w_292_708, w_292_707);
  not1 I292_707(w_292_709, w_292_708);
  not1 I292_708(w_292_710, w_292_709);
  and2 I292_709(w_292_711, w_292_710, w_126_166);
  not1 I292_710(w_292_712, w_292_711);
  and2 I292_711(w_292_713, w_284_092, w_292_712);
  not1 I292_712(w_292_714, w_292_713);
  or2  I292_713(w_292_705, w_292_714, w_029_016);
  or2  I293_051(w_293_051, w_145_050, w_281_029);
  not1 I293_087(w_293_087, w_191_118);
  and2 I293_573(w_293_573, w_064_789, w_142_208);
  or2  I293_625(w_293_625, w_139_013, w_250_420);
  not1 I293_697(w_293_697, w_023_186);
  and2 I294_010(w_294_010, w_262_059, w_006_141);
  nand2 I294_038(w_294_038, w_049_602, w_219_277);
  or2  I294_279(w_294_279, w_104_169, w_111_101);
  not1 I294_644(w_294_644, w_031_399);
  and2 I294_710(w_294_710, w_197_422, w_227_067);
  or2  I295_009(w_295_009, w_100_305, w_051_438);
  or2  I295_080(w_295_080, w_186_070, w_267_076);
  nand2 I295_116(w_295_116, w_063_064, w_178_600);
  nand2 I295_170(w_295_170, w_227_522, w_182_115);
  and2 I296_000(w_296_000, w_146_073, w_150_160);
  or2  I296_017(w_296_017, w_001_570, w_024_070);
  nand2 I296_067(w_296_067, w_243_075, w_233_078);
  and2 I297_114(w_297_114, w_292_235, w_180_333);
  nand2 I297_117(w_297_117, w_032_588, w_101_120);
  and2 I297_138(w_297_138, w_283_335, w_171_472);
  not1 I297_150(w_297_150, w_243_141);
  not1 I297_196(w_297_196, w_146_328);
  or2  I298_205(w_298_205, w_194_909, w_059_169);
  or2  I299_079(w_299_079, w_086_059, w_059_177);
  or2  I299_134(w_299_134, w_048_050, w_029_110);
  and2 I300_036(w_300_036, w_297_138, w_145_029);
  and2 I300_208(w_300_208, w_287_395, w_010_086);
  or2  I300_507(w_300_507, w_246_002, w_130_925);
  or2  I300_631(w_300_631, w_098_222, w_201_514);
  and2 I300_854(w_300_854, w_259_234, w_050_311);
  not1 I301_070(w_301_070, w_044_159);
  nand2 I301_356(w_301_356, w_252_383, w_091_145);
  and2 I301_478(w_301_478, w_257_271, w_071_363);
  or2  I302_000(w_302_000, w_257_402, w_211_040);
  nand2 I302_016(w_302_016, w_246_287, w_136_307);
  and2 I302_020(w_302_020, w_019_417, w_291_707);
  not1 I302_023(w_302_023, w_214_107);
  or2  I302_029(w_302_029, w_068_212, w_276_645);
  not1 I304_041(w_304_041, w_207_244);
  not1 I304_046(w_304_046, w_270_681);
  or2  I304_064(w_304_064, w_296_000, w_076_616);
  nand2 I304_079(w_304_079, w_224_041, w_297_114);
  not1 I305_009(w_305_009, w_173_110);
  or2  I305_046(w_305_046, w_140_308, w_152_479);
  not1 I305_083(w_305_083, w_123_025);
  or2  I305_091(w_305_091, w_190_289, w_064_448);
  not1 I305_093(w_305_093, w_164_129);
  not1 I305_097(w_305_097, w_116_007);
  or2  I305_151(w_305_151, w_001_397, w_264_439);
  nand2 I306_015(w_306_015, w_138_145, w_032_424);
  not1 I306_018(w_306_018, w_038_101);
  nand2 I306_028(w_306_028, w_112_071, w_104_159);
  nand2 I306_072(w_306_072, w_098_257, w_201_076);
  not1 I306_088(w_306_088, w_146_170);
  not1 I306_091(w_306_091, w_221_070);
  or2  I306_137(w_306_137, w_250_059, w_295_116);
  not1 I307_312(w_307_312, w_052_108);
  not1 I308_061(w_308_061, w_026_430);
  nand2 I308_084(w_308_084, w_252_358, w_263_093);
  or2  I309_002(w_309_002, w_191_174, w_079_000);
  or2  I309_115(w_309_115, w_109_169, w_143_549);
  or2  I309_151(w_309_151, w_097_260, w_113_070);
  or2  I309_164(w_309_164, w_263_189, w_265_528);
  not1 I309_193(w_309_193, w_048_161);
  or2  I310_259(w_310_259, w_075_179, w_181_234);
  not1 I311_140(w_311_140, w_051_317);
  or2  I311_169(w_311_169, w_011_032, w_131_632);
  nand2 I312_051(w_312_051, w_016_328, w_094_078);
  and2 I312_791(w_312_791, w_026_029, w_134_203);
  and2 I312_894(w_312_894, w_116_038, w_146_129);
  or2  I313_027(w_313_027, w_144_282, w_031_089);
  nand2 I313_166(w_313_166, w_024_402, w_297_150);
  and2 I313_170(w_313_170, w_156_302, w_226_005);
  not1 I313_228(w_313_228, w_038_448);
  not1 I313_246(w_313_246, w_054_102);
  not1 I313_446(w_313_446, w_034_127);
  nand2 I313_477(w_313_477, w_253_003, w_134_097);
  and2 I314_086(w_314_086, w_114_356, w_014_453);
  nand2 I314_388(w_314_388, w_255_033, w_123_048);
  nand2 I314_765(w_314_765, w_014_086, w_231_057);
  not1 I315_105(w_315_105, w_123_160);
  and2 I315_129(w_315_129, w_291_052, w_188_161);
  not1 I315_455(w_315_455, w_140_630);
  and2 I315_491(w_315_491, w_006_073, w_184_157);
  nand2 I316_056(w_316_056, w_012_086, w_005_191);
  nand2 I316_137(w_316_137, w_152_696, w_143_356);
  nand2 I316_320(w_316_320, w_139_007, w_247_498);
  nand2 I316_635(w_316_635, w_219_217, w_158_145);
  and2 I316_731(w_316_731, w_145_097, w_060_178);
  nand2 I316_851(w_316_853, w_191_036, w_316_852);
  and2 I316_852(w_316_854, w_316_853, w_314_388);
  not1 I316_853(w_316_855, w_316_854);
  or2  I316_854(w_316_856, w_316_855, w_145_091);
  or2  I316_855(w_316_857, w_316_856, w_049_250);
  not1 I316_856(w_316_858, w_316_857);
  and2 I316_857(w_316_859, w_316_858, w_117_290);
  and2 I316_858(w_316_860, w_316_859, w_060_242);
  not1 I316_859(w_316_861, w_316_860);
  not1 I316_860(w_316_862, w_316_861);
  and2 I316_861(w_316_852, w_158_198, w_316_862);
  and2 I317_043(w_317_043, w_238_053, w_271_157);
  or2  I317_059(w_317_059, w_110_581, w_067_229);
  or2  I317_533(w_317_533, w_192_002, w_074_254);
  and2 I317_562(w_317_562, w_013_042, w_312_791);
  not1 I317_740(w_317_740, w_038_168);
  and2 I318_024(w_318_024, w_216_129, w_037_013);
  not1 I318_026(w_318_026, w_297_196);
  not1 I318_031(w_318_031, w_211_276);
  nand2 I318_038(w_318_038, w_041_014, w_182_274);
  not1 I318_051(w_318_051, w_177_095);
  or2  I318_062(w_318_064, w_318_063, w_260_510);
  not1 I318_063(w_318_065, w_318_064);
  nand2 I318_064(w_318_066, w_138_183, w_318_065);
  not1 I318_065(w_318_067, w_318_066);
  not1 I318_066(w_318_068, w_318_067);
  and2 I318_067(w_318_069, w_004_009, w_318_068);
  and2 I318_068(w_318_070, w_119_119, w_318_069);
  nand2 I318_069(w_318_071, w_318_070, w_026_387);
  not1 I318_070(w_318_072, w_318_071);
  not1 I318_071(w_318_063, w_318_072);
  not1 I319_072(w_319_072, w_074_963);
  or2  I319_254(w_319_254, w_130_917, w_027_437);
  not1 I320_029(w_320_029, w_040_338);
  and2 I320_101(w_320_101, w_106_418, w_159_192);
  or2  I320_365(w_320_365, w_099_038, w_017_016);
  and2 I320_609(w_320_609, w_200_683, w_016_461);
  not1 I321_011(w_321_011, w_141_078);
  and2 I321_277(w_321_277, w_233_342, w_049_649);
  nand2 I321_543(w_321_543, w_144_128, w_065_527);
  or2  I321_763(w_321_763, w_305_151, w_195_335);
  or2  I322_585(w_322_585, w_248_299, w_194_011);
  not1 I323_219(w_323_219, w_050_264);
  and2 I323_372(w_323_372, w_019_314, w_271_002);
  and2 I323_678(w_323_678, w_271_107, w_186_544);
  not1 I323_902(w_323_902, w_255_007);
  nand2 I324_020(w_324_020, w_023_106, w_250_445);
  and2 I324_030(w_324_030, w_172_388, w_267_550);
  nand2 I324_151(w_324_151, w_203_110, w_049_654);
  nand2 I324_589(w_324_589, w_246_276, w_223_840);
  not1 I325_027(w_325_027, w_270_174);
  or2  I325_156(w_325_156, w_289_480, w_236_315);
  not1 I325_265(w_325_265, w_000_958);
  nand2 I326_011(w_326_011, w_224_058, w_064_668);
  nand2 I326_193(w_326_193, w_061_410, w_059_230);
  or2  I327_007(w_327_007, w_238_389, w_072_020);
  or2  I327_025(w_327_025, w_115_019, w_250_055);
  not1 I327_728(w_327_728, w_120_035);
  not1 I327_873(w_327_873, w_146_065);
  or2  I328_273(w_328_273, w_293_087, w_090_209);
  nand2 I329_037(w_329_037, w_038_135, w_107_190);
  and2 I329_379(w_329_379, w_324_020, w_049_003);
  or2  I329_502(w_329_502, w_315_455, w_323_219);
  or2  I330_072(w_330_072, w_188_427, w_077_266);
  or2  I330_107(w_330_107, w_131_682, w_072_003);
  nand2 I330_151(w_330_151, w_110_005, w_052_145);
  nand2 I331_007(w_331_007, w_102_094, w_311_140);
  and2 I331_050(w_331_050, w_149_065, w_281_706);
  nand2 I331_087(w_331_087, w_080_114, w_250_003);
  nand2 I331_095(w_331_095, w_007_307, w_096_255);
  nand2 I332_075(w_332_075, w_307_312, w_187_022);
  nand2 I332_147(w_332_147, w_284_312, w_294_710);
  nand2 I332_161(w_332_161, w_325_156, w_150_154);
  not1 I332_184(w_332_184, w_271_074);
  not1 I332_407(w_332_407, w_198_741);
  not1 I333_108(w_333_108, w_182_228);
  and2 I333_374(w_333_374, w_284_462, w_139_012);
  nand2 I333_540(w_333_540, w_162_466, w_316_056);
  or2  I334_000(w_334_000, w_231_026, w_217_819);
  nand2 I334_002(w_334_002, w_176_180, w_121_485);
  nand2 I335_094(w_335_094, w_195_029, w_262_035);
  not1 I335_105(w_335_105, w_038_560);
  nand2 I336_047(w_336_047, w_020_008, w_276_686);
  not1 I336_056(w_336_056, w_323_372);
  nand2 I338_448(w_338_448, w_297_117, w_176_154);
  not1 I338_783(w_338_783, w_261_469);
  not1 I339_117(w_339_117, w_064_610);
  and2 I340_120(w_340_120, w_001_277, w_069_146);
  and2 I340_224(w_340_224, w_120_068, w_197_352);
  and2 I340_315(w_340_315, w_230_295, w_118_102);
  and2 I340_328(w_340_328, w_194_219, w_106_016);
  not1 I341_018(w_341_018, w_057_010);
  not1 I341_025(w_341_025, w_162_427);
  nand2 I341_044(w_341_044, w_108_000, w_306_088);
  and2 I341_045(w_341_045, w_182_193, w_010_044);
  nand2 I341_046(w_341_046, w_294_010, w_319_254);
  not1 I342_109(w_342_109, w_077_491);
  not1 I342_140(w_342_140, w_091_182);
  or2  I342_172(w_342_172, w_251_229, w_260_751);
  or2  I342_504(w_342_504, w_305_097, w_133_266);
  nand2 I343_076(w_343_076, w_139_006, w_009_042);
  not1 I343_160(w_343_160, w_019_152);
  not1 I343_172(w_343_172, w_084_131);
  not1 I344_000(w_344_000, w_259_308);
  not1 I344_001(w_344_001, w_192_002);
  and2 I345_197(w_345_197, w_009_002, w_254_057);
  or2  I346_012(w_346_012, w_151_000, w_058_071);
  or2  I346_022(w_346_022, w_142_567, w_166_360);
  nand2 I346_024(w_346_024, w_342_172, w_056_039);
  or2  I346_038(w_346_038, w_151_298, w_305_091);
  nand2 I347_123(w_347_123, w_068_283, w_080_092);
  or2  I347_130(w_347_130, w_006_162, w_018_054);
  or2  I348_000(w_348_000, w_263_174, w_302_000);
  not1 I349_067(w_349_067, w_117_196);
  and2 I349_088(w_349_088, w_071_366, w_275_003);
  or2  I350_011(w_350_011, w_190_000, w_156_456);
  nand2 I350_226(w_350_226, w_208_267, w_027_712);
  not1 I351_002(w_351_002, w_195_082);
  and2 I351_004(w_351_004, w_299_079, w_277_109);
  or2  I351_041(w_351_041, w_081_041, w_231_049);
  nand2 I351_044(w_351_044, w_331_095, w_227_547);
  and2 I351_045(w_351_045, w_070_154, w_127_077);
  or2  I352_075(w_352_075, w_348_000, w_037_128);
  nand2 I352_100(w_352_100, w_003_084, w_120_110);
  and2 I353_055(w_353_055, w_267_088, w_013_011);
  not1 I353_057(w_353_057, w_189_298);
  or2  I353_080(w_353_080, w_153_415, w_177_030);
  and2 I353_088(w_353_088, w_083_137, w_336_056);
  and2 I353_102(w_353_102, w_024_040, w_326_193);
  nand2 I354_345(w_354_345, w_016_122, w_151_109);
  or2  I354_649(w_354_649, w_280_023, w_316_320);
  and2 I355_160(w_355_160, w_030_246, w_000_868);
  not1 I356_012(w_356_012, w_125_089);
  and2 I356_475(w_356_475, w_295_170, w_354_649);
  or2  I356_701(w_356_701, w_044_198, w_192_002);
  not1 I356_756(w_356_756, w_038_037);
  or2  I357_147(w_357_147, w_194_471, w_127_130);
  and2 I358_031(w_358_031, w_289_304, w_238_159);
  or2  I358_421(w_358_421, w_341_044, w_074_297);
  not1 I358_438(w_358_438, w_041_122);
  not1 I358_607(w_358_607, w_267_111);
  nand2 I358_750(w_358_750, w_083_302, w_059_264);
  or2  I359_460(w_359_460, w_216_126, w_039_310);
  nand2 I360_035(w_360_035, w_058_009, w_045_076);
  and2 I361_000(w_361_000, w_321_277, w_047_327);
  or2  I361_026(w_361_026, w_306_028, w_185_277);
  nand2 I361_029(w_361_029, w_262_086, w_321_543);
  or2  I361_032(w_361_032, w_212_013, w_017_020);
  nand2 I361_059(w_361_059, w_215_267, w_285_158);
  or2  I362_019(w_362_019, w_083_619, w_107_046);
  nand2 I362_069(w_362_069, w_277_033, w_144_347);
  and2 I362_083(w_362_083, w_068_039, w_265_075);
  and2 I363_006(w_363_006, w_306_015, w_089_113);
  and2 I364_383(w_364_383, w_013_121, w_102_298);
  not1 I364_803(w_364_803, w_234_554);
  or2  I365_043(w_365_043, w_264_371, w_214_005);
  not1 I365_069(w_365_069, w_184_039);
  not1 I365_145(w_365_145, w_321_011);
  not1 I366_160(w_366_160, w_075_114);
  not1 I366_444(w_366_444, w_141_707);
  and2 I367_053(w_367_053, w_233_391, w_167_275);
  and2 I367_133(w_367_133, w_024_112, w_049_739);
  or2  I367_180(w_367_180, w_014_354, w_247_496);
  nand2 I367_243(w_367_243, w_284_430, w_366_160);
  nand2 I368_005(w_368_005, w_046_179, w_057_121);
  nand2 I368_006(w_368_006, w_027_584, w_223_925);
  not1 I369_005(w_369_005, w_230_048);
  or2  I369_081(w_369_081, w_356_012, w_162_210);
  and2 I369_305(w_369_305, w_309_002, w_338_783);
  not1 I370_154(w_370_154, w_178_016);
  not1 I371_053(w_371_053, w_247_610);
  and2 I372_378(w_372_378, w_275_000, w_362_069);
  nand2 I372_442(w_372_442, w_248_648, w_128_216);
  not1 I372_455(w_372_455, w_278_224);
  and2 I373_024(w_373_024, w_332_407, w_351_045);
  or2  I373_069(w_373_069, w_368_005, w_284_102);
  or2  I374_011(w_374_011, w_312_894, w_237_379);
  and2 I374_012(w_374_012, w_021_051, w_232_363);
  nand2 I375_045(w_375_045, w_022_177, w_007_333);
  not1 I376_277(w_376_277, w_141_342);
  and2 I376_391(w_376_391, w_068_303, w_166_015);
  and2 I377_168(w_377_168, w_278_216, w_261_418);
  not1 I377_284(w_377_284, w_190_348);
  or2  I377_395(w_377_395, w_096_380, w_329_037);
  not1 I377_418(w_377_418, w_224_042);
  or2  I378_247(w_378_247, w_245_090, w_319_072);
  nand2 I379_001(w_379_001, w_332_147, w_194_211);
  not1 I379_050(w_379_050, w_299_134);
  or2  I379_060(w_379_060, w_254_269, w_187_022);
  or2  I380_030(w_380_030, w_053_816, w_145_062);
  nand2 I380_104(w_380_104, w_347_130, w_351_044);
  and2 I380_107(w_380_107, w_296_067, w_377_395);
  nand2 I380_238(w_380_238, w_230_082, w_175_456);
  or2  I381_222(w_381_222, w_082_015, w_101_083);
  and2 I381_632(w_381_632, w_173_043, w_096_229);
  or2  I382_232(w_382_232, w_259_099, w_020_077);
  nand2 I382_405(w_382_405, w_128_201, w_233_128);
  and2 I382_610(w_382_610, w_241_336, w_249_255);
  and2 I383_005(w_383_005, w_021_230, w_241_276);
  or2  I383_095(w_383_095, w_313_477, w_151_196);
  or2  I383_156(w_383_156, w_218_004, w_304_046);
  not1 I383_337(w_383_337, w_379_060);
  not1 I383_420(w_383_420, w_147_152);
  or2  I385_375(w_385_375, w_028_895, w_135_006);
  or2  I386_036(w_386_036, w_041_070, w_013_058);
  not1 I386_195(w_386_195, w_046_393);
  nand2 I386_630(w_386_630, w_021_186, w_201_655);
  and2 I387_049(w_387_049, w_061_432, w_138_738);
  and2 I388_023(w_388_023, w_104_246, w_122_472);
  and2 I388_079(w_388_079, w_169_022, w_224_009);
  not1 I388_098(w_388_098, w_320_365);
  or2  I388_100(w_388_100, w_361_026, w_290_115);
  not1 I388_223(w_388_223, w_181_495);
  not1 I388_244(w_388_244, w_071_329);
  nand2 I389_061(w_389_061, w_275_000, w_232_202);
  or2  I389_068(w_389_068, w_263_069, w_206_126);
  not1 I389_092(w_389_092, w_116_038);
  or2  I389_335(w_389_335, w_353_102, w_177_395);
  nand2 I390_033(w_390_033, w_203_082, w_356_475);
  nand2 I391_028(w_391_028, w_185_078, w_035_009);
  not1 I392_000(w_392_000, w_167_458);
  or2  I393_163(w_393_163, w_388_223, w_003_067);
  and2 I393_323(w_393_323, w_255_003, w_159_064);
  nand2 I394_103(w_394_103, w_073_156, w_308_084);
  nand2 I394_118(w_394_118, w_331_050, w_230_252);
  nand2 I394_129(w_394_129, w_152_621, w_345_197);
  nand2 I394_195(w_394_195, w_347_123, w_224_038);
  or2  I395_026(w_395_026, w_342_504, w_332_184);
  and2 I395_081(w_395_081, w_381_222, w_394_118);
  or2  I395_103(w_395_103, w_045_560, w_221_136);
  or2  I395_161(w_395_161, w_085_044, w_216_050);
  or2  I396_533(w_396_533, w_389_068, w_135_221);
  nand2 I397_098(w_397_098, w_260_616, w_285_102);
  or2  I397_194(w_397_194, w_162_244, w_238_251);
  and2 I397_197(w_397_197, w_018_076, w_311_169);
  and2 I397_322(w_397_322, w_389_061, w_248_327);
  nand2 I398_362(w_398_362, w_144_323, w_187_011);
  nand2 I399_008(w_399_008, w_190_237, w_196_712);
  or2  I399_050(w_399_050, w_259_505, w_309_115);
  and2 I399_061(w_399_061, w_062_371, w_220_257);
  not1 I399_064(w_399_064, w_039_232);
  and2 I399_091(w_399_091, w_344_000, w_294_644);
  nand2 I400_025(w_400_025, w_217_372, w_094_817);
  or2  I400_203(w_400_203, w_132_300, w_183_041);
  or2  I400_789(w_400_791, w_174_538, w_400_790);
  and2 I400_790(w_400_792, w_400_791, w_310_259);
  or2  I400_791(w_400_793, w_400_792, w_353_055);
  not1 I400_792(w_400_794, w_400_793);
  nand2 I400_793(w_400_795, w_166_219, w_400_794);
  nand2 I400_794(w_400_796, w_150_140, w_400_795);
  not1 I400_795(w_400_797, w_400_796);
  nand2 I400_796(w_400_798, w_400_797, w_394_195);
  not1 I400_797(w_400_790, w_400_798);
  or2  I401_500(w_401_500, w_369_305, w_178_590);
  not1 I401_636(w_401_636, w_238_033);
  not1 I401_729(w_401_729, w_196_045);
  nand2 I401_785(w_401_785, w_188_430, w_193_340);
  nand2 I402_188(w_402_188, w_259_372, w_322_585);
  or2  I402_217(w_402_217, w_387_049, w_038_591);
  not1 I403_085(w_403_085, w_129_004);
  nand2 I403_140(w_403_140, w_171_359, w_058_072);
  not1 I403_276(w_403_276, w_245_297);
  and2 I403_277(w_403_277, w_374_011, w_038_118);
  and2 I403_278(w_403_278, w_280_019, w_008_428);
  or2  I404_022(w_404_022, w_358_607, w_147_213);
  nand2 I404_049(w_404_049, w_270_166, w_386_036);
  not1 I405_131(w_405_131, w_236_151);
  not1 I405_146(w_405_146, w_171_042);
  and2 I405_393(w_405_393, w_302_016, w_277_088);
  not1 I405_439(w_405_439, w_087_263);
  and2 I405_808(w_405_808, w_305_083, w_271_038);
  nand2 I406_013(w_406_013, w_351_002, w_273_366);
  and2 I406_047(w_406_047, w_264_132, w_043_015);
  not1 I406_263(w_406_263, w_404_022);
  and2 I406_437(w_406_437, w_316_635, w_036_040);
  not1 I406_577(w_406_577, w_094_726);
  or2  I407_039(w_407_039, w_338_448, w_132_367);
  not1 I407_066(w_407_066, w_139_007);
  not1 I408_011(w_408_011, w_107_180);
  and2 I408_090(w_408_090, w_388_079, w_023_594);
  not1 I410_001(w_410_001, w_237_228);
  or2  I410_093(w_410_093, w_174_516, w_376_277);
  or2  I411_948(w_411_948, w_260_154, w_312_051);
  or2  I412_106(w_412_106, w_174_762, w_230_248);
  not1 I412_147(w_412_147, w_228_637);
  or2  I412_746(w_412_746, w_246_253, w_282_103);
  not1 I413_287(w_413_287, w_195_487);
  or2  I413_446(w_413_446, w_163_181, w_006_157);
  not1 I414_008(w_414_008, w_255_036);
  not1 I414_153(w_414_153, w_193_416);
  or2  I414_162(w_414_162, w_131_070, w_130_262);
  and2 I415_059(w_415_059, w_192_001, w_055_688);
  and2 I415_247(w_415_247, w_177_524, w_243_205);
  not1 I415_370(w_415_370, w_329_379);
  not1 I416_134(w_416_134, w_162_396);
  or2  I416_301(w_416_301, w_117_148, w_364_803);
  nand2 I416_719(w_416_719, w_300_507, w_235_019);
  not1 I416_775(w_416_777, w_416_776);
  and2 I416_776(w_416_778, w_330_107, w_416_777);
  and2 I416_777(w_416_779, w_395_081, w_416_778);
  or2  I416_778(w_416_780, w_416_779, w_247_091);
  nand2 I416_779(w_416_781, w_346_012, w_416_780);
  and2 I416_780(w_416_776, w_416_781, w_298_205);
  nand2 I417_005(w_417_005, w_366_444, w_053_551);
  and2 I417_149(w_417_149, w_341_045, w_115_030);
  nand2 I417_156(w_417_156, w_293_051, w_358_750);
  and2 I418_005(w_418_005, w_365_043, w_393_163);
  or2  I418_034(w_418_034, w_122_366, w_103_825);
  not1 I420_527(w_420_527, w_233_319);
  or2  I421_003(w_421_003, w_063_198, w_203_304);
  and2 I421_146(w_421_146, w_321_763, w_020_024);
  and2 I421_159(w_421_159, w_333_108, w_324_151);
  nand2 I422_026(w_422_026, w_067_746, w_066_475);
  nand2 I422_041(w_422_041, w_227_408, w_414_162);
  and2 I423_027(w_423_027, w_317_740, w_246_107);
  nand2 I423_151(w_423_151, w_316_137, w_218_141);
  or2  I423_235(w_423_235, w_306_018, w_329_502);
  nand2 I424_038(w_424_038, w_149_161, w_418_005);
  and2 I424_083(w_424_083, w_083_164, w_192_000);
  and2 I424_336(w_424_336, w_288_203, w_078_211);
  or2  I424_509(w_424_509, w_043_038, w_100_172);
  or2  I427_082(w_427_082, w_162_321, w_009_017);
  nand2 I427_096(w_427_096, w_236_162, w_084_062);
  nand2 I427_358(w_427_358, w_318_031, w_097_183);
  and2 I428_557(w_428_557, w_405_131, w_047_066);
  and2 I428_765(w_428_765, w_304_041, w_061_267);
  nand2 I429_111(w_429_111, w_026_361, w_253_009);
  nand2 I429_135(w_429_135, w_109_130, w_179_724);
  and2 I429_153(w_429_153, w_352_075, w_376_391);
  or2  I429_244(w_429_244, w_207_005, w_098_410);
  not1 I430_279(w_430_279, w_281_197);
  and2 I431_019(w_431_019, w_127_076, w_179_218);
  or2  I431_024(w_431_024, w_383_156, w_149_069);
  nand2 I431_025(w_431_025, w_429_244, w_258_122);
  nand2 I432_022(w_432_022, w_088_534, w_332_161);
  nand2 I432_026(w_432_026, w_340_224, w_255_000);
  and2 I433_066(w_433_066, w_218_016, w_149_239);
  or2  I433_391(w_433_391, w_102_611, w_363_006);
  or2  I435_077(w_435_077, w_044_051, w_326_011);
  and2 I435_087(w_435_087, w_107_021, w_197_746);
  nand2 I435_090(w_435_090, w_427_358, w_101_133);
  and2 I436_087(w_436_087, w_085_057, w_305_046);
  or2  I436_096(w_436_096, w_202_003, w_380_238);
  not1 I436_111(w_436_111, w_018_177);
  nand2 I437_005(w_437_005, w_004_023, w_294_038);
  or2  I437_050(w_437_050, w_379_050, w_003_057);
  nand2 I437_069(w_437_069, w_034_422, w_313_246);
  or2  I438_352(w_438_352, w_018_092, w_079_121);
  and2 I439_237(w_439_237, w_400_025, w_416_134);
  not1 I440_157(w_440_157, w_340_328);
  nand2 I440_458(w_440_458, w_243_003, w_171_215);
  or2  I440_479(w_440_479, w_272_135, w_212_084);
  not1 I440_495(w_440_495, w_178_351);
  nand2 I441_004(w_441_004, w_142_087, w_231_002);
  and2 I441_011(w_441_011, w_364_383, w_168_767);
  nand2 I441_013(w_441_013, w_091_552, w_023_188);
  or2  I442_003(w_442_003, w_225_026, w_250_287);
  and2 I442_014(w_442_014, w_044_107, w_399_061);
  nand2 I442_020(w_442_020, w_367_180, w_408_090);
  not1 I442_053(w_442_053, w_424_336);
  not1 I442_089(w_442_089, w_327_025);
  and2 I444_000(w_444_000, w_191_385, w_172_315);
  or2  I444_005(w_444_005, w_408_011, w_229_274);
  not1 I444_007(w_444_007, w_013_002);
  or2  I445_010(w_445_010, w_232_146, w_273_127);
  and2 I445_017(w_445_017, w_269_035, w_128_239);
  or2  I445_024(w_445_024, w_383_420, w_386_630);
  nand2 I445_037(w_445_037, w_019_116, w_026_311);
  or2  I446_650(w_446_650, w_279_032, w_248_014);
  nand2 I447_210(w_447_210, w_390_033, w_218_582);
  not1 I447_349(w_447_349, w_085_056);
  or2  I447_499(w_447_499, w_132_166, w_157_539);
  not1 I449_078(w_449_078, w_417_149);
  not1 I449_110(w_449_110, w_268_172);
  not1 I450_081(w_450_081, w_122_270);
  nand2 I450_115(w_450_117, w_373_024, w_450_116);
  nand2 I450_116(w_450_118, w_450_117, w_389_092);
  not1 I450_117(w_450_119, w_450_118);
  not1 I450_118(w_450_120, w_450_119);
  or2  I450_119(w_450_121, w_183_110, w_450_120);
  nand2 I450_120(w_450_122, w_246_274, w_450_121);
  nand2 I450_121(w_450_123, w_450_122, w_369_081);
  nand2 I450_122(w_450_116, w_450_123, w_158_546);
  or2  I451_379(w_451_379, w_445_017, w_401_785);
  not1 I452_044(w_452_044, w_021_340);
  or2  I452_487(w_452_487, w_102_721, w_017_009);
  and2 I453_179(w_453_179, w_412_147, w_358_438);
  or2  I454_165(w_454_165, w_318_024, w_176_361);
  nand2 I454_685(w_454_685, w_372_442, w_107_206);
  nand2 I455_040(w_455_040, w_184_049, w_009_007);
  or2  I455_105(w_455_105, w_412_746, w_137_165);
  and2 I455_112(w_455_112, w_104_176, w_241_344);
  not1 I457_023(w_457_023, w_032_180);
  and2 I457_071(w_457_071, w_090_244, w_242_223);
  nand2 I457_092(w_457_092, w_413_446, w_020_063);
  nand2 I459_131(w_459_131, w_093_484, w_044_012);
  nand2 I460_255(w_460_255, w_231_036, w_140_219);
  nand2 I460_536(w_460_536, w_163_002, w_128_146);
  and2 I461_112(w_461_112, w_040_126, w_334_002);
  not1 I461_186(w_461_186, w_431_019);
  or2  I462_369(w_462_369, w_123_062, w_113_041);
  and2 I464_156(w_464_156, w_141_088, w_070_388);
  not1 I465_326(w_465_326, w_026_239);
  or2  I465_523(w_465_523, w_120_102, w_350_011);
  not1 I466_177(w_466_177, w_447_349);
  nand2 I466_287(w_466_287, w_048_320, w_042_055);
  not1 I467_016(w_467_016, w_239_648);
  and2 I467_042(w_467_042, w_232_008, w_275_002);
  and2 I468_004(w_468_004, w_264_782, w_300_854);
  and2 I468_052(w_468_052, w_271_039, w_068_024);
  or2  I468_080(w_468_080, w_113_239, w_227_408);
  or2  I469_058(w_469_058, w_046_422, w_388_098);
  nand2 I469_209(w_469_209, w_110_123, w_130_213);
  not1 I469_565(w_469_565, w_046_733);
  or2  I470_021(w_470_021, w_284_229, w_222_045);
  and2 I471_332(w_471_332, w_253_005, w_257_512);
  and2 I471_893(w_471_893, w_306_091, w_327_007);
  or2  I474_405(w_474_405, w_030_462, w_382_610);
  and2 I474_429(w_474_431, w_474_449, w_474_430);
  nand2 I474_430(w_474_432, w_474_431, w_283_373);
  nand2 I474_431(w_474_433, w_474_432, w_344_000);
  nand2 I474_432(w_474_434, w_325_265, w_474_433);
  or2  I474_433(w_474_430, w_133_416, w_474_434);
  not1 I474_434(w_474_439, w_474_438);
  or2  I474_435(w_474_440, w_106_622, w_474_439);
  and2 I474_436(w_474_441, w_123_011, w_474_440);
  or2  I474_437(w_474_442, w_474_441, w_372_378);
  or2  I474_438(w_474_443, w_194_077, w_474_442);
  nand2 I474_439(w_474_444, w_445_024, w_474_443);
  nand2 I474_440(w_474_445, w_164_042, w_474_444);
  and2 I474_441(w_474_446, w_461_186, w_474_445);
  and2 I474_442(w_474_447, w_474_446, w_127_141);
  not1 I474_443(w_474_438, w_474_431);
  and2 I474_444(w_474_449, w_301_478, w_474_447);
  or2  I476_110(w_476_110, w_080_102, w_324_589);
  nand2 I476_174(w_476_174, w_356_701, w_132_529);
  nand2 I476_782(w_476_782, w_343_076, w_421_003);
  or2  I477_060(w_477_060, w_131_120, w_291_035);
  and2 I477_460(w_477_460, w_333_540, w_351_004);
  and2 I477_648(w_477_648, w_273_061, w_119_046);
  and2 I477_713(w_477_713, w_400_203, w_013_485);
  nand2 I478_050(w_478_050, w_260_578, w_228_329);
  not1 I479_086(w_479_086, w_229_076);
  not1 I479_183(w_479_183, w_125_007);
  and2 I479_188(w_479_188, w_011_193, w_219_069);
  or2  I480_046(w_480_046, w_477_713, w_058_015);
  nand2 I480_285(w_480_285, w_397_194, w_039_413);
  nand2 I482_031(w_482_031, w_281_115, w_109_283);
  nand2 I483_180(w_483_180, w_452_487, w_361_029);
  or2  I483_215(w_483_217, w_034_113, w_483_216);
  or2  I483_216(w_483_218, w_483_217, w_260_812);
  and2 I483_217(w_483_219, w_483_218, w_146_106);
  and2 I483_218(w_483_220, w_053_404, w_483_219);
  or2  I483_219(w_483_221, w_442_003, w_483_220);
  and2 I483_220(w_483_222, w_223_023, w_483_221);
  and2 I483_221(w_483_223, w_483_222, w_293_625);
  and2 I483_222(w_483_224, w_269_031, w_483_223);
  or2  I483_223(w_483_225, w_483_224, w_137_579);
  and2 I483_224(w_483_226, w_483_225, w_270_103);
  and2 I483_225(w_483_227, w_483_226, w_444_007);
  nand2 I483_226(w_483_216, w_019_353, w_483_227);
  or2  I484_159(w_484_159, w_423_235, w_183_053);
  nand2 I484_422(w_484_422, w_377_168, w_088_618);
  and2 I484_522(w_484_522, w_476_782, w_135_083);
  and2 I484_601(w_484_601, w_353_088, w_096_218);
  not1 I486_233(w_486_233, w_207_353);
  and2 I487_023(w_487_023, w_467_016, w_076_175);
  nand2 I487_195(w_487_195, w_470_021, w_440_458);
  or2  I487_231(w_487_231, w_325_027, w_300_631);
  not1 I488_004(w_488_004, w_442_089);
  not1 I488_061(w_488_061, w_239_183);
  or2  I488_066(w_488_066, w_407_066, w_422_041);
  nand2 I488_117(w_488_117, w_134_267, w_415_059);
  not1 I489_029(w_489_029, w_406_263);
  or2  I490_392(w_490_392, w_102_779, w_344_000);
  or2  I491_184(w_491_184, w_182_091, w_440_157);
  nand2 I491_222(w_491_222, w_454_165, w_104_024);
  not1 I491_453(w_491_453, w_295_009);
  nand2 I493_023(w_493_023, w_081_026, w_382_232);
  not1 I494_418(w_494_418, w_265_059);
  or2  I494_428(w_494_428, w_214_070, w_341_025);
  nand2 I495_061(w_495_061, w_142_130, w_068_329);
  not1 I497_072(w_497_072, w_327_728);
  nand2 I497_367(w_497_367, w_428_557, w_075_180);
  not1 I498_003(w_498_003, w_152_278);
  or2  I498_527(w_498_527, w_027_659, w_102_754);
  not1 I499_113(w_499_113, w_017_003);
  and2 I499_268(w_499_268, w_254_184, w_016_313);
  or2  I499_278(w_499_278, w_172_030, w_078_044);
  not1 I500_173(w_500_173, w_149_315);
  or2  I501_029(w_501_029, w_236_300, w_147_047);
  nand2 I501_049(w_501_049, w_053_289, w_389_335);
  and2 I502_002(w_502_002, w_175_551, w_262_110);
  nand2 I502_014(w_502_014, w_235_058, w_288_353);
  and2 I503_031(w_503_031, w_241_027, w_008_147);
  and2 I503_729(w_503_731, w_503_730, w_257_044);
  not1 I503_730(w_503_732, w_503_731);
  not1 I503_731(w_503_733, w_503_732);
  or2  I503_732(w_503_734, w_410_093, w_503_733);
  or2  I503_733(w_503_735, w_097_329, w_503_734);
  or2  I503_734(w_503_736, w_133_177, w_503_735);
  or2  I503_735(w_503_737, w_503_736, w_025_146);
  and2 I503_736(w_503_738, w_503_737, w_497_072);
  or2  I503_737(w_503_739, w_503_754, w_503_738);
  nand2 I503_738(w_503_730, w_406_437, w_503_739);
  nand2 I503_739(w_503_744, w_503_743, w_059_272);
  and2 I503_740(w_503_745, w_107_072, w_503_744);
  not1 I503_741(w_503_746, w_503_745);
  nand2 I503_742(w_503_747, w_381_632, w_503_746);
  and2 I503_743(w_503_748, w_099_070, w_503_747);
  and2 I503_744(w_503_749, w_493_023, w_503_748);
  nand2 I503_745(w_503_750, w_503_749, w_394_118);
  not1 I503_746(w_503_751, w_503_750);
  not1 I503_747(w_503_752, w_503_751);
  not1 I503_748(w_503_743, w_503_739);
  and2 I503_749(w_503_754, w_488_004, w_503_752);
  and2 I504_203(w_504_203, w_323_902, w_365_145);
  and2 I505_085(w_505_085, w_251_026, w_309_164);
  and2 I505_686(w_505_686, w_316_731, w_306_072);
  not1 I508_000(w_508_000, w_368_006);
  nand2 I509_022(w_509_022, w_105_346, w_216_102);
  and2 I509_040(w_509_040, w_094_884, w_126_118);
  not1 I510_377(w_510_377, w_442_020);
  nand2 I510_748(w_510_748, w_027_014, w_111_206);
  not1 I511_108(w_511_108, w_232_029);
  nand2 I511_753(w_511_753, w_257_146, w_269_017);
  nand2 I512_001(w_512_001, w_075_144, w_207_147);
  or2  I512_120(w_512_120, w_279_344, w_262_146);
  or2  I512_345(w_512_345, w_160_072, w_287_110);
  or2  I513_218(w_513_218, w_391_028, w_243_147);
  or2  I514_204(w_514_204, w_209_180, w_263_077);
  not1 I515_129(w_515_129, w_330_072);
  and2 I515_169(w_515_169, w_498_003, w_486_233);
  nand2 I515_535(w_515_535, w_122_208, w_380_107);
  or2  I517_397(w_517_397, w_199_419, w_383_095);
  and2 I518_369(w_518_369, w_196_728, w_439_237);
  not1 I518_760(w_518_760, w_511_753);
  not1 I519_060(w_519_060, w_422_026);
  nand2 I519_098(w_519_098, w_514_204, w_165_098);
  not1 I520_251(w_520_251, w_109_145);
  nand2 I520_860(w_520_860, w_078_053, w_159_149);
  not1 I521_000(w_521_000, w_283_079);
  not1 I524_068(w_524_068, w_309_193);
  or2  I524_639(w_524_639, w_171_280, w_494_428);
  nand2 I525_019(w_525_019, w_115_073, w_290_260);
  nand2 I525_027(w_525_027, w_211_150, w_421_159);
  not1 I526_150(w_526_150, w_435_087);
  not1 I527_041(w_527_041, w_362_083);
  and2 I527_056(w_527_056, w_166_531, w_151_034);
  not1 I527_095(w_527_095, w_452_044);
  nand2 I527_113(w_527_113, w_335_094, w_385_375);
  and2 I528_000(w_528_000, w_129_006, w_341_046);
  or2  I528_087(w_528_087, w_509_022, w_488_066);
  or2  I529_240(w_529_240, w_515_129, w_197_541);
  nand2 I529_542(w_529_542, w_089_107, w_484_422);
  not1 I529_947(w_529_947, w_313_027);
  and2 I530_171(w_530_171, w_274_000, w_469_565);
  nand2 I530_524(w_530_524, w_292_109, w_397_322);
  nand2 I531_104(w_531_104, w_453_179, w_407_039);
  not1 I531_273(w_531_273, w_140_333);
  and2 I531_352(w_531_352, w_355_160, w_477_460);
  not1 I534_277(w_534_277, w_247_611);
  not1 I536_295(w_536_295, w_340_315);
  nand2 I537_074(w_537_074, w_101_047, w_358_421);
  and2 I538_778(w_538_778, w_095_165, w_350_226);
  nand2 I539_036(w_539_036, w_109_083, w_388_100);
  not1 I539_064(w_539_064, w_015_322);
  nand2 I541_008(w_541_008, w_197_140, w_133_057);
  and2 I541_013(w_541_013, w_041_048, w_170_045);
  not1 I541_068(w_541_068, w_113_220);
  or2  I543_064(w_543_064, w_438_352, w_057_092);
  and2 I545_264(w_545_264, w_455_105, w_057_039);
  and2 I545_270(w_545_270, w_414_008, w_190_261);
  and2 I546_205(w_546_205, w_217_209, w_143_253);
  not1 I547_131(w_547_131, w_331_007);
  not1 I547_377(w_547_377, w_417_156);
  or2  I547_427(w_547_427, w_222_477, w_405_146);
  not1 I550_001(w_550_001, w_209_203);
  or2  I550_051(w_550_051, w_488_061, w_192_000);
  and2 I551_922(w_551_922, w_112_049, w_204_218);
  not1 I552_506(w_552_506, w_098_025);
  not1 I552_556(w_552_556, w_503_031);
  or2  I553_655(w_553_655, w_423_027, w_398_362);
  and2 I555_112(w_555_112, w_203_258, w_534_277);
  and2 I556_244(w_556_244, w_251_262, w_055_233);
  and2 I558_351(w_558_351, w_212_102, w_023_181);
  or2  I559_126(w_559_126, w_302_029, w_397_197);
  not1 I559_352(w_559_352, w_105_017);
  nand2 I560_550(w_560_550, w_050_370, w_539_064);
  not1 I560_731(w_560_731, w_107_025);
  and2 I561_112(w_561_112, w_154_113, w_026_056);
  and2 I562_064(w_562_064, w_460_536, w_521_000);
  not1 I563_002(w_563_002, w_016_424);
  or2  I563_007(w_563_007, w_436_111, w_154_297);
  and2 I563_029(w_563_029, w_025_022, w_394_103);
  or2  I564_518(w_564_518, w_089_088, w_318_051);
  not1 I564_612(w_564_612, w_203_156);
  not1 I565_169(w_565_169, w_477_648);
  or2  I565_447(w_565_447, w_491_453, w_465_523);
  and2 I565_579(w_565_579, w_344_001, w_060_229);
  not1 I565_627(w_565_627, w_228_288);
  nand2 I565_653(w_565_653, w_283_250, w_372_455);
  or2  I566_252(w_566_252, w_177_549, w_200_262);
  nand2 I566_464(w_566_464, w_313_170, w_172_299);
  nand2 I567_204(w_567_204, w_063_110, w_288_135);
  not1 I567_775(w_567_775, w_251_259);
  nand2 I568_144(w_568_144, w_388_244, w_193_290);
  not1 I569_371(w_569_371, w_462_369);
  not1 I570_277(w_570_277, w_146_296);
  nand2 I571_125(w_571_125, w_041_119, w_405_393);
  not1 I572_339(w_572_339, w_343_160);
  and2 I572_469(w_572_469, w_565_447, w_029_050);
  nand2 I573_015(w_573_015, w_215_092, w_238_312);
  not1 I576_060(w_576_060, w_360_035);
  nand2 I576_076(w_576_076, w_465_326, w_395_161);
  not1 I577_770(w_577_770, w_191_083);
  not1 I578_013(w_578_013, w_367_053);
  nand2 I578_116(w_578_116, w_088_189, w_280_002);
  or2  I578_266(w_578_266, w_167_416, w_314_765);
  and2 I580_001(w_580_001, w_165_187, w_331_087);
  nand2 I580_034(w_580_034, w_565_169, w_565_579);
  and2 I581_048(w_581_048, w_033_397, w_411_948);
  and2 I581_068(w_581_068, w_115_075, w_468_080);
  nand2 I581_206(w_581_206, w_027_041, w_515_169);
  or2  I582_163(w_582_163, w_099_077, w_071_436);
  nand2 I584_143(w_584_143, w_265_065, w_581_206);
  and2 I584_242(w_584_242, w_095_153, w_550_051);
  or2  I585_305(w_585_305, w_191_316, w_510_748);
  or2  I586_005(w_586_005, w_346_022, w_240_178);
  nand2 I588_655(w_588_655, w_546_205, w_351_041);
  nand2 I588_660(w_588_660, w_194_699, w_484_601);
  and2 I588_885(w_588_885, w_031_409, w_254_306);
  not1 I589_435(w_589_435, w_027_459);
  nand2 I589_696(w_589_696, w_071_286, w_051_002);
  nand2 I590_483(w_590_483, w_075_043, w_589_696);
  or2  I592_237(w_592_237, w_447_499, w_568_144);
  not1 I593_338(w_593_338, w_519_060);
  and2 I593_555(w_593_555, w_112_048, w_140_101);
  nand2 I594_047(w_594_047, w_446_650, w_301_070);
  not1 I594_071(w_594_071, w_099_082);
  not1 I594_088(w_594_088, w_412_106);
  and2 I595_052(w_595_052, w_505_085, w_578_013);
  not1 I595_289(w_595_289, w_436_087);
  and2 I597_010(w_597_010, w_256_047, w_491_184);
  and2 I597_154(w_597_154, w_402_217, w_382_405);
  not1 I597_305(w_597_305, w_519_098);
  or2  I597_328(w_597_330, w_597_329, w_597_351);
  and2 I597_329(w_597_331, w_597_330, w_362_019);
  not1 I597_330(w_597_332, w_597_331);
  nand2 I597_331(w_597_333, w_435_090, w_597_332);
  or2  I597_332(w_597_334, w_597_333, w_468_004);
  not1 I597_333(w_597_335, w_597_334);
  or2  I597_334(w_597_336, w_227_199, w_597_335);
  or2  I597_335(w_597_337, w_003_003, w_597_336);
  and2 I597_336(w_597_329, w_597_337, w_543_064);
  or2  I597_337(w_597_342, w_597_341, w_166_020);
  nand2 I597_338(w_597_343, w_558_351, w_597_342);
  nand2 I597_339(w_597_344, w_597_343, w_561_112);
  not1 I597_340(w_597_345, w_597_344);
  nand2 I597_341(w_597_346, w_530_524, w_597_345);
  and2 I597_342(w_597_347, w_167_069, w_597_346);
  and2 I597_343(w_597_348, w_597_347, w_405_439);
  not1 I597_344(w_597_349, w_597_348);
  not1 I597_345(w_597_341, w_597_330);
  and2 I597_346(w_597_351, w_277_106, w_597_349);
  nand2 I600_055(w_600_055, w_079_015, w_157_528);
  and2 I601_099(w_601_099, w_588_885, w_334_000);
  not1 I604_292(w_604_292, w_094_506);
  not1 I604_585(w_604_585, w_067_077);
  and2 I604_740(w_604_740, w_515_535, w_361_032);
  or2  I606_125(w_606_125, w_403_140, w_424_509);
  nand2 I606_297(w_606_297, w_527_113, w_108_000);
  and2 I606_398(w_606_398, w_317_533, w_447_349);
  or2  I610_161(w_610_161, w_502_002, w_527_095);
  nand2 I610_178(w_610_178, w_085_024, w_478_050);
  nand2 I611_013(w_611_013, w_188_073, w_104_042);
  and2 I612_023(w_612_023, w_604_292, w_198_322);
  and2 I613_169(w_613_169, w_173_069, w_314_086);
  or2  I613_372(w_613_372, w_093_130, w_094_124);
  not1 I614_603(w_614_603, w_499_268);
  or2  I615_006(w_615_006, w_263_199, w_025_071);
  nand2 I617_055(w_617_055, w_071_011, w_512_345);
  nand2 I618_328(w_618_328, w_219_064, w_406_047);
  nand2 I619_158(w_619_158, w_178_014, w_499_278);
  and2 I620_386(w_620_386, w_445_010, w_294_279);
  or2  I620_448(w_620_448, w_092_034, w_527_056);
  not1 I622_073(w_622_073, w_457_092);
  not1 I623_290(w_623_290, w_131_181);
  and2 I624_007(w_624_007, w_494_418, w_222_259);
  not1 I624_026(w_624_026, w_318_026);
  nand2 I625_023(w_625_023, w_624_007, w_038_388);
  or2  I626_001(w_626_001, w_342_140, w_336_047);
  or2  I628_163(w_628_163, w_185_149, w_116_011);
  not1 I630_006(w_630_006, w_620_386);
  and2 I630_101(w_630_101, w_461_112, w_296_017);
  not1 I633_074(w_633_074, w_404_049);
  nand2 I633_156(w_633_156, w_308_061, w_157_038);
  nand2 I635_153(w_635_153, w_320_101, w_501_029);
  or2  I637_226(w_637_226, w_186_618, w_162_326);
  not1 I637_537(w_637_537, w_369_005);
  nand2 I638_381(w_638_381, w_547_377, w_595_052);
  and2 I639_173(w_639_173, w_313_166, w_000_188);
  nand2 I643_784(w_643_784, w_095_163, w_614_603);
  not1 I643_889(w_643_889, w_606_297);
  and2 I644_029(w_644_029, w_630_101, w_488_117);
  and2 I644_288(w_644_288, w_163_237, w_367_243);
  and2 I644_363(w_644_363, w_210_523, w_094_415);
  and2 I644_394(w_644_394, w_356_756, w_034_792);
  and2 I646_006(w_646_006, w_521_000, w_536_295);
  not1 I646_027(w_646_027, w_388_023);
  or2  I651_087(w_651_087, w_318_038, w_646_006);
  nand2 I652_169(w_652_169, w_223_379, w_281_344);
  not1 I652_187(w_652_187, w_306_137);
  or2  I654_033(w_654_033, w_144_299, w_132_338);
  or2  I656_184(w_656_184, w_501_049, w_101_148);
  and2 I657_576(w_657_576, w_626_001, w_437_050);
  not1 I658_148(w_658_148, w_221_396);
  and2 I665_155(w_665_155, w_242_106, w_196_274);
  or2  I667_474(w_667_474, w_244_160, w_188_087);
  and2 I671_004(w_671_004, w_075_052, w_401_636);
  nand2 I671_349(w_671_349, w_566_464, w_258_236);
  nand2 I673_893(w_673_893, w_592_237, w_665_155);
  and2 I675_073(w_675_073, w_131_578, w_415_370);
  not1 I677_133(w_677_133, w_563_029);
  and2 I679_446(w_679_446, w_332_075, w_017_027);
  or2  I681_125(w_681_125, w_220_604, w_235_140);
  or2  I684_004(w_684_004, w_100_201, w_370_154);
  and2 I684_012(w_684_012, w_170_275, w_202_019);
  and2 I684_680(w_684_680, w_279_088, w_204_363);
  not1 I685_052(w_685_052, w_416_301);
  not1 I685_145(w_685_145, w_447_210);
  not1 I686_000(w_686_000, w_191_135);
  not1 I686_047(w_686_047, w_667_474);
  not1 I687_067(w_687_067, w_401_729);
  not1 I687_271(w_687_271, w_433_391);
  or2  I689_222(w_689_222, w_406_013, w_035_335);
  not1 I689_272(w_689_272, w_361_059);
  or2  I689_291(w_689_291, w_466_177, w_159_192);
  and2 I690_226(w_690_226, w_592_237, w_606_398);
  not1 I690_459(w_690_459, w_531_352);
  and2 I691_066(w_691_066, w_142_011, w_302_020);
  or2  I692_415(w_692_415, w_444_000, w_180_269);
  and2 I693_100(w_693_100, w_459_131, w_581_048);
  and2 I694_016(w_694_016, w_187_175, w_168_412);
  nand2 I698_419(w_698_419, w_037_115, w_633_074);
  not1 I700_169(w_700_169, w_162_181);
  not1 I701_285(w_701_285, w_353_057);
  and2 I701_509(w_701_509, w_637_537, w_214_092);
  not1 I702_177(w_702_177, w_180_210);
  not1 I703_212(w_703_212, w_061_070);
  and2 I703_394(w_703_396, w_703_395, w_518_369);
  and2 I703_395(w_703_397, w_703_396, w_480_285);
  or2  I703_396(w_703_398, w_703_397, w_611_013);
  nand2 I703_397(w_703_399, w_500_173, w_703_398);
  nand2 I703_398(w_703_400, w_169_034, w_703_399);
  not1 I703_399(w_703_401, w_703_400);
  nand2 I703_400(w_703_402, w_703_401, w_686_000);
  not1 I703_401(w_703_403, w_703_402);
  not1 I703_402(w_703_404, w_703_403);
  nand2 I703_403(w_703_405, w_091_002, w_703_404);
  and2 I703_404(w_703_406, w_058_128, w_703_405);
  and2 I703_405(w_703_395, w_703_406, w_428_765);
  or2  I705_598(w_705_598, w_570_277, w_004_016);
  or2  I706_150(w_706_150, w_440_495, w_098_465);
  and2 I706_155(w_706_155, w_237_423, w_034_260);
  nand2 I707_071(w_707_071, w_681_125, w_346_038);
  not1 I707_146(w_707_146, w_541_013);
  nand2 I713_009(w_713_009, w_225_026, w_241_065);
  and2 I713_132(w_713_134, w_713_151, w_713_133);
  not1 I713_133(w_713_135, w_713_134);
  or2  I713_134(w_713_133, w_713_135, w_578_266);
  nand2 I713_135(w_713_140, w_713_139, w_076_044);
  not1 I713_136(w_713_141, w_713_140);
  not1 I713_137(w_713_142, w_713_141);
  or2  I713_138(w_713_143, w_713_142, w_580_001);
  nand2 I713_139(w_713_144, w_208_026, w_713_143);
  nand2 I713_140(w_713_145, w_073_413, w_713_144);
  or2  I713_141(w_713_146, w_713_145, w_343_172);
  or2  I713_142(w_713_147, w_009_048, w_713_146);
  and2 I713_143(w_713_148, w_713_147, w_639_173);
  and2 I713_144(w_713_149, w_013_067, w_713_148);
  not1 I713_145(w_713_139, w_713_134);
  and2 I713_146(w_713_151, w_686_047, w_713_149);
  not1 I716_133(w_716_133, w_375_045);
  and2 I718_257(w_718_257, w_197_189, w_026_068);
  and2 I719_614(w_719_616, w_203_512, w_719_615);
  and2 I719_615(w_719_617, w_719_616, w_392_000);
  not1 I719_616(w_719_618, w_719_617);
  or2  I719_617(w_719_619, w_719_618, w_258_754);
  not1 I719_618(w_719_620, w_719_619);
  or2  I719_619(w_719_621, w_283_283, w_719_620);
  nand2 I719_620(w_719_622, w_300_208, w_719_621);
  nand2 I719_621(w_719_623, w_719_622, w_520_860);
  and2 I719_622(w_719_615, w_259_461, w_719_623);
  nand2 I720_811(w_720_812, w_720_811, w_365_069);
  not1 I720_812(w_720_813, w_720_812);
  not1 I720_813(w_720_814, w_720_813);
  and2 I720_814(w_720_815, w_720_814, w_179_713);
  and2 I720_815(w_720_816, w_267_225, w_720_815);
  not1 I720_816(w_720_811, w_720_816);
  not1 I721_179(w_721_179, w_654_033);
  not1 I721_271(w_721_271, w_128_094);
  not1 I722_521(w_722_521, w_593_555);
  not1 I723_185(w_723_185, w_116_032);
  or2  I729_129(w_729_129, w_637_226, w_265_068);
  not1 I730_090(w_730_090, w_283_498);
  or2  I731_104(w_731_104, w_440_479, w_716_133);
  nand2 I732_078(w_732_078, w_646_027, w_508_000);
  nand2 I737_368(w_737_368, w_525_019, w_652_169);
  not1 I737_554(w_737_556, w_737_555);
  or2  I737_555(w_737_557, w_059_214, w_737_556);
  not1 I737_556(w_737_558, w_737_557);
  or2  I737_557(w_737_559, w_223_141, w_737_558);
  or2  I737_558(w_737_560, w_096_475, w_737_559);
  nand2 I737_559(w_737_561, w_737_560, w_157_180);
  not1 I737_560(w_737_555, w_737_561);
  and2 I739_365(w_739_365, w_442_014, w_594_088);
  or2  I740_340(w_740_340, w_673_893, w_487_231);
  or2  I742_037(w_742_037, w_528_087, w_513_218);
  not1 I742_744(w_742_744, w_220_608);
  not1 I743_141(w_743_143, w_743_142);
  or2  I743_142(w_743_144, w_743_143, w_510_377);
  and2 I743_143(w_743_145, w_143_279, w_743_144);
  or2  I743_144(w_743_146, w_743_145, w_430_279);
  or2  I743_145(w_743_142, w_138_690, w_743_146);
  and2 I745_143(w_745_143, w_361_000, w_079_199);
  or2  I746_004(w_746_004, w_292_160, w_138_084);
  or2  I749_165(w_749_165, w_238_231, w_317_059);
  or2  I751_361(w_751_361, w_604_585, w_429_111);
  nand2 I753_047(w_753_047, w_495_061, w_399_050);
  nand2 I754_035(w_754_035, w_159_285, w_225_002);
  and2 I754_554(w_754_554, w_198_220, w_497_367);
  not1 I755_022(w_755_022, w_030_019);
  or2  I756_019(w_756_019, w_656_184, w_537_074);
  nand2 I757_254(w_757_254, w_189_071, w_065_855);
  nand2 I759_380(w_759_380, w_441_013, w_193_197);
  not1 I761_008(w_761_008, w_029_134);
  or2  I762_761(w_762_761, w_754_554, w_131_081);
  or2  I764_052(w_764_052, w_613_372, w_309_151);
  not1 I764_518(w_764_518, w_403_277);
  and2 I768_177(w_768_177, w_454_685, w_432_026);
  nand2 I771_065(w_771_065, w_581_068, w_072_021);
  not1 I775_531(w_775_531, w_445_037);
  nand2 I775_618(w_775_618, w_644_288, w_196_306);
  nand2 I777_041(w_777_041, w_466_287, w_433_066);
  and2 I778_142(w_778_142, w_111_162, w_143_002);
  or2  I778_263(w_778_263, w_685_052, w_413_287);
  nand2 I780_073(w_780_073, w_559_126, w_685_145);
  nand2 I783_313(w_783_313, w_414_153, w_778_142);
  or2  I784_017(w_784_017, w_524_068, w_266_451);
  nand2 I787_430(w_787_430, w_287_695, w_315_491);
  or2  I788_200(w_788_202, w_788_201, w_751_361);
  or2  I788_201(w_788_203, w_357_147, w_788_202);
  or2  I788_202(w_788_204, w_788_203, w_788_219);
  nand2 I788_203(w_788_205, w_705_598, w_788_204);
  and2 I788_204(w_788_201, w_706_150, w_788_205);
  nand2 I788_205(w_788_210, w_194_453, w_788_209);
  nand2 I788_206(w_788_211, w_788_210, w_125_190);
  nand2 I788_207(w_788_212, w_730_090, w_788_211);
  nand2 I788_208(w_788_213, w_788_212, w_764_052);
  and2 I788_209(w_788_214, w_066_210, w_788_213);
  or2  I788_210(w_788_215, w_209_171, w_788_214);
  and2 I788_211(w_788_216, w_788_215, w_138_191);
  or2  I788_212(w_788_217, w_788_216, w_759_380);
  not1 I788_213(w_788_209, w_788_204);
  and2 I788_214(w_788_219, w_045_149, w_788_217);
  or2  I789_570(w_789_570, w_143_241, w_633_156);
  nand2 I790_729(w_790_729, w_529_947, w_577_770);
  and2 I791_166(w_791_166, w_188_123, w_207_104);
  or2  I795_038(w_795_038, w_547_131, w_003_018);
  not1 I795_155(w_795_155, w_399_091);
  and2 I796_256(w_796_256, w_565_653, w_597_154);
  or2  I797_385(w_797_385, w_141_706, w_707_071);
  not1 I802_627(w_802_629, w_802_628);
  nand2 I802_628(w_802_630, w_802_629, w_344_001);
  nand2 I802_629(w_802_631, w_802_630, w_256_124);
  and2 I802_630(w_802_632, w_042_065, w_802_631);
  nand2 I802_631(w_802_633, w_423_151, w_802_632);
  and2 I802_632(w_802_634, w_802_633, w_402_188);
  nand2 I802_633(w_802_628, w_564_518, w_802_634);
  or2  I804_005(w_804_005, w_295_080, w_405_808);
  not1 I805_240(w_805_240, w_756_019);
  not1 I807_002(w_807_002, w_721_179);
  nand2 I809_082(w_809_082, w_403_276, w_315_129);
  not1 I813_317(w_813_317, w_403_085);
  and2 I820_016(w_820_016, w_199_056, w_135_123);
  or2  I821_033(w_821_033, w_584_143, w_199_131);
  not1 I822_987(w_822_989, w_822_988);
  nand2 I822_988(w_822_990, w_239_728, w_822_989);
  or2  I822_989(w_822_988, w_822_990, w_623_290);
  nand2 I826_020(w_826_020, w_253_000, w_479_086);
  or2  I826_130(w_826_130, w_749_165, w_718_257);
  and2 I828_076(w_828_076, w_499_113, w_643_784);
  not1 I828_088(w_828_088, w_286_249);
  or2  I829_086(w_829_086, w_046_546, w_186_609);
  or2  I829_467(w_829_467, w_441_004, w_504_203);
  or2  I832_482(w_832_482, w_477_060, w_630_006);
  or2  I838_328(w_838_328, w_677_133, w_215_422);
  nand2 I842_229(w_842_229, w_373_069, w_740_340);
  nand2 I843_544(w_843_544, w_092_122, w_165_120);
  or2  I844_288(w_844_288, w_761_008, w_502_014);
  nand2 I845_074(w_845_074, w_469_058, w_075_111);
  not1 I846_004(w_846_004, w_805_240);
  nand2 I847_001(w_847_003, w_197_778, w_847_002);
  nand2 I847_002(w_847_004, w_826_130, w_847_003);
  nand2 I847_003(w_847_005, w_847_004, w_004_033);
  and2 I847_004(w_847_006, w_076_422, w_847_005);
  and2 I847_005(w_847_002, w_847_006, w_202_012);
  not1 I848_326(w_848_326, w_689_222);
  and2 I848_335(w_848_335, w_778_263, w_096_160);
  nand2 I850_023(w_850_023, w_104_250, w_232_235);
  nand2 I853_747(w_853_747, w_796_256, w_687_271);
  or2  I856_011(w_856_011, w_564_612, w_418_034);
  nand2 I860_088(w_860_088, w_594_071, w_742_037);
  and2 I860_491(w_860_491, w_566_252, w_559_352);
  not1 I863_324(w_863_324, w_706_155);
  and2 I866_111(w_866_111, w_790_729, w_264_796);
  and2 I869_114(w_869_114, w_415_247, w_077_219);
  or2  I871_145(w_871_145, w_313_446, w_120_016);
  nand2 I871_351(w_871_351, w_809_082, w_324_030);
  not1 I873_255(w_873_255, w_033_630);
  nand2 I875_165(w_875_165, w_652_187, w_593_338);
  nand2 I875_251(w_875_251, w_431_024, w_383_337);
  not1 I876_001(w_876_001, w_551_922);
  not1 I878_548(w_878_548, w_043_063);
  not1 I878_681(w_878_681, w_528_000);
  not1 I878_747(w_878_749, w_878_748);
  or2  I878_748(w_878_750, w_878_749, w_635_153);
  nand2 I878_749(w_878_751, w_520_251, w_878_750);
  not1 I878_750(w_878_752, w_878_751);
  and2 I878_751(w_878_753, w_033_352, w_878_752);
  or2  I878_752(w_878_754, w_878_753, w_878_766);
  or2  I878_753(w_878_755, w_539_036, w_878_754);
  and2 I878_754(w_878_748, w_451_379, w_878_755);
  not1 I878_755(w_878_760, w_878_759);
  nand2 I878_756(w_878_761, w_878_760, w_396_533);
  nand2 I878_757(w_878_762, w_658_148, w_878_761);
  nand2 I878_758(w_878_763, w_878_762, w_527_041);
  or2  I878_759(w_878_764, w_878_763, w_155_027);
  not1 I878_760(w_878_759, w_878_754);
  and2 I878_761(w_878_766, w_529_542, w_878_764);
  not1 I881_105(w_881_105, w_550_001);
  not1 I882_423(w_882_423, w_144_234);
  nand2 I883_420(w_883_420, w_742_744, w_320_029);
  nand2 I887_066(w_887_066, w_578_116, w_222_662);
  nand2 I888_266(w_888_266, w_563_002, w_221_550);
  nand2 I889_143(w_889_143, w_856_011, w_871_145);
  and2 I889_239(w_889_239, w_393_323, w_207_023);
  and2 I889_352(w_889_352, w_484_159, w_062_252);
  and2 I891_119(w_891_119, w_245_277, w_889_352);
  nand2 I891_163(w_891_163, w_397_098, w_302_023);
  not1 I893_103(w_893_103, w_846_004);
  not1 I893_145(w_893_145, w_606_125);
  not1 I894_261(w_894_263, w_894_262);
  not1 I894_262(w_894_264, w_894_263);
  and2 I894_263(w_894_265, w_305_093, w_894_264);
  or2  I894_264(w_894_266, w_894_265, w_437_069);
  nand2 I894_265(w_894_267, w_125_022, w_894_266);
  or2  I894_266(w_894_268, w_894_267, w_206_334);
  nand2 I894_267(w_894_269, w_894_268, w_624_026);
  nand2 I894_268(w_894_270, w_894_269, w_894_287);
  or2  I894_269(w_894_271, w_894_270, w_468_052);
  and2 I894_270(w_894_272, w_894_271, w_395_103);
  and2 I894_271(w_894_273, w_130_002, w_894_272);
  nand2 I894_272(w_894_262, w_894_273, w_620_448);
  not1 I894_273(w_894_278, w_894_277);
  and2 I894_274(w_894_279, w_894_278, w_511_108);
  not1 I894_275(w_894_280, w_894_279);
  not1 I894_276(w_894_281, w_894_280);
  or2  I894_277(w_894_282, w_894_281, w_449_078);
  or2  I894_278(w_894_283, w_095_040, w_894_282);
  or2  I894_279(w_894_284, w_068_024, w_894_283);
  and2 I894_280(w_894_285, w_280_023, w_894_284);
  not1 I894_281(w_894_277, w_894_270);
  and2 I894_282(w_894_287, w_008_129, w_894_285);
  and2 I896_754(w_896_756, w_896_755, w_149_392);
  not1 I896_755(w_896_757, w_896_756);
  nand2 I896_756(w_896_758, w_896_757, w_300_036);
  nand2 I896_757(w_896_755, w_182_210, w_896_758);
  and2 I899_530(w_899_532, w_899_531, w_476_174);
  and2 I899_531(w_899_533, w_597_010, w_899_532);
  and2 I899_532(w_899_534, w_427_082, w_899_533);
  and2 I899_533(w_899_535, w_553_655, w_899_534);
  nand2 I899_534(w_899_536, w_745_143, w_899_535);
  not1 I899_535(w_899_537, w_899_536);
  or2  I899_536(w_899_538, w_266_295, w_899_537);
  and2 I899_537(w_899_539, w_899_538, w_471_893);
  or2  I899_538(w_899_540, w_129_011, w_899_539);
  and2 I899_539(w_899_531, w_899_540, w_754_035);
  not1 I901_380(w_901_380, w_529_240);
  or2  I904_126(w_904_126, w_420_527, w_152_059);
  or2  I905_809(w_905_811, w_905_810, w_320_609);
  and2 I905_810(w_905_812, w_905_823, w_905_811);
  or2  I905_811(w_905_810, w_905_812, w_580_034);
  and2 I905_812(w_905_817, w_156_622, w_905_816);
  nand2 I905_813(w_905_818, w_905_817, w_377_284);
  or2  I905_814(w_905_819, w_905_818, w_205_113);
  and2 I905_815(w_905_820, w_721_271, w_905_819);
  nand2 I905_816(w_905_821, w_842_229, w_905_820);
  not1 I905_817(w_905_816, w_905_812);
  and2 I905_818(w_905_823, w_572_339, w_905_821);
  nand2 I907_282(w_907_282, w_342_109, w_713_009);
  nand2 I908_298(w_908_298, w_134_203, w_585_305);
  nand2 I914_427(w_914_427, w_908_298, w_904_126);
  and2 I916_185(w_916_185, w_317_562, w_882_423);
  or2  I916_358(w_916_358, w_878_681, w_341_018);
  or2  I919_108(w_919_108, w_059_154, w_813_317);
  not1 I919_354(w_919_354, w_916_185);
  and2 I921_163(w_921_163, w_073_114, w_379_001);
  nand2 I924_279(w_924_279, w_121_124, w_029_082);
  nand2 I924_298(w_924_298, w_619_158, w_317_043);
  and2 I927_320(w_927_320, w_919_354, w_293_573);
  and2 I928_157(w_928_157, w_349_067, w_590_483);
  or2  I930_000(w_930_000, w_293_697, w_588_660);
  nand2 I931_517(w_931_517, w_457_071, w_111_146);
  nand2 I933_375(w_933_375, w_436_096, w_571_125);
  nand2 I935_942(w_935_942, w_694_016, w_200_166);
  nand2 I935_968(w_935_970, w_610_178, w_935_969);
  nand2 I935_969(w_935_971, w_935_970, w_498_527);
  and2 I935_970(w_935_972, w_804_005, w_935_971);
  nand2 I935_971(w_935_973, w_567_775, w_935_972);
  or2  I935_972(w_935_969, w_935_973, w_935_981);
  nand2 I935_973(w_935_978, w_927_320, w_935_977);
  and2 I935_974(w_935_979, w_538_778, w_935_978);
  not1 I935_975(w_935_977, w_935_969);
  and2 I935_976(w_935_981, w_552_506, w_935_979);
  and2 I938_341(w_938_341, w_613_169, w_891_119);
  not1 I942_549(w_942_549, w_193_042);
  or2  I943_456(w_943_456, w_058_191, w_126_112);
  or2  I945_256(w_945_256, w_930_000, w_687_067);
  or2  I949_032(w_949_032, w_893_103, w_601_099);
  or2  I952_565(w_952_565, w_247_092, w_707_146);
  or2  I952_772(w_952_772, w_178_943, w_517_397);
  nand2 I954_012(w_954_012, w_185_202, w_829_467);
  nand2 I955_092(w_955_092, w_401_500, w_238_285);
  and2 I955_347(w_955_349, w_955_348, w_287_109);
  and2 I955_348(w_955_350, w_689_291, w_955_349);
  or2  I955_349(w_955_351, w_450_081, w_955_350);
  not1 I955_350(w_955_352, w_955_351);
  and2 I955_351(w_955_353, w_289_855, w_955_352);
  and2 I955_352(w_955_354, w_628_163, w_955_353);
  not1 I955_353(w_955_355, w_955_354);
  not1 I955_354(w_955_356, w_955_355);
  and2 I955_355(w_955_357, w_132_166, w_955_356);
  or2  I955_356(w_955_348, w_509_040, w_955_357);
  or2  I966_010(w_966_010, w_086_652, w_139_001);
  nand2 I966_534(w_966_534, w_572_469, w_304_064);
  or2  I967_137(w_967_137, w_025_225, w_358_031);
  and2 I968_915(w_968_917, w_968_936, w_968_916);
  or2  I968_916(w_968_918, w_968_917, w_097_495);
  not1 I968_917(w_968_919, w_968_918);
  nand2 I968_918(w_968_920, w_968_919, w_146_314);
  or2  I968_919(w_968_921, w_691_066, w_968_920);
  nand2 I968_920(w_968_922, w_076_142, w_968_921);
  or2  I968_921(w_968_923, w_968_922, w_280_016);
  or2  I968_922(w_968_924, w_968_923, w_560_550);
  nand2 I968_923(w_968_925, w_238_080, w_968_924);
  not1 I968_924(w_968_926, w_968_925);
  not1 I968_925(w_968_927, w_968_926);
  not1 I968_926(w_968_916, w_968_927);
  and2 I968_927(w_968_932, w_556_244, w_968_931);
  and2 I968_928(w_968_933, w_292_413, w_968_932);
  and2 I968_929(w_968_934, w_644_363, w_968_933);
  not1 I968_930(w_968_931, w_968_917);
  and2 I968_931(w_968_936, w_170_407, w_968_934);
  nand2 I971_279(w_971_281, w_971_280, w_340_120);
  nand2 I971_280(w_971_282, w_210_681, w_971_281);
  not1 I971_281(w_971_283, w_971_282);
  or2  I971_282(w_971_284, w_971_283, w_367_133);
  or2  I971_283(w_971_285, w_187_161, w_971_284);
  nand2 I971_284(w_971_286, w_971_285, w_484_522);
  or2  I971_285(w_971_287, w_214_075, w_971_286);
  or2  I971_286(w_971_288, w_971_287, w_154_004);
  or2  I971_287(w_971_280, w_971_288, w_444_005);
  not1 I973_121(w_973_121, w_863_324);
  nand2 I974_075(w_974_075, w_479_183, w_198_315);
  and2 I975_059(w_975_059, w_158_356, w_380_030);
  nand2 I977_099(w_977_099, w_137_554, w_073_292);
  or2  I978_339(w_978_339, w_643_889, w_679_446);
  and2 I980_815(w_980_815, w_768_177, w_866_111);
  and2 I982_324(w_982_324, w_070_256, w_176_201);
  nand2 I986_106(w_986_106, w_780_073, w_722_521);
  nand2 I986_714(w_986_714, w_881_105, w_876_001);
  nand2 I991_282(w_991_282, w_197_237, w_427_096);
  and2 I996_052(w_996_052, w_889_143, w_417_005);
  or2  I1000_000(w_1000_000, w_545_264, w_919_108);
  or2  I1000_001(w_1000_001, w_921_163, w_060_246);
  not1 I1000_002(w_1000_002, w_512_001);
  and2 I1000_003(w_1000_003, w_192_000, w_037_067);
  and2 I1000_004(w_1000_004, w_251_208, w_239_678);
  and2 I1000_005(w_1000_005, w_431_025, w_690_226);
  and2 I1000_006(w_1000_006, w_887_066, w_845_074);
  and2 I1000_007(w_1000_007, w_764_518, w_505_686);
  not1 I1000_008(w_1000_008, w_565_627);
  or2  I1000_009(w_1000_009, w_429_135, w_109_049);
  or2  I1000_010(w_1000_010, w_146_274, w_017_022);
  or2  I1000_011(w_1000_011, w_257_428, w_198_040);
  and2 I1000_012(w_1000_012, w_888_266, w_304_079);
  not1 I1000_013(w_1000_013, w_149_559);
  not1 I1000_014(w_1000_014, w_266_429);
  nand2 I1000_015(w_1000_015, w_952_772, w_112_013);
  or2  I1000_016(w_1000_016, w_541_068, w_234_515);
  nand2 I1000_017(w_1000_017, w_732_078, w_832_482);
  not1 I1000_018(w_1000_018, w_441_011);
  and2 I1000_019(w_1000_019, w_482_031, w_693_100);
  nand2 I1000_020(w_1000_020, w_820_016, w_176_380);
  and2 I1000_021(w_1000_021, w_442_053, w_211_050);
  or2  I1000_022(w_1000_022, w_323_678, w_410_001);
  nand2 I1000_023(w_1000_023, w_996_052, w_186_042);
  or2  I1000_024(w_1000_024, w_371_053, w_479_188);
  not1 I1000_025(w_1000_025, w_284_079);
  or2  I1000_026(w_1000_026, w_977_099, w_576_076);
  or2  I1000_027(w_1000_027, w_753_047, w_386_195);
  nand2 I1000_028(w_1000_028, w_949_032, w_328_273);
  and2 I1000_029(w_1000_029, w_739_365, w_991_282);
  not1 I1000_030(w_1000_030, w_530_171);
  nand2 I1000_031(w_1000_031, w_901_380, w_278_065);
  not1 I1000_032(w_1000_032, w_562_064);
  and2 I1000_033(w_1000_033, w_891_163, w_684_004);
  and2 I1000_034(w_1000_034, w_789_570, w_974_075);
  or2  I1000_035(w_1000_035, w_924_279, w_942_549);
  nand2 I1000_036(w_1000_036, w_033_391, w_594_047);
  or2  I1000_037(w_1000_037, w_476_110, w_116_041);
  or2  I1000_038(w_1000_038, w_746_004, w_875_251);
  nand2 I1000_039(w_1000_039, w_335_105, w_374_012);
  or2  I1000_040(w_1000_040, w_610_161, w_164_131);
  not1 I1000_041(w_1000_041, w_777_041);
  or2  I1000_042(w_1000_042, w_071_058, w_380_104);
  or2  I1000_043(w_1000_043, w_327_873, w_118_190);
  not1 I1000_044(w_1000_044, w_586_005);
  nand2 I1000_045(w_1000_045, w_684_680, w_354_345);
  nand2 I1000_046(w_1000_046, w_042_018, w_265_414);
  nand2 I1000_047(w_1000_047, w_875_165, w_359_460);
  not1 I1000_048(w_1000_048, w_489_029);
  nand2 I1000_049(w_1000_049, w_560_731, w_288_665);
  and2 I1000_050(w_1000_050, w_615_006, w_002_272);
  and2 I1000_051(w_1000_051, w_588_655, w_531_273);
  nand2 I1000_052(w_1000_052, w_237_376, w_226_013);
  and2 I1000_053(w_1000_053, w_491_222, w_416_719);
  or2  I1000_054(w_1000_054, w_775_531, w_399_064);
  or2  I1000_055(w_1000_055, w_954_012, w_584_242);
  not1 I1000_056(w_1000_056, w_469_209);
  and2 I1000_057(w_1000_057, w_471_332, w_432_022);
  nand2 I1000_058(w_1000_058, w_315_105, w_675_073);
  nand2 I1000_059(w_1000_059, w_253_048, w_228_745);
  or2  I1000_060(w_1000_060, w_644_394, w_850_023);
  nand2 I1000_061(w_1000_061, w_249_036, w_552_556);
  or2  I1000_062(w_1000_062, w_137_150, w_703_212);
  and2 I1000_063(w_1000_063, w_435_077, w_044_219);
  or2  I1000_064(w_1000_064, w_383_005, w_526_150);
  not1 I1000_065(w_1000_065, w_182_038);
  not1 I1000_066(w_1000_066, w_762_761);
  and2 I1000_067(w_1000_067, w_406_577, w_702_177);
  and2 I1000_068(w_1000_068, w_952_565, w_829_086);
  not1 I1000_069(w_1000_069, w_966_010);
  or2  I1000_070(w_1000_070, w_924_298, w_268_353);
  not1 I1000_071(w_1000_071, w_487_195);
  not1 I1000_072(w_1000_072, w_021_360);
  and2 I1000_073(w_1000_073, w_460_255, w_928_157);
  or2  I1000_074(w_1000_074, w_689_272, w_775_618);
  or2  I1000_075(w_1000_075, w_305_009, w_237_276);
  and2 I1000_076(w_1000_076, w_449_110, w_690_459);
  not1 I1000_077(w_1000_077, w_966_534);
  nand2 I1000_078(w_1000_078, w_671_004, w_238_218);
  not1 I1000_079(w_1000_079, w_612_023);
  nand2 I1000_080(w_1000_080, w_072_008, w_755_022);
  or2  I1000_081(w_1000_081, w_797_385, w_692_415);
  not1 I1000_082(w_1000_082, w_349_088);
  nand2 I1000_083(w_1000_083, w_220_034, w_060_183);
  and2 I1000_084(w_1000_084, w_871_351, w_042_057);
  not1 I1000_085(w_1000_085, w_066_249);
  or2  I1000_086(w_1000_086, w_284_405, w_657_576);
  nand2 I1000_087(w_1000_087, w_729_129, w_555_112);
  or2  I1000_088(w_1000_088, w_352_100, w_437_005);
  not1 I1000_089(w_1000_089, w_787_430);
  or2  I1000_090(w_1000_090, w_007_464, w_313_228);
  or2  I1000_091(w_1000_091, w_185_061, w_935_942);
  not1 I1000_092(w_1000_092, w_001_056);
  nand2 I1000_093(w_1000_093, w_638_381, w_088_214);
  and2 I1000_094(w_1000_094, w_169_042, w_087_052);
  nand2 I1000_095(w_1000_095, w_791_166, w_873_255);
  nand2 I1000_096(w_1000_096, w_012_341, w_569_371);
  or2  I1000_097(w_1000_097, w_234_050, w_698_419);
  not1 I1000_098(w_1000_098, w_986_714);
  and2 I1000_099(w_1000_099, w_339_117, w_403_278);
  nand2 I1000_100(w_1000_100, w_843_544, w_684_012);
  not1 I1000_101(w_1000_101, w_771_065);
  not1 I1000_102(w_1000_102, w_563_007);
  nand2 I1000_103(w_1000_103, w_474_405, w_259_167);
  not1 I1000_104(w_1000_104, w_982_324);
  or2  I1000_105(w_1000_105, w_933_375, w_980_815);
  or2  I1000_106(w_1000_106, w_046_006, w_700_169);
  nand2 I1000_107(w_1000_107, w_030_176, w_035_574);
  and2 I1000_108(w_1000_108, w_399_008, w_480_046);
  not1 I1000_109(w_1000_109, w_395_026);
  or2  I1000_110(w_1000_110, w_869_114, w_040_026);
  not1 I1000_111(w_1000_111, w_022_159);
  nand2 I1000_112(w_1000_112, w_955_092, w_828_076);
  and2 I1000_113(w_1000_113, w_226_001, w_853_747);
  not1 I1000_114(w_1000_114, w_883_420);
  or2  I1000_115(w_1000_115, w_457_023, w_889_239);
  and2 I1000_116(w_1000_116, w_353_080, w_003_034);
  or2  I1000_117(w_1000_117, w_224_052, w_622_073);
  not1 I1000_118(w_1000_118, w_644_029);
  not1 I1000_119(w_1000_119, w_600_055);
  not1 I1000_120(w_1000_120, w_723_185);
  and2 I1000_121(w_1000_121, w_986_106, w_860_088);
  or2  I1000_122(w_1000_122, w_280_018, w_518_760);
  nand2 I1000_123(w_1000_123, w_487_023, w_524_639);
  and2 I1000_124(w_1000_124, w_784_017, w_301_356);
  nand2 I1000_125(w_1000_125, w_265_202, w_191_294);
  or2  I1000_126(w_1000_126, w_143_115, w_455_040);
  and2 I1000_127(w_1000_127, w_567_204, w_914_427);
  or2  I1000_128(w_1000_128, w_975_059, w_223_493);
  and2 I1000_129(w_1000_129, w_394_129, w_541_008);
  and2 I1000_130(w_1000_130, w_617_055, w_545_270);
  nand2 I1000_131(w_1000_131, w_092_033, w_626_001);
  not1 I1000_132(w_1000_132, w_547_427);
  or2  I1000_133(w_1000_133, w_002_147, w_737_368);
  not1 I1000_134(w_1000_134, w_003_023);
  nand2 I1000_135(w_1000_135, w_978_339, w_070_823);
  or2  I1000_136(w_1000_136, w_464_156, w_826_020);
  and2 I1000_137(w_1000_137, w_795_155, w_377_418);
  or2  I1000_138(w_1000_138, w_821_033, w_531_104);
  and2 I1000_139(w_1000_139, w_079_112, w_194_433);
  or2  I1000_140(w_1000_140, w_283_355, w_731_104);
  or2  I1000_141(w_1000_141, w_226_013, w_170_199);
  or2  I1000_142(w_1000_142, w_455_112, w_597_305);
  not1 I1000_143(w_1000_143, w_429_153);
  and2 I1000_144(w_1000_144, w_158_198, w_893_145);
  and2 I1000_145(w_1000_145, w_424_083, w_049_855);
  nand2 I1000_146(w_1000_146, w_595_289, w_848_326);
  and2 I1000_147(w_1000_147, w_931_517, w_701_509);
  nand2 I1000_148(w_1000_148, w_223_157, w_576_060);
  or2  I1000_149(w_1000_149, w_525_027, w_467_042);
  and2 I1000_150(w_1000_150, w_807_002, w_290_052);
  nand2 I1000_151(w_1000_151, w_147_140, w_878_548);
  and2 I1000_152(w_1000_152, w_197_143, w_973_121);
  or2  I1000_153(w_1000_153, w_618_328, w_243_109);
  or2  I1000_154(w_1000_154, w_378_247, w_346_024);
  or2  I1000_155(w_1000_155, w_967_137, w_589_435);
  or2  I1000_156(w_1000_156, w_033_594, w_249_065);
  nand2 I1000_157(w_1000_157, w_044_174, w_828_088);
  not1 I1000_158(w_1000_158, w_512_120);
  or2  I1000_159(w_1000_159, w_838_328, w_943_456);
  not1 I1000_160(w_1000_160, w_186_479);
  nand2 I1000_161(w_1000_161, w_916_358, w_086_222);
  and2 I1000_162(w_1000_162, w_053_053, w_945_256);
  not1 I1000_163(w_1000_163, w_330_151);
  nand2 I1000_164(w_1000_164, w_005_211, w_483_180);
  not1 I1000_165(w_1000_165, w_757_254);
  not1 I1000_166(w_1000_166, w_229_125);
  and2 I1000_167(w_1000_167, w_099_059, w_124_649);
  or2  I1000_168(w_1000_168, w_604_740, w_573_015);
  not1 I1000_169(w_1000_169, w_795_038);
  and2 I1000_170(w_1000_170, w_848_335, w_424_038);
  or2  I1000_171(w_1000_171, w_211_133, w_671_349);
  and2 I1000_172(w_1000_172, w_203_407, w_421_146);
  not1 I1000_173(w_1000_173, w_651_087);
  not1 I1000_174(w_1000_174, w_102_400);
  nand2 I1000_175(w_1000_175, w_103_057, w_191_325);
  not1 I1000_176(w_1000_176, w_225_022);
  or2  I1000_177(w_1000_177, w_264_606, w_625_023);
  not1 I1000_178(w_1000_178, w_015_265);
  not1 I1000_179(w_1000_179, w_844_288);
  nand2 I1000_180(w_1000_180, w_860_491, w_907_282);
  and2 I1000_181(w_1000_181, w_701_285, w_582_163);
  nand2 I1000_182(w_1000_182, w_334_002, w_490_392);
  or2  I1000_183(w_1000_183, w_333_374, w_167_042);
  and2 I1000_184(w_1000_184, w_783_313, w_129_006);
  and2 I1000_185(w_1000_185, w_145_054, w_938_341);

  initial begin
    $get_module_info();
  end
endmodule

// ****** Combined Logic Module Defination ******

// ****** TestBench Module Defination ******

/*
module tb();
  wire  w_000_000, w_000_001, w_000_002, w_000_003, w_000_004, w_000_005, w_000_006, w_000_007, w_000_008, w_000_009, w_000_010, w_000_011, w_000_012, w_000_013, w_000_014, w_000_015, w_000_016, w_000_017, w_000_018, w_000_019, w_000_020, w_000_021, w_000_022, w_000_023, w_000_024, w_000_025, w_000_026, w_000_027, w_000_028, w_000_029, w_000_030, w_000_031, w_000_032, w_000_033, w_000_034, w_000_035, w_000_036, w_000_037, w_000_038, w_000_039, w_000_040, w_000_041, w_000_042, w_000_043, w_000_044, w_000_045, w_000_046, w_000_047, w_000_048, w_000_049, w_000_050, w_000_051, w_000_052, w_000_053, w_000_054, w_000_055, w_000_056, w_000_057, w_000_058, w_000_059, w_000_060, w_000_061, w_000_062, w_000_063, w_000_064, w_000_065, w_000_066, w_000_067, w_000_068, w_000_069, w_000_070, w_000_071, w_000_072, w_000_073, w_000_074, w_000_075, w_000_076, w_000_077, w_000_078, w_000_079, w_000_080, w_000_081, w_000_082, w_000_083, w_000_084, w_000_085, w_000_086, w_000_087, w_000_088, w_000_089, w_000_090, w_000_091, w_000_092, w_000_093, w_000_094, w_000_095, w_000_096, w_000_097, w_000_098, w_000_099, w_000_100, w_000_101, w_000_102, w_000_103, w_000_104, w_000_105, w_000_106, w_000_107, w_000_108, w_000_109, w_000_110, w_000_111, w_000_112, w_000_113, w_000_114, w_000_115, w_000_116, w_000_117, w_000_118, w_000_119, w_000_120, w_000_121, w_000_122, w_000_123, w_000_124, w_000_125, w_000_126, w_000_127, w_000_128, w_000_129, w_000_130, w_000_131, w_000_132, w_000_133, w_000_134, w_000_135, w_000_136, w_000_137, w_000_138, w_000_139, w_000_140, w_000_141, w_000_142, w_000_143, w_000_144, w_000_145, w_000_146, w_000_147, w_000_148, w_000_149, w_000_150, w_000_151, w_000_152, w_000_153, w_000_154, w_000_155, w_000_156, w_000_157, w_000_158, w_000_159, w_000_160, w_000_161, w_000_162, w_000_163, w_000_164, w_000_165, w_000_166, w_000_167, w_000_168, w_000_169, w_000_170, w_000_171, w_000_172, w_000_173, w_000_174, w_000_175, w_000_176, w_000_177, w_000_178, w_000_179, w_000_180, w_000_181, w_000_182, w_000_183, w_000_184, w_000_185, w_000_186, w_000_187, w_000_188, w_000_189, w_000_190, w_000_191, w_000_192, w_000_193, w_000_194, w_000_195, w_000_196, w_000_197, w_000_198, w_000_199, w_000_200, w_000_201, w_000_202, w_000_203, w_000_204, w_000_205, w_000_206, w_000_207, w_000_208, w_000_209, w_000_210, w_000_211, w_000_212, w_000_213, w_000_214, w_000_215, w_000_216, w_000_217, w_000_218, w_000_219, w_000_220, w_000_221, w_000_222, w_000_223, w_000_224, w_000_225, w_000_226, w_000_227, w_000_228, w_000_230, w_000_231, w_000_232, w_000_233, w_000_234, w_000_235, w_000_236, w_000_237, w_000_238, w_000_239, w_000_240, w_000_241, w_000_242, w_000_243, w_000_244, w_000_245, w_000_246, w_000_247, w_000_248, w_000_249, w_000_250, w_000_251, w_000_252, w_000_253, w_000_254, w_000_255, w_000_256, w_000_257, w_000_258, w_000_259, w_000_260, w_000_262, w_000_263, w_000_264, w_000_265, w_000_266, w_000_267, w_000_268, w_000_269, w_000_270, w_000_271, w_000_272, w_000_273, w_000_274, w_000_275, w_000_276, w_000_277, w_000_278, w_000_279, w_000_280, w_000_281, w_000_282, w_000_283, w_000_284, w_000_285, w_000_286, w_000_287, w_000_288, w_000_289, w_000_290, w_000_291, w_000_292, w_000_293, w_000_294, w_000_295, w_000_296, w_000_297, w_000_298, w_000_299, w_000_300, w_000_301, w_000_302, w_000_303, w_000_304, w_000_305, w_000_306, w_000_307, w_000_308, w_000_309, w_000_310, w_000_311, w_000_312, w_000_313, w_000_314, w_000_315, w_000_316, w_000_317, w_000_318, w_000_319, w_000_320, w_000_321, w_000_322, w_000_323, w_000_324, w_000_325, w_000_326, w_000_327, w_000_328, w_000_329, w_000_330, w_000_331, w_000_332, w_000_333, w_000_334, w_000_335, w_000_336, w_000_337, w_000_338, w_000_339, w_000_340, w_000_341, w_000_342, w_000_343, w_000_344, w_000_345, w_000_346, w_000_347, w_000_348, w_000_349, w_000_350, w_000_351, w_000_352, w_000_353, w_000_354, w_000_355, w_000_356, w_000_357, w_000_358, w_000_359, w_000_360, w_000_361, w_000_362, w_000_364, w_000_365, w_000_366, w_000_367, w_000_369, w_000_370, w_000_371, w_000_372, w_000_373, w_000_374, w_000_375, w_000_376, w_000_377, w_000_378, w_000_379, w_000_380, w_000_381, w_000_382, w_000_383, w_000_384, w_000_385, w_000_386, w_000_387, w_000_388, w_000_389, w_000_390, w_000_391, w_000_392, w_000_393, w_000_394, w_000_395, w_000_396, w_000_397, w_000_398, w_000_399, w_000_400, w_000_401, w_000_402, w_000_403, w_000_404, w_000_405, w_000_406, w_000_407, w_000_408, w_000_409, w_000_410, w_000_411, w_000_412, w_000_413, w_000_414, w_000_415, w_000_416, w_000_417, w_000_418, w_000_419, w_000_420, w_000_421, w_000_422, w_000_423, w_000_424, w_000_425, w_000_426, w_000_427, w_000_428, w_000_429, w_000_430, w_000_431, w_000_432, w_000_433, w_000_434, w_000_435, w_000_436, w_000_437, w_000_438, w_000_439, w_000_440, w_000_441, w_000_442, w_000_443, w_000_444, w_000_445, w_000_446, w_000_447, w_000_448, w_000_449, w_000_450, w_000_451, w_000_452, w_000_453, w_000_454, w_000_455, w_000_456, w_000_457, w_000_458, w_000_459, w_000_460, w_000_461, w_000_462, w_000_463, w_000_464, w_000_465, w_000_466, w_000_467, w_000_468, w_000_469, w_000_470, w_000_471, w_000_472, w_000_473, w_000_474, w_000_475, w_000_476, w_000_477, w_000_478, w_000_479, w_000_480, w_000_481, w_000_482, w_000_483, w_000_484, w_000_485, w_000_486, w_000_487, w_000_488, w_000_489, w_000_490, w_000_491, w_000_492, w_000_493, w_000_494, w_000_495, w_000_496, w_000_497, w_000_498, w_000_499, w_000_500, w_000_501, w_000_502, w_000_503, w_000_504, w_000_505, w_000_506, w_000_507, w_000_508, w_000_509, w_000_510, w_000_511, w_000_512, w_000_513, w_000_514, w_000_515, w_000_516, w_000_517, w_000_518, w_000_519, w_000_520, w_000_521, w_000_522, w_000_523, w_000_524, w_000_525, w_000_526, w_000_527, w_000_528, w_000_529, w_000_530, w_000_531, w_000_532, w_000_533, w_000_534, w_000_535, w_000_536, w_000_537, w_000_538, w_000_539, w_000_540, w_000_541, w_000_542, w_000_543, w_000_544, w_000_545, w_000_546, w_000_547, w_000_548, w_000_549, w_000_550, w_000_551, w_000_552, w_000_553, w_000_554, w_000_555, w_000_556, w_000_557, w_000_558, w_000_559, w_000_560, w_000_561, w_000_562, w_000_563, w_000_564, w_000_565, w_000_566, w_000_567, w_000_568, w_000_569, w_000_570, w_000_571, w_000_572, w_000_573, w_000_574, w_000_575, w_000_576, w_000_577, w_000_578, w_000_579, w_000_580, w_000_581, w_000_582, w_000_583, w_000_584, w_000_585, w_000_586, w_000_587, w_000_588, w_000_589, w_000_590, w_000_591, w_000_592, w_000_593, w_000_594, w_000_595, w_000_596, w_000_597, w_000_598, w_000_599, w_000_600, w_000_601, w_000_602, w_000_603, w_000_604, w_000_605, w_000_606, w_000_607, w_000_608, w_000_609, w_000_610, w_000_611, w_000_612, w_000_613, w_000_614, w_000_615, w_000_616, w_000_617, w_000_618, w_000_619, w_000_620, w_000_621, w_000_622, w_000_623, w_000_624, w_000_625, w_000_626, w_000_627, w_000_628, w_000_629, w_000_630, w_000_631, w_000_632, w_000_633, w_000_634, w_000_635, w_000_636, w_000_637, w_000_638, w_000_639, w_000_640, w_000_641, w_000_642, w_000_643, w_000_644, w_000_645, w_000_646, w_000_647, w_000_648, w_000_649, w_000_650, w_000_651, w_000_652, w_000_653, w_000_654, w_000_655, w_000_656, w_000_657, w_000_658, w_000_659, w_000_660, w_000_661, w_000_662, w_000_663, w_000_664, w_000_665, w_000_666, w_000_667, w_000_669, w_000_670, w_000_671, w_000_672, w_000_673, w_000_674, w_000_675, w_000_676, w_000_677, w_000_678, w_000_679, w_000_680, w_000_681, w_000_682, w_000_683, w_000_684, w_000_685, w_000_686, w_000_687, w_000_688, w_000_689, w_000_690, w_000_691, w_000_692, w_000_693, w_000_694, w_000_695, w_000_696, w_000_697, w_000_698, w_000_699, w_000_700, w_000_701, w_000_702, w_000_703, w_000_704, w_000_705, w_000_706, w_000_707, w_000_708, w_000_709, w_000_710, w_000_711, w_000_712, w_000_713, w_000_714, w_000_715, w_000_716, w_000_717, w_000_718, w_000_719, w_000_720, w_000_721, w_000_722, w_000_723, w_000_724, w_000_725, w_000_726, w_000_727, w_000_728, w_000_729, w_000_730, w_000_731, w_000_732, w_000_733, w_000_734, w_000_735, w_000_736, w_000_737, w_000_738, w_000_739, w_000_740, w_000_741, w_000_742, w_000_743, w_000_744, w_000_745, w_000_746, w_000_747, w_000_748, w_000_749, w_000_750, w_000_751, w_000_752, w_000_753, w_000_754, w_000_755, w_000_756, w_000_757, w_000_758, w_000_759, w_000_760, w_000_761, w_000_762, w_000_763, w_000_765, w_000_766, w_000_767, w_000_769, w_000_770, w_000_772, w_000_773, w_000_774, w_000_775, w_000_776, w_000_777, w_000_779, w_000_780, w_000_781, w_000_782, w_000_783, w_000_784, w_000_785, w_000_786, w_000_787, w_000_788, w_000_789, w_000_790, w_000_791, w_000_792, w_000_793, w_000_794, w_000_795, w_000_796, w_000_797, w_000_798, w_000_799, w_000_801, w_000_802, w_000_803, w_000_804, w_000_805, w_000_806, w_000_807, w_000_808, w_000_809, w_000_810, w_000_811, w_000_812, w_000_813, w_000_814, w_000_815, w_000_816, w_000_817, w_000_818, w_000_819, w_000_820, w_000_821, w_000_822, w_000_823, w_000_824, w_000_825, w_000_826, w_000_827, w_000_828, w_000_829, w_000_830, w_000_831, w_000_832, w_000_833, w_000_834, w_000_835, w_000_836, w_000_837, w_000_838, w_000_839, w_000_840, w_000_841, w_000_842, w_000_843, w_000_844, w_000_845, w_000_846, w_000_847, w_000_848, w_000_849, w_000_850, w_000_851, w_000_852, w_000_853, w_000_854, w_000_855, w_000_856, w_000_857, w_000_858, w_000_859, w_000_860, w_000_861, w_000_862, w_000_863, w_000_864, w_000_865, w_000_866, w_000_867, w_000_868, w_000_869, w_000_870, w_000_871, w_000_872, w_000_873, w_000_874, w_000_875, w_000_876, w_000_877, w_000_878, w_000_879, w_000_880, w_000_881, w_000_882, w_000_883, w_000_885, w_000_886, w_000_887, w_000_889, w_000_890, w_000_891, w_000_893, w_000_894, w_000_895, w_000_896, w_000_897, w_000_898, w_000_899, w_000_900, w_000_901, w_000_903, w_000_904, w_000_905, w_000_906, w_000_907, w_000_908, w_000_909, w_000_910, w_000_912, w_000_914, w_000_915, w_000_916, w_000_917, w_000_918, w_000_919, w_000_923, w_000_924, w_000_925, w_000_926, w_000_928, w_000_929, w_000_930, w_000_931, w_000_932, w_000_934, w_000_935, w_000_936, w_000_937, w_000_938, w_000_939, w_000_943, w_000_944, w_000_945, w_000_947, w_000_949, w_000_950, w_000_952, w_000_953, w_000_954, w_000_955, w_000_956, w_000_958, w_000_959, w_000_960, w_000_963, w_000_964, w_000_965, w_000_967, w_000_968, w_000_969, w_000_970, w_000_971, w_000_977, w_000_979, w_000_980, w_000_981, w_000_982, w_000_983, w_1000_000, w_1000_001, w_1000_002, w_1000_003, w_1000_004, w_1000_005, w_1000_006, w_1000_007, w_1000_008, w_1000_009, w_1000_010, w_1000_011, w_1000_012, w_1000_013, w_1000_014, w_1000_015, w_1000_016, w_1000_017, w_1000_018, w_1000_019, w_1000_020, w_1000_021, w_1000_022, w_1000_023, w_1000_024, w_1000_025, w_1000_026, w_1000_027, w_1000_028, w_1000_029, w_1000_030, w_1000_031, w_1000_032, w_1000_033, w_1000_034, w_1000_035, w_1000_036, w_1000_037, w_1000_038, w_1000_039, w_1000_040, w_1000_041, w_1000_042, w_1000_043, w_1000_044, w_1000_045, w_1000_046, w_1000_047, w_1000_048, w_1000_049, w_1000_050, w_1000_051, w_1000_052, w_1000_053, w_1000_054, w_1000_055, w_1000_056, w_1000_057, w_1000_058, w_1000_059, w_1000_060, w_1000_061, w_1000_062, w_1000_063, w_1000_064, w_1000_065, w_1000_066, w_1000_067, w_1000_068, w_1000_069, w_1000_070, w_1000_071, w_1000_072, w_1000_073, w_1000_074, w_1000_075, w_1000_076, w_1000_077, w_1000_078, w_1000_079, w_1000_080, w_1000_081, w_1000_082, w_1000_083, w_1000_084, w_1000_085, w_1000_086, w_1000_087, w_1000_088, w_1000_089, w_1000_090, w_1000_091, w_1000_092, w_1000_093, w_1000_094, w_1000_095, w_1000_096, w_1000_097, w_1000_098, w_1000_099, w_1000_100, w_1000_101, w_1000_102, w_1000_103, w_1000_104, w_1000_105, w_1000_106, w_1000_107, w_1000_108, w_1000_109, w_1000_110, w_1000_111, w_1000_112, w_1000_113, w_1000_114, w_1000_115, w_1000_116, w_1000_117, w_1000_118, w_1000_119, w_1000_120, w_1000_121, w_1000_122, w_1000_123, w_1000_124, w_1000_125, w_1000_126, w_1000_127, w_1000_128, w_1000_129, w_1000_130, w_1000_131, w_1000_132, w_1000_133, w_1000_134, w_1000_135, w_1000_136, w_1000_137, w_1000_138, w_1000_139, w_1000_140, w_1000_141, w_1000_142, w_1000_143, w_1000_144, w_1000_145, w_1000_146, w_1000_147, w_1000_148, w_1000_149, w_1000_150, w_1000_151, w_1000_152, w_1000_153, w_1000_154, w_1000_155, w_1000_156, w_1000_157, w_1000_158, w_1000_159, w_1000_160, w_1000_161, w_1000_162, w_1000_163, w_1000_164, w_1000_165, w_1000_166, w_1000_167, w_1000_168, w_1000_169, w_1000_170, w_1000_171, w_1000_172, w_1000_173, w_1000_174, w_1000_175, w_1000_176, w_1000_177, w_1000_178, w_1000_179, w_1000_180, w_1000_181, w_1000_182, w_1000_183, w_1000_184, w_1000_185 ;
  combLogic I0(  w_000_000, w_000_001, w_000_002, w_000_003, w_000_004, w_000_005, w_000_006, w_000_007, w_000_008, w_000_009, w_000_010, w_000_011, w_000_012, w_000_013, w_000_014, w_000_015, w_000_016, w_000_017, w_000_018, w_000_019, w_000_020, w_000_021, w_000_022, w_000_023, w_000_024, w_000_025, w_000_026, w_000_027, w_000_028, w_000_029, w_000_030, w_000_031, w_000_032, w_000_033, w_000_034, w_000_035, w_000_036, w_000_037, w_000_038, w_000_039, w_000_040, w_000_041, w_000_042, w_000_043, w_000_044, w_000_045, w_000_046, w_000_047, w_000_048, w_000_049, w_000_050, w_000_051, w_000_052, w_000_053, w_000_054, w_000_055, w_000_056, w_000_057, w_000_058, w_000_059, w_000_060, w_000_061, w_000_062, w_000_063, w_000_064, w_000_065, w_000_066, w_000_067, w_000_068, w_000_069, w_000_070, w_000_071, w_000_072, w_000_073, w_000_074, w_000_075, w_000_076, w_000_077, w_000_078, w_000_079, w_000_080, w_000_081, w_000_082, w_000_083, w_000_084, w_000_085, w_000_086, w_000_087, w_000_088, w_000_089, w_000_090, w_000_091, w_000_092, w_000_093, w_000_094, w_000_095, w_000_096, w_000_097, w_000_098, w_000_099, w_000_100, w_000_101, w_000_102, w_000_103, w_000_104, w_000_105, w_000_106, w_000_107, w_000_108, w_000_109, w_000_110, w_000_111, w_000_112, w_000_113, w_000_114, w_000_115, w_000_116, w_000_117, w_000_118, w_000_119, w_000_120, w_000_121, w_000_122, w_000_123, w_000_124, w_000_125, w_000_126, w_000_127, w_000_128, w_000_129, w_000_130, w_000_131, w_000_132, w_000_133, w_000_134, w_000_135, w_000_136, w_000_137, w_000_138, w_000_139, w_000_140, w_000_141, w_000_142, w_000_143, w_000_144, w_000_145, w_000_146, w_000_147, w_000_148, w_000_149, w_000_150, w_000_151, w_000_152, w_000_153, w_000_154, w_000_155, w_000_156, w_000_157, w_000_158, w_000_159, w_000_160, w_000_161, w_000_162, w_000_163, w_000_164, w_000_165, w_000_166, w_000_167, w_000_168, w_000_169, w_000_170, w_000_171, w_000_172, w_000_173, w_000_174, w_000_175, w_000_176, w_000_177, w_000_178, w_000_179, w_000_180, w_000_181, w_000_182, w_000_183, w_000_184, w_000_185, w_000_186, w_000_187, w_000_188, w_000_189, w_000_190, w_000_191, w_000_192, w_000_193, w_000_194, w_000_195, w_000_196, w_000_197, w_000_198, w_000_199, w_000_200, w_000_201, w_000_202, w_000_203, w_000_204, w_000_205, w_000_206, w_000_207, w_000_208, w_000_209, w_000_210, w_000_211, w_000_212, w_000_213, w_000_214, w_000_215, w_000_216, w_000_217, w_000_218, w_000_219, w_000_220, w_000_221, w_000_222, w_000_223, w_000_224, w_000_225, w_000_226, w_000_227, w_000_228, w_000_230, w_000_231, w_000_232, w_000_233, w_000_234, w_000_235, w_000_236, w_000_237, w_000_238, w_000_239, w_000_240, w_000_241, w_000_242, w_000_243, w_000_244, w_000_245, w_000_246, w_000_247, w_000_248, w_000_249, w_000_250, w_000_251, w_000_252, w_000_253, w_000_254, w_000_255, w_000_256, w_000_257, w_000_258, w_000_259, w_000_260, w_000_262, w_000_263, w_000_264, w_000_265, w_000_266, w_000_267, w_000_268, w_000_269, w_000_270, w_000_271, w_000_272, w_000_273, w_000_274, w_000_275, w_000_276, w_000_277, w_000_278, w_000_279, w_000_280, w_000_281, w_000_282, w_000_283, w_000_284, w_000_285, w_000_286, w_000_287, w_000_288, w_000_289, w_000_290, w_000_291, w_000_292, w_000_293, w_000_294, w_000_295, w_000_296, w_000_297, w_000_298, w_000_299, w_000_300, w_000_301, w_000_302, w_000_303, w_000_304, w_000_305, w_000_306, w_000_307, w_000_308, w_000_309, w_000_310, w_000_311, w_000_312, w_000_313, w_000_314, w_000_315, w_000_316, w_000_317, w_000_318, w_000_319, w_000_320, w_000_321, w_000_322, w_000_323, w_000_324, w_000_325, w_000_326, w_000_327, w_000_328, w_000_329, w_000_330, w_000_331, w_000_332, w_000_333, w_000_334, w_000_335, w_000_336, w_000_337, w_000_338, w_000_339, w_000_340, w_000_341, w_000_342, w_000_343, w_000_344, w_000_345, w_000_346, w_000_347, w_000_348, w_000_349, w_000_350, w_000_351, w_000_352, w_000_353, w_000_354, w_000_355, w_000_356, w_000_357, w_000_358, w_000_359, w_000_360, w_000_361, w_000_362, w_000_364, w_000_365, w_000_366, w_000_367, w_000_369, w_000_370, w_000_371, w_000_372, w_000_373, w_000_374, w_000_375, w_000_376, w_000_377, w_000_378, w_000_379, w_000_380, w_000_381, w_000_382, w_000_383, w_000_384, w_000_385, w_000_386, w_000_387, w_000_388, w_000_389, w_000_390, w_000_391, w_000_392, w_000_393, w_000_394, w_000_395, w_000_396, w_000_397, w_000_398, w_000_399, w_000_400, w_000_401, w_000_402, w_000_403, w_000_404, w_000_405, w_000_406, w_000_407, w_000_408, w_000_409, w_000_410, w_000_411, w_000_412, w_000_413, w_000_414, w_000_415, w_000_416, w_000_417, w_000_418, w_000_419, w_000_420, w_000_421, w_000_422, w_000_423, w_000_424, w_000_425, w_000_426, w_000_427, w_000_428, w_000_429, w_000_430, w_000_431, w_000_432, w_000_433, w_000_434, w_000_435, w_000_436, w_000_437, w_000_438, w_000_439, w_000_440, w_000_441, w_000_442, w_000_443, w_000_444, w_000_445, w_000_446, w_000_447, w_000_448, w_000_449, w_000_450, w_000_451, w_000_452, w_000_453, w_000_454, w_000_455, w_000_456, w_000_457, w_000_458, w_000_459, w_000_460, w_000_461, w_000_462, w_000_463, w_000_464, w_000_465, w_000_466, w_000_467, w_000_468, w_000_469, w_000_470, w_000_471, w_000_472, w_000_473, w_000_474, w_000_475, w_000_476, w_000_477, w_000_478, w_000_479, w_000_480, w_000_481, w_000_482, w_000_483, w_000_484, w_000_485, w_000_486, w_000_487, w_000_488, w_000_489, w_000_490, w_000_491, w_000_492, w_000_493, w_000_494, w_000_495, w_000_496, w_000_497, w_000_498, w_000_499, w_000_500, w_000_501, w_000_502, w_000_503, w_000_504, w_000_505, w_000_506, w_000_507, w_000_508, w_000_509, w_000_510, w_000_511, w_000_512, w_000_513, w_000_514, w_000_515, w_000_516, w_000_517, w_000_518, w_000_519, w_000_520, w_000_521, w_000_522, w_000_523, w_000_524, w_000_525, w_000_526, w_000_527, w_000_528, w_000_529, w_000_530, w_000_531, w_000_532, w_000_533, w_000_534, w_000_535, w_000_536, w_000_537, w_000_538, w_000_539, w_000_540, w_000_541, w_000_542, w_000_543, w_000_544, w_000_545, w_000_546, w_000_547, w_000_548, w_000_549, w_000_550, w_000_551, w_000_552, w_000_553, w_000_554, w_000_555, w_000_556, w_000_557, w_000_558, w_000_559, w_000_560, w_000_561, w_000_562, w_000_563, w_000_564, w_000_565, w_000_566, w_000_567, w_000_568, w_000_569, w_000_570, w_000_571, w_000_572, w_000_573, w_000_574, w_000_575, w_000_576, w_000_577, w_000_578, w_000_579, w_000_580, w_000_581, w_000_582, w_000_583, w_000_584, w_000_585, w_000_586, w_000_587, w_000_588, w_000_589, w_000_590, w_000_591, w_000_592, w_000_593, w_000_594, w_000_595, w_000_596, w_000_597, w_000_598, w_000_599, w_000_600, w_000_601, w_000_602, w_000_603, w_000_604, w_000_605, w_000_606, w_000_607, w_000_608, w_000_609, w_000_610, w_000_611, w_000_612, w_000_613, w_000_614, w_000_615, w_000_616, w_000_617, w_000_618, w_000_619, w_000_620, w_000_621, w_000_622, w_000_623, w_000_624, w_000_625, w_000_626, w_000_627, w_000_628, w_000_629, w_000_630, w_000_631, w_000_632, w_000_633, w_000_634, w_000_635, w_000_636, w_000_637, w_000_638, w_000_639, w_000_640, w_000_641, w_000_642, w_000_643, w_000_644, w_000_645, w_000_646, w_000_647, w_000_648, w_000_649, w_000_650, w_000_651, w_000_652, w_000_653, w_000_654, w_000_655, w_000_656, w_000_657, w_000_658, w_000_659, w_000_660, w_000_661, w_000_662, w_000_663, w_000_664, w_000_665, w_000_666, w_000_667, w_000_669, w_000_670, w_000_671, w_000_672, w_000_673, w_000_674, w_000_675, w_000_676, w_000_677, w_000_678, w_000_679, w_000_680, w_000_681, w_000_682, w_000_683, w_000_684, w_000_685, w_000_686, w_000_687, w_000_688, w_000_689, w_000_690, w_000_691, w_000_692, w_000_693, w_000_694, w_000_695, w_000_696, w_000_697, w_000_698, w_000_699, w_000_700, w_000_701, w_000_702, w_000_703, w_000_704, w_000_705, w_000_706, w_000_707, w_000_708, w_000_709, w_000_710, w_000_711, w_000_712, w_000_713, w_000_714, w_000_715, w_000_716, w_000_717, w_000_718, w_000_719, w_000_720, w_000_721, w_000_722, w_000_723, w_000_724, w_000_725, w_000_726, w_000_727, w_000_728, w_000_729, w_000_730, w_000_731, w_000_732, w_000_733, w_000_734, w_000_735, w_000_736, w_000_737, w_000_738, w_000_739, w_000_740, w_000_741, w_000_742, w_000_743, w_000_744, w_000_745, w_000_746, w_000_747, w_000_748, w_000_749, w_000_750, w_000_751, w_000_752, w_000_753, w_000_754, w_000_755, w_000_756, w_000_757, w_000_758, w_000_759, w_000_760, w_000_761, w_000_762, w_000_763, w_000_765, w_000_766, w_000_767, w_000_769, w_000_770, w_000_772, w_000_773, w_000_774, w_000_775, w_000_776, w_000_777, w_000_779, w_000_780, w_000_781, w_000_782, w_000_783, w_000_784, w_000_785, w_000_786, w_000_787, w_000_788, w_000_789, w_000_790, w_000_791, w_000_792, w_000_793, w_000_794, w_000_795, w_000_796, w_000_797, w_000_798, w_000_799, w_000_801, w_000_802, w_000_803, w_000_804, w_000_805, w_000_806, w_000_807, w_000_808, w_000_809, w_000_810, w_000_811, w_000_812, w_000_813, w_000_814, w_000_815, w_000_816, w_000_817, w_000_818, w_000_819, w_000_820, w_000_821, w_000_822, w_000_823, w_000_824, w_000_825, w_000_826, w_000_827, w_000_828, w_000_829, w_000_830, w_000_831, w_000_832, w_000_833, w_000_834, w_000_835, w_000_836, w_000_837, w_000_838, w_000_839, w_000_840, w_000_841, w_000_842, w_000_843, w_000_844, w_000_845, w_000_846, w_000_847, w_000_848, w_000_849, w_000_850, w_000_851, w_000_852, w_000_853, w_000_854, w_000_855, w_000_856, w_000_857, w_000_858, w_000_859, w_000_860, w_000_861, w_000_862, w_000_863, w_000_864, w_000_865, w_000_866, w_000_867, w_000_868, w_000_869, w_000_870, w_000_871, w_000_872, w_000_873, w_000_874, w_000_875, w_000_876, w_000_877, w_000_878, w_000_879, w_000_880, w_000_881, w_000_882, w_000_883, w_000_885, w_000_886, w_000_887, w_000_889, w_000_890, w_000_891, w_000_893, w_000_894, w_000_895, w_000_896, w_000_897, w_000_898, w_000_899, w_000_900, w_000_901, w_000_903, w_000_904, w_000_905, w_000_906, w_000_907, w_000_908, w_000_909, w_000_910, w_000_912, w_000_914, w_000_915, w_000_916, w_000_917, w_000_918, w_000_919, w_000_923, w_000_924, w_000_925, w_000_926, w_000_928, w_000_929, w_000_930, w_000_931, w_000_932, w_000_934, w_000_935, w_000_936, w_000_937, w_000_938, w_000_939, w_000_943, w_000_944, w_000_945, w_000_947, w_000_949, w_000_950, w_000_952, w_000_953, w_000_954, w_000_955, w_000_956, w_000_958, w_000_959, w_000_960, w_000_963, w_000_964, w_000_965, w_000_967, w_000_968, w_000_969, w_000_970, w_000_971, w_000_977, w_000_979, w_000_980, w_000_981, w_000_982, w_000_983, w_1000_000, w_1000_001, w_1000_002, w_1000_003, w_1000_004, w_1000_005, w_1000_006, w_1000_007, w_1000_008, w_1000_009, w_1000_010, w_1000_011, w_1000_012, w_1000_013, w_1000_014, w_1000_015, w_1000_016, w_1000_017, w_1000_018, w_1000_019, w_1000_020, w_1000_021, w_1000_022, w_1000_023, w_1000_024, w_1000_025, w_1000_026, w_1000_027, w_1000_028, w_1000_029, w_1000_030, w_1000_031, w_1000_032, w_1000_033, w_1000_034, w_1000_035, w_1000_036, w_1000_037, w_1000_038, w_1000_039, w_1000_040, w_1000_041, w_1000_042, w_1000_043, w_1000_044, w_1000_045, w_1000_046, w_1000_047, w_1000_048, w_1000_049, w_1000_050, w_1000_051, w_1000_052, w_1000_053, w_1000_054, w_1000_055, w_1000_056, w_1000_057, w_1000_058, w_1000_059, w_1000_060, w_1000_061, w_1000_062, w_1000_063, w_1000_064, w_1000_065, w_1000_066, w_1000_067, w_1000_068, w_1000_069, w_1000_070, w_1000_071, w_1000_072, w_1000_073, w_1000_074, w_1000_075, w_1000_076, w_1000_077, w_1000_078, w_1000_079, w_1000_080, w_1000_081, w_1000_082, w_1000_083, w_1000_084, w_1000_085, w_1000_086, w_1000_087, w_1000_088, w_1000_089, w_1000_090, w_1000_091, w_1000_092, w_1000_093, w_1000_094, w_1000_095, w_1000_096, w_1000_097, w_1000_098, w_1000_099, w_1000_100, w_1000_101, w_1000_102, w_1000_103, w_1000_104, w_1000_105, w_1000_106, w_1000_107, w_1000_108, w_1000_109, w_1000_110, w_1000_111, w_1000_112, w_1000_113, w_1000_114, w_1000_115, w_1000_116, w_1000_117, w_1000_118, w_1000_119, w_1000_120, w_1000_121, w_1000_122, w_1000_123, w_1000_124, w_1000_125, w_1000_126, w_1000_127, w_1000_128, w_1000_129, w_1000_130, w_1000_131, w_1000_132, w_1000_133, w_1000_134, w_1000_135, w_1000_136, w_1000_137, w_1000_138, w_1000_139, w_1000_140, w_1000_141, w_1000_142, w_1000_143, w_1000_144, w_1000_145, w_1000_146, w_1000_147, w_1000_148, w_1000_149, w_1000_150, w_1000_151, w_1000_152, w_1000_153, w_1000_154, w_1000_155, w_1000_156, w_1000_157, w_1000_158, w_1000_159, w_1000_160, w_1000_161, w_1000_162, w_1000_163, w_1000_164, w_1000_165, w_1000_166, w_1000_167, w_1000_168, w_1000_169, w_1000_170, w_1000_171, w_1000_172, w_1000_173, w_1000_174, w_1000_175, w_1000_176, w_1000_177, w_1000_178, w_1000_179, w_1000_180, w_1000_181, w_1000_182, w_1000_183, w_1000_184, w_1000_185  );

  reg r0, r1, r2, r3, r4, r5, r6, r7, r8, r9, r10, r11, r12, r13, r14, r15, r16, r17, r18, r19, r20, r21, r22, r23, r24, r25, r26, r27, r28, r29, r30, r31, r32, r33, r34, r35, r36, r37, r38, r39, r40, r41, r42, r43, r44, r45, r46, r47, r48, r49, r50, r51, r52, r53, r54, r55, r56, r57, r58, r59, r60, r61, r62, r63, r64, r65, r66, r67, r68, r69, r70, r71, r72, r73, r74, r75, r76, r77, r78, r79, r80, r81, r82, r83, r84, r85, r86, r87, r88, r89, r90, r91, r92, r93, r94, r95, r96, r97, r98, r99, r100, r101, r102, r103, r104, r105, r106, r107, r108, r109, r110, r111, r112, r113, r114, r115, r116, r117, r118, r119, r120, r121, r122, r123, r124, r125, r126, r127, r128, r129, r130, r131, r132, r133, r134, r135, r136, r137, r138, r139, r140, r141, r142, r143, r144, r145, r146, r147, r148, r149, r150, r151, r152, r153, r154, r155, r156, r157, r158, r159, r160, r161, r162, r163, r164, r165, r166, r167, r168, r169, r170, r171, r172, r173, r174, r175, r176, r177, r178, r179, r180, r181, r182, r183, r184, r185, r186, r187, r188, r189, r190, r191, r192, r193, r194, r195, r196, r197, r198, r199, r200, r201, r202, r203, r204, r205, r206, r207, r208, r209, r210, r211, r212, r213, r214, r215, r216, r217, r218, r219, r220, r221, r222, r223, r224, r225, r226, r227, r228, r229, r230, r231, r232, r233, r234, r235, r236, r237, r238, r239, r240, r241, r242, r243, r244, r245, r246, r247, r248, r249, r250, r251, r252, r253, r254, r255, r256, r257, r258, r259, r260, r261, r262, r263, r264, r265, r266, r267, r268, r269, r270, r271, r272, r273, r274, r275, r276, r277, r278, r279, r280, r281, r282, r283, r284, r285, r286, r287, r288, r289, r290, r291, r292, r293, r294, r295, r296, r297, r298, r299, r300, r301, r302, r303, r304, r305, r306, r307, r308, r309, r310, r311, r312, r313, r314, r315, r316, r317, r318, r319, r320, r321, r322, r323, r324, r325, r326, r327, r328, r329, r330, r331, r332, r333, r334, r335, r336, r337, r338, r339, r340, r341, r342, r343, r344, r345, r346, r347, r348, r349, r350, r351, r352, r353, r354, r355, r356, r357, r358, r359, r360, r361, r362, r363, r364, r365, r366, r367, r368, r369, r370, r371, r372, r373, r374, r375, r376, r377, r378, r379, r380, r381, r382, r383, r384, r385, r386, r387, r388, r389, r390, r391, r392, r393, r394, r395, r396, r397, r398, r399, r400, r401, r402, r403, r404, r405, r406, r407, r408, r409, r410, r411, r412, r413, r414, r415, r416, r417, r418, r419, r420, r421, r422, r423, r424, r425, r426, r427, r428, r429, r430, r431, r432, r433, r434, r435, r436, r437, r438, r439, r440, r441, r442, r443, r444, r445, r446, r447, r448, r449, r450, r451, r452, r453, r454, r455, r456, r457, r458, r459, r460, r461, r462, r463, r464, r465, r466, r467, r468, r469, r470, r471, r472, r473, r474, r475, r476, r477, r478, r479, r480, r481, r482, r483, r484, r485, r486, r487, r488, r489, r490, r491, r492, r493, r494, r495, r496, r497, r498, r499, r500, r501, r502, r503, r504, r505, r506, r507, r508, r509, r510, r511, r512, r513, r514, r515, r516, r517, r518, r519, r520, r521, r522, r523, r524, r525, r526, r527, r528, r529, r530, r531, r532, r533, r534, r535, r536, r537, r538, r539, r540, r541, r542, r543, r544, r545, r546, r547, r548, r549, r550, r551, r552, r553, r554, r555, r556, r557, r558, r559, r560, r561, r562, r563, r564, r565, r566, r567, r568, r569, r570, r571, r572, r573, r574, r575, r576, r577, r578, r579, r580, r581, r582, r583, r584, r585, r586, r587, r588, r589, r590, r591, r592, r593, r594, r595, r596, r597, r598, r599, r600, r601, r602, r603, r604, r605, r606, r607, r608, r609, r610, r611, r612, r613, r614, r615, r616, r617, r618, r619, r620, r621, r622, r623, r624, r625, r626, r627, r628, r629, r630, r631, r632, r633, r634, r635, r636, r637, r638, r639, r640, r641, r642, r643, r644, r645, r646, r647, r648, r649, r650, r651, r652, r653, r654, r655, r656, r657, r658, r659, r660, r661, r662, r663, r664, r665, r666, r667, r668, r669, r670, r671, r672, r673, r674, r675, r676, r677, r678, r679, r680, r681, r682, r683, r684, r685, r686, r687, r688, r689, r690, r691, r692, r693, r694, r695, r696, r697, r698, r699, r700, r701, r702, r703, r704, r705, r706, r707, r708, r709, r710, r711, r712, r713, r714, r715, r716, r717, r718, r719, r720, r721, r722, r723, r724, r725, r726, r727, r728, r729, r730, r731, r732, r733, r734, r735, r736, r737, r738, r739, r740, r741, r742, r743, r744, r745, r746, r747, r748, r749, r750, r751, r752, r753, r754, r755, r756, r757, r758, r759, r760, r761, r762, r763, r764, r765, r766, r767, r768, r769, r770, r771, r772, r773, r774, r775, r776, r777, r778, r779, r780, r781, r782, r783, r784, r785, r786, r787, r788, r789, r790, r791, r792, r793, r794, r795, r796, r797, r798, r799, r800, r801, r802, r803, r804, r805, r806, r807, r808, r809, r810, r811, r812, r813, r814, r815, r816, r817, r818, r819, r820, r821, r822, r823, r824, r825, r826, r827, r828, r829, r830, r831, r832, r833, r834, r835, r836, r837, r838, r839, r840, r841, r842, r843, r844, r845, r846, r847, r848, r849, r850, r851, r852, r853, r854, r855, r856, r857, r858, r859, r860, r861, r862, r863, r864, r865, r866, r867, r868, r869, r870, r871, r872, r873, r874, r875, r876, r877, r878, r879, r880, r881, r882, r883, r884, r885, r886, r887, r888, r889, r890, r891, r892, r893, r894, r895, r896, r897, r898, r899, r900, r901, r902, r903, r904, r905, r906, r907, r908, r909, r910, r911, r912, r913, r914, r915, r916, r917, r918, r919, r920, r921, r922, r923, r924, r925, r926, r927, r928, r929, r930, r931, r932, r933, r934, r935, r936, r937, r938, r939, r940, r941, r942, r943, r944, r945, r946, r947, r948, r949, r950, r951, r952, r953, r954, r955, r956, r957, r958, r959, r960, r961, r962, r963, r964, r965, r966, r967, r968, r969, r970, r971, r972, r973, r974, r975, r976, r977, r978, r979, r980, r981, r982, r983, r984, r985, r986, r987, r988, r989, r990, r991, r992, r993, r994, r995, r996, r997, r998, r999, rEnd; 

  assign w_000_000 = r0;
  assign w_000_001 = r1;
  assign w_000_002 = r2;
  assign w_000_003 = r3;
  assign w_000_004 = r4;
  assign w_000_005 = r5;
  assign w_000_006 = r6;
  assign w_000_007 = r7;
  assign w_000_008 = r8;
  assign w_000_009 = r9;
  assign w_000_010 = r10;
  assign w_000_011 = r11;
  assign w_000_012 = r12;
  assign w_000_013 = r13;
  assign w_000_014 = r14;
  assign w_000_015 = r15;
  assign w_000_016 = r16;
  assign w_000_017 = r17;
  assign w_000_018 = r18;
  assign w_000_019 = r19;
  assign w_000_020 = r20;
  assign w_000_021 = r21;
  assign w_000_022 = r22;
  assign w_000_023 = r23;
  assign w_000_024 = r24;
  assign w_000_025 = r25;
  assign w_000_026 = r26;
  assign w_000_027 = r27;
  assign w_000_028 = r28;
  assign w_000_029 = r29;
  assign w_000_030 = r30;
  assign w_000_031 = r31;
  assign w_000_032 = r32;
  assign w_000_033 = r33;
  assign w_000_034 = r34;
  assign w_000_035 = r35;
  assign w_000_036 = r36;
  assign w_000_037 = r37;
  assign w_000_038 = r38;
  assign w_000_039 = r39;
  assign w_000_040 = r40;
  assign w_000_041 = r41;
  assign w_000_042 = r42;
  assign w_000_043 = r43;
  assign w_000_044 = r44;
  assign w_000_045 = r45;
  assign w_000_046 = r46;
  assign w_000_047 = r47;
  assign w_000_048 = r48;
  assign w_000_049 = r49;
  assign w_000_050 = r50;
  assign w_000_051 = r51;
  assign w_000_052 = r52;
  assign w_000_053 = r53;
  assign w_000_054 = r54;
  assign w_000_055 = r55;
  assign w_000_056 = r56;
  assign w_000_057 = r57;
  assign w_000_058 = r58;
  assign w_000_059 = r59;
  assign w_000_060 = r60;
  assign w_000_061 = r61;
  assign w_000_062 = r62;
  assign w_000_063 = r63;
  assign w_000_064 = r64;
  assign w_000_065 = r65;
  assign w_000_066 = r66;
  assign w_000_067 = r67;
  assign w_000_068 = r68;
  assign w_000_069 = r69;
  assign w_000_070 = r70;
  assign w_000_071 = r71;
  assign w_000_072 = r72;
  assign w_000_073 = r73;
  assign w_000_074 = r74;
  assign w_000_075 = r75;
  assign w_000_076 = r76;
  assign w_000_077 = r77;
  assign w_000_078 = r78;
  assign w_000_079 = r79;
  assign w_000_080 = r80;
  assign w_000_081 = r81;
  assign w_000_082 = r82;
  assign w_000_083 = r83;
  assign w_000_084 = r84;
  assign w_000_085 = r85;
  assign w_000_086 = r86;
  assign w_000_087 = r87;
  assign w_000_088 = r88;
  assign w_000_089 = r89;
  assign w_000_090 = r90;
  assign w_000_091 = r91;
  assign w_000_092 = r92;
  assign w_000_093 = r93;
  assign w_000_094 = r94;
  assign w_000_095 = r95;
  assign w_000_096 = r96;
  assign w_000_097 = r97;
  assign w_000_098 = r98;
  assign w_000_099 = r99;
  assign w_000_100 = r100;
  assign w_000_101 = r101;
  assign w_000_102 = r102;
  assign w_000_103 = r103;
  assign w_000_104 = r104;
  assign w_000_105 = r105;
  assign w_000_106 = r106;
  assign w_000_107 = r107;
  assign w_000_108 = r108;
  assign w_000_109 = r109;
  assign w_000_110 = r110;
  assign w_000_111 = r111;
  assign w_000_112 = r112;
  assign w_000_113 = r113;
  assign w_000_114 = r114;
  assign w_000_115 = r115;
  assign w_000_116 = r116;
  assign w_000_117 = r117;
  assign w_000_118 = r118;
  assign w_000_119 = r119;
  assign w_000_120 = r120;
  assign w_000_121 = r121;
  assign w_000_122 = r122;
  assign w_000_123 = r123;
  assign w_000_124 = r124;
  assign w_000_125 = r125;
  assign w_000_126 = r126;
  assign w_000_127 = r127;
  assign w_000_128 = r128;
  assign w_000_129 = r129;
  assign w_000_130 = r130;
  assign w_000_131 = r131;
  assign w_000_132 = r132;
  assign w_000_133 = r133;
  assign w_000_134 = r134;
  assign w_000_135 = r135;
  assign w_000_136 = r136;
  assign w_000_137 = r137;
  assign w_000_138 = r138;
  assign w_000_139 = r139;
  assign w_000_140 = r140;
  assign w_000_141 = r141;
  assign w_000_142 = r142;
  assign w_000_143 = r143;
  assign w_000_144 = r144;
  assign w_000_145 = r145;
  assign w_000_146 = r146;
  assign w_000_147 = r147;
  assign w_000_148 = r148;
  assign w_000_149 = r149;
  assign w_000_150 = r150;
  assign w_000_151 = r151;
  assign w_000_152 = r152;
  assign w_000_153 = r153;
  assign w_000_154 = r154;
  assign w_000_155 = r155;
  assign w_000_156 = r156;
  assign w_000_157 = r157;
  assign w_000_158 = r158;
  assign w_000_159 = r159;
  assign w_000_160 = r160;
  assign w_000_161 = r161;
  assign w_000_162 = r162;
  assign w_000_163 = r163;
  assign w_000_164 = r164;
  assign w_000_165 = r165;
  assign w_000_166 = r166;
  assign w_000_167 = r167;
  assign w_000_168 = r168;
  assign w_000_169 = r169;
  assign w_000_170 = r170;
  assign w_000_171 = r171;
  assign w_000_172 = r172;
  assign w_000_173 = r173;
  assign w_000_174 = r174;
  assign w_000_175 = r175;
  assign w_000_176 = r176;
  assign w_000_177 = r177;
  assign w_000_178 = r178;
  assign w_000_179 = r179;
  assign w_000_180 = r180;
  assign w_000_181 = r181;
  assign w_000_182 = r182;
  assign w_000_183 = r183;
  assign w_000_184 = r184;
  assign w_000_185 = r185;
  assign w_000_186 = r186;
  assign w_000_187 = r187;
  assign w_000_188 = r188;
  assign w_000_189 = r189;
  assign w_000_190 = r190;
  assign w_000_191 = r191;
  assign w_000_192 = r192;
  assign w_000_193 = r193;
  assign w_000_194 = r194;
  assign w_000_195 = r195;
  assign w_000_196 = r196;
  assign w_000_197 = r197;
  assign w_000_198 = r198;
  assign w_000_199 = r199;
  assign w_000_200 = r200;
  assign w_000_201 = r201;
  assign w_000_202 = r202;
  assign w_000_203 = r203;
  assign w_000_204 = r204;
  assign w_000_205 = r205;
  assign w_000_206 = r206;
  assign w_000_207 = r207;
  assign w_000_208 = r208;
  assign w_000_209 = r209;
  assign w_000_210 = r210;
  assign w_000_211 = r211;
  assign w_000_212 = r212;
  assign w_000_213 = r213;
  assign w_000_214 = r214;
  assign w_000_215 = r215;
  assign w_000_216 = r216;
  assign w_000_217 = r217;
  assign w_000_218 = r218;
  assign w_000_219 = r219;
  assign w_000_220 = r220;
  assign w_000_221 = r221;
  assign w_000_222 = r222;
  assign w_000_223 = r223;
  assign w_000_224 = r224;
  assign w_000_225 = r225;
  assign w_000_226 = r226;
  assign w_000_227 = r227;
  assign w_000_228 = r228;
  assign w_000_229 = r229;
  assign w_000_230 = r230;
  assign w_000_231 = r231;
  assign w_000_232 = r232;
  assign w_000_233 = r233;
  assign w_000_234 = r234;
  assign w_000_235 = r235;
  assign w_000_236 = r236;
  assign w_000_237 = r237;
  assign w_000_238 = r238;
  assign w_000_239 = r239;
  assign w_000_240 = r240;
  assign w_000_241 = r241;
  assign w_000_242 = r242;
  assign w_000_243 = r243;
  assign w_000_244 = r244;
  assign w_000_245 = r245;
  assign w_000_246 = r246;
  assign w_000_247 = r247;
  assign w_000_248 = r248;
  assign w_000_249 = r249;
  assign w_000_250 = r250;
  assign w_000_251 = r251;
  assign w_000_252 = r252;
  assign w_000_253 = r253;
  assign w_000_254 = r254;
  assign w_000_255 = r255;
  assign w_000_256 = r256;
  assign w_000_257 = r257;
  assign w_000_258 = r258;
  assign w_000_259 = r259;
  assign w_000_260 = r260;
  assign w_000_261 = r261;
  assign w_000_262 = r262;
  assign w_000_263 = r263;
  assign w_000_264 = r264;
  assign w_000_265 = r265;
  assign w_000_266 = r266;
  assign w_000_267 = r267;
  assign w_000_268 = r268;
  assign w_000_269 = r269;
  assign w_000_270 = r270;
  assign w_000_271 = r271;
  assign w_000_272 = r272;
  assign w_000_273 = r273;
  assign w_000_274 = r274;
  assign w_000_275 = r275;
  assign w_000_276 = r276;
  assign w_000_277 = r277;
  assign w_000_278 = r278;
  assign w_000_279 = r279;
  assign w_000_280 = r280;
  assign w_000_281 = r281;
  assign w_000_282 = r282;
  assign w_000_283 = r283;
  assign w_000_284 = r284;
  assign w_000_285 = r285;
  assign w_000_286 = r286;
  assign w_000_287 = r287;
  assign w_000_288 = r288;
  assign w_000_289 = r289;
  assign w_000_290 = r290;
  assign w_000_291 = r291;
  assign w_000_292 = r292;
  assign w_000_293 = r293;
  assign w_000_294 = r294;
  assign w_000_295 = r295;
  assign w_000_296 = r296;
  assign w_000_297 = r297;
  assign w_000_298 = r298;
  assign w_000_299 = r299;
  assign w_000_300 = r300;
  assign w_000_301 = r301;
  assign w_000_302 = r302;
  assign w_000_303 = r303;
  assign w_000_304 = r304;
  assign w_000_305 = r305;
  assign w_000_306 = r306;
  assign w_000_307 = r307;
  assign w_000_308 = r308;
  assign w_000_309 = r309;
  assign w_000_310 = r310;
  assign w_000_311 = r311;
  assign w_000_312 = r312;
  assign w_000_313 = r313;
  assign w_000_314 = r314;
  assign w_000_315 = r315;
  assign w_000_316 = r316;
  assign w_000_317 = r317;
  assign w_000_318 = r318;
  assign w_000_319 = r319;
  assign w_000_320 = r320;
  assign w_000_321 = r321;
  assign w_000_322 = r322;
  assign w_000_323 = r323;
  assign w_000_324 = r324;
  assign w_000_325 = r325;
  assign w_000_326 = r326;
  assign w_000_327 = r327;
  assign w_000_328 = r328;
  assign w_000_329 = r329;
  assign w_000_330 = r330;
  assign w_000_331 = r331;
  assign w_000_332 = r332;
  assign w_000_333 = r333;
  assign w_000_334 = r334;
  assign w_000_335 = r335;
  assign w_000_336 = r336;
  assign w_000_337 = r337;
  assign w_000_338 = r338;
  assign w_000_339 = r339;
  assign w_000_340 = r340;
  assign w_000_341 = r341;
  assign w_000_342 = r342;
  assign w_000_343 = r343;
  assign w_000_344 = r344;
  assign w_000_345 = r345;
  assign w_000_346 = r346;
  assign w_000_347 = r347;
  assign w_000_348 = r348;
  assign w_000_349 = r349;
  assign w_000_350 = r350;
  assign w_000_351 = r351;
  assign w_000_352 = r352;
  assign w_000_353 = r353;
  assign w_000_354 = r354;
  assign w_000_355 = r355;
  assign w_000_356 = r356;
  assign w_000_357 = r357;
  assign w_000_358 = r358;
  assign w_000_359 = r359;
  assign w_000_360 = r360;
  assign w_000_361 = r361;
  assign w_000_362 = r362;
  assign w_000_363 = r363;
  assign w_000_364 = r364;
  assign w_000_365 = r365;
  assign w_000_366 = r366;
  assign w_000_367 = r367;
  assign w_000_368 = r368;
  assign w_000_369 = r369;
  assign w_000_370 = r370;
  assign w_000_371 = r371;
  assign w_000_372 = r372;
  assign w_000_373 = r373;
  assign w_000_374 = r374;
  assign w_000_375 = r375;
  assign w_000_376 = r376;
  assign w_000_377 = r377;
  assign w_000_378 = r378;
  assign w_000_379 = r379;
  assign w_000_380 = r380;
  assign w_000_381 = r381;
  assign w_000_382 = r382;
  assign w_000_383 = r383;
  assign w_000_384 = r384;
  assign w_000_385 = r385;
  assign w_000_386 = r386;
  assign w_000_387 = r387;
  assign w_000_388 = r388;
  assign w_000_389 = r389;
  assign w_000_390 = r390;
  assign w_000_391 = r391;
  assign w_000_392 = r392;
  assign w_000_393 = r393;
  assign w_000_394 = r394;
  assign w_000_395 = r395;
  assign w_000_396 = r396;
  assign w_000_397 = r397;
  assign w_000_398 = r398;
  assign w_000_399 = r399;
  assign w_000_400 = r400;
  assign w_000_401 = r401;
  assign w_000_402 = r402;
  assign w_000_403 = r403;
  assign w_000_404 = r404;
  assign w_000_405 = r405;
  assign w_000_406 = r406;
  assign w_000_407 = r407;
  assign w_000_408 = r408;
  assign w_000_409 = r409;
  assign w_000_410 = r410;
  assign w_000_411 = r411;
  assign w_000_412 = r412;
  assign w_000_413 = r413;
  assign w_000_414 = r414;
  assign w_000_415 = r415;
  assign w_000_416 = r416;
  assign w_000_417 = r417;
  assign w_000_418 = r418;
  assign w_000_419 = r419;
  assign w_000_420 = r420;
  assign w_000_421 = r421;
  assign w_000_422 = r422;
  assign w_000_423 = r423;
  assign w_000_424 = r424;
  assign w_000_425 = r425;
  assign w_000_426 = r426;
  assign w_000_427 = r427;
  assign w_000_428 = r428;
  assign w_000_429 = r429;
  assign w_000_430 = r430;
  assign w_000_431 = r431;
  assign w_000_432 = r432;
  assign w_000_433 = r433;
  assign w_000_434 = r434;
  assign w_000_435 = r435;
  assign w_000_436 = r436;
  assign w_000_437 = r437;
  assign w_000_438 = r438;
  assign w_000_439 = r439;
  assign w_000_440 = r440;
  assign w_000_441 = r441;
  assign w_000_442 = r442;
  assign w_000_443 = r443;
  assign w_000_444 = r444;
  assign w_000_445 = r445;
  assign w_000_446 = r446;
  assign w_000_447 = r447;
  assign w_000_448 = r448;
  assign w_000_449 = r449;
  assign w_000_450 = r450;
  assign w_000_451 = r451;
  assign w_000_452 = r452;
  assign w_000_453 = r453;
  assign w_000_454 = r454;
  assign w_000_455 = r455;
  assign w_000_456 = r456;
  assign w_000_457 = r457;
  assign w_000_458 = r458;
  assign w_000_459 = r459;
  assign w_000_460 = r460;
  assign w_000_461 = r461;
  assign w_000_462 = r462;
  assign w_000_463 = r463;
  assign w_000_464 = r464;
  assign w_000_465 = r465;
  assign w_000_466 = r466;
  assign w_000_467 = r467;
  assign w_000_468 = r468;
  assign w_000_469 = r469;
  assign w_000_470 = r470;
  assign w_000_471 = r471;
  assign w_000_472 = r472;
  assign w_000_473 = r473;
  assign w_000_474 = r474;
  assign w_000_475 = r475;
  assign w_000_476 = r476;
  assign w_000_477 = r477;
  assign w_000_478 = r478;
  assign w_000_479 = r479;
  assign w_000_480 = r480;
  assign w_000_481 = r481;
  assign w_000_482 = r482;
  assign w_000_483 = r483;
  assign w_000_484 = r484;
  assign w_000_485 = r485;
  assign w_000_486 = r486;
  assign w_000_487 = r487;
  assign w_000_488 = r488;
  assign w_000_489 = r489;
  assign w_000_490 = r490;
  assign w_000_491 = r491;
  assign w_000_492 = r492;
  assign w_000_493 = r493;
  assign w_000_494 = r494;
  assign w_000_495 = r495;
  assign w_000_496 = r496;
  assign w_000_497 = r497;
  assign w_000_498 = r498;
  assign w_000_499 = r499;
  assign w_000_500 = r500;
  assign w_000_501 = r501;
  assign w_000_502 = r502;
  assign w_000_503 = r503;
  assign w_000_504 = r504;
  assign w_000_505 = r505;
  assign w_000_506 = r506;
  assign w_000_507 = r507;
  assign w_000_508 = r508;
  assign w_000_509 = r509;
  assign w_000_510 = r510;
  assign w_000_511 = r511;
  assign w_000_512 = r512;
  assign w_000_513 = r513;
  assign w_000_514 = r514;
  assign w_000_515 = r515;
  assign w_000_516 = r516;
  assign w_000_517 = r517;
  assign w_000_518 = r518;
  assign w_000_519 = r519;
  assign w_000_520 = r520;
  assign w_000_521 = r521;
  assign w_000_522 = r522;
  assign w_000_523 = r523;
  assign w_000_524 = r524;
  assign w_000_525 = r525;
  assign w_000_526 = r526;
  assign w_000_527 = r527;
  assign w_000_528 = r528;
  assign w_000_529 = r529;
  assign w_000_530 = r530;
  assign w_000_531 = r531;
  assign w_000_532 = r532;
  assign w_000_533 = r533;
  assign w_000_534 = r534;
  assign w_000_535 = r535;
  assign w_000_536 = r536;
  assign w_000_537 = r537;
  assign w_000_538 = r538;
  assign w_000_539 = r539;
  assign w_000_540 = r540;
  assign w_000_541 = r541;
  assign w_000_542 = r542;
  assign w_000_543 = r543;
  assign w_000_544 = r544;
  assign w_000_545 = r545;
  assign w_000_546 = r546;
  assign w_000_547 = r547;
  assign w_000_548 = r548;
  assign w_000_549 = r549;
  assign w_000_550 = r550;
  assign w_000_551 = r551;
  assign w_000_552 = r552;
  assign w_000_553 = r553;
  assign w_000_554 = r554;
  assign w_000_555 = r555;
  assign w_000_556 = r556;
  assign w_000_557 = r557;
  assign w_000_558 = r558;
  assign w_000_559 = r559;
  assign w_000_560 = r560;
  assign w_000_561 = r561;
  assign w_000_562 = r562;
  assign w_000_563 = r563;
  assign w_000_564 = r564;
  assign w_000_565 = r565;
  assign w_000_566 = r566;
  assign w_000_567 = r567;
  assign w_000_568 = r568;
  assign w_000_569 = r569;
  assign w_000_570 = r570;
  assign w_000_571 = r571;
  assign w_000_572 = r572;
  assign w_000_573 = r573;
  assign w_000_574 = r574;
  assign w_000_575 = r575;
  assign w_000_576 = r576;
  assign w_000_577 = r577;
  assign w_000_578 = r578;
  assign w_000_579 = r579;
  assign w_000_580 = r580;
  assign w_000_581 = r581;
  assign w_000_582 = r582;
  assign w_000_583 = r583;
  assign w_000_584 = r584;
  assign w_000_585 = r585;
  assign w_000_586 = r586;
  assign w_000_587 = r587;
  assign w_000_588 = r588;
  assign w_000_589 = r589;
  assign w_000_590 = r590;
  assign w_000_591 = r591;
  assign w_000_592 = r592;
  assign w_000_593 = r593;
  assign w_000_594 = r594;
  assign w_000_595 = r595;
  assign w_000_596 = r596;
  assign w_000_597 = r597;
  assign w_000_598 = r598;
  assign w_000_599 = r599;
  assign w_000_600 = r600;
  assign w_000_601 = r601;
  assign w_000_602 = r602;
  assign w_000_603 = r603;
  assign w_000_604 = r604;
  assign w_000_605 = r605;
  assign w_000_606 = r606;
  assign w_000_607 = r607;
  assign w_000_608 = r608;
  assign w_000_609 = r609;
  assign w_000_610 = r610;
  assign w_000_611 = r611;
  assign w_000_612 = r612;
  assign w_000_613 = r613;
  assign w_000_614 = r614;
  assign w_000_615 = r615;
  assign w_000_616 = r616;
  assign w_000_617 = r617;
  assign w_000_618 = r618;
  assign w_000_619 = r619;
  assign w_000_620 = r620;
  assign w_000_621 = r621;
  assign w_000_622 = r622;
  assign w_000_623 = r623;
  assign w_000_624 = r624;
  assign w_000_625 = r625;
  assign w_000_626 = r626;
  assign w_000_627 = r627;
  assign w_000_628 = r628;
  assign w_000_629 = r629;
  assign w_000_630 = r630;
  assign w_000_631 = r631;
  assign w_000_632 = r632;
  assign w_000_633 = r633;
  assign w_000_634 = r634;
  assign w_000_635 = r635;
  assign w_000_636 = r636;
  assign w_000_637 = r637;
  assign w_000_638 = r638;
  assign w_000_639 = r639;
  assign w_000_640 = r640;
  assign w_000_641 = r641;
  assign w_000_642 = r642;
  assign w_000_643 = r643;
  assign w_000_644 = r644;
  assign w_000_645 = r645;
  assign w_000_646 = r646;
  assign w_000_647 = r647;
  assign w_000_648 = r648;
  assign w_000_649 = r649;
  assign w_000_650 = r650;
  assign w_000_651 = r651;
  assign w_000_652 = r652;
  assign w_000_653 = r653;
  assign w_000_654 = r654;
  assign w_000_655 = r655;
  assign w_000_656 = r656;
  assign w_000_657 = r657;
  assign w_000_658 = r658;
  assign w_000_659 = r659;
  assign w_000_660 = r660;
  assign w_000_661 = r661;
  assign w_000_662 = r662;
  assign w_000_663 = r663;
  assign w_000_664 = r664;
  assign w_000_665 = r665;
  assign w_000_666 = r666;
  assign w_000_667 = r667;
  assign w_000_668 = r668;
  assign w_000_669 = r669;
  assign w_000_670 = r670;
  assign w_000_671 = r671;
  assign w_000_672 = r672;
  assign w_000_673 = r673;
  assign w_000_674 = r674;
  assign w_000_675 = r675;
  assign w_000_676 = r676;
  assign w_000_677 = r677;
  assign w_000_678 = r678;
  assign w_000_679 = r679;
  assign w_000_680 = r680;
  assign w_000_681 = r681;
  assign w_000_682 = r682;
  assign w_000_683 = r683;
  assign w_000_684 = r684;
  assign w_000_685 = r685;
  assign w_000_686 = r686;
  assign w_000_687 = r687;
  assign w_000_688 = r688;
  assign w_000_689 = r689;
  assign w_000_690 = r690;
  assign w_000_691 = r691;
  assign w_000_692 = r692;
  assign w_000_693 = r693;
  assign w_000_694 = r694;
  assign w_000_695 = r695;
  assign w_000_696 = r696;
  assign w_000_697 = r697;
  assign w_000_698 = r698;
  assign w_000_699 = r699;
  assign w_000_700 = r700;
  assign w_000_701 = r701;
  assign w_000_702 = r702;
  assign w_000_703 = r703;
  assign w_000_704 = r704;
  assign w_000_705 = r705;
  assign w_000_706 = r706;
  assign w_000_707 = r707;
  assign w_000_708 = r708;
  assign w_000_709 = r709;
  assign w_000_710 = r710;
  assign w_000_711 = r711;
  assign w_000_712 = r712;
  assign w_000_713 = r713;
  assign w_000_714 = r714;
  assign w_000_715 = r715;
  assign w_000_716 = r716;
  assign w_000_717 = r717;
  assign w_000_718 = r718;
  assign w_000_719 = r719;
  assign w_000_720 = r720;
  assign w_000_721 = r721;
  assign w_000_722 = r722;
  assign w_000_723 = r723;
  assign w_000_724 = r724;
  assign w_000_725 = r725;
  assign w_000_726 = r726;
  assign w_000_727 = r727;
  assign w_000_728 = r728;
  assign w_000_729 = r729;
  assign w_000_730 = r730;
  assign w_000_731 = r731;
  assign w_000_732 = r732;
  assign w_000_733 = r733;
  assign w_000_734 = r734;
  assign w_000_735 = r735;
  assign w_000_736 = r736;
  assign w_000_737 = r737;
  assign w_000_738 = r738;
  assign w_000_739 = r739;
  assign w_000_740 = r740;
  assign w_000_741 = r741;
  assign w_000_742 = r742;
  assign w_000_743 = r743;
  assign w_000_744 = r744;
  assign w_000_745 = r745;
  assign w_000_746 = r746;
  assign w_000_747 = r747;
  assign w_000_748 = r748;
  assign w_000_749 = r749;
  assign w_000_750 = r750;
  assign w_000_751 = r751;
  assign w_000_752 = r752;
  assign w_000_753 = r753;
  assign w_000_754 = r754;
  assign w_000_755 = r755;
  assign w_000_756 = r756;
  assign w_000_757 = r757;
  assign w_000_758 = r758;
  assign w_000_759 = r759;
  assign w_000_760 = r760;
  assign w_000_761 = r761;
  assign w_000_762 = r762;
  assign w_000_763 = r763;
  assign w_000_764 = r764;
  assign w_000_765 = r765;
  assign w_000_766 = r766;
  assign w_000_767 = r767;
  assign w_000_768 = r768;
  assign w_000_769 = r769;
  assign w_000_770 = r770;
  assign w_000_771 = r771;
  assign w_000_772 = r772;
  assign w_000_773 = r773;
  assign w_000_774 = r774;
  assign w_000_775 = r775;
  assign w_000_776 = r776;
  assign w_000_777 = r777;
  assign w_000_778 = r778;
  assign w_000_779 = r779;
  assign w_000_780 = r780;
  assign w_000_781 = r781;
  assign w_000_782 = r782;
  assign w_000_783 = r783;
  assign w_000_784 = r784;
  assign w_000_785 = r785;
  assign w_000_786 = r786;
  assign w_000_787 = r787;
  assign w_000_788 = r788;
  assign w_000_789 = r789;
  assign w_000_790 = r790;
  assign w_000_791 = r791;
  assign w_000_792 = r792;
  assign w_000_793 = r793;
  assign w_000_794 = r794;
  assign w_000_795 = r795;
  assign w_000_796 = r796;
  assign w_000_797 = r797;
  assign w_000_798 = r798;
  assign w_000_799 = r799;
  assign w_000_800 = r800;
  assign w_000_801 = r801;
  assign w_000_802 = r802;
  assign w_000_803 = r803;
  assign w_000_804 = r804;
  assign w_000_805 = r805;
  assign w_000_806 = r806;
  assign w_000_807 = r807;
  assign w_000_808 = r808;
  assign w_000_809 = r809;
  assign w_000_810 = r810;
  assign w_000_811 = r811;
  assign w_000_812 = r812;
  assign w_000_813 = r813;
  assign w_000_814 = r814;
  assign w_000_815 = r815;
  assign w_000_816 = r816;
  assign w_000_817 = r817;
  assign w_000_818 = r818;
  assign w_000_819 = r819;
  assign w_000_820 = r820;
  assign w_000_821 = r821;
  assign w_000_822 = r822;
  assign w_000_823 = r823;
  assign w_000_824 = r824;
  assign w_000_825 = r825;
  assign w_000_826 = r826;
  assign w_000_827 = r827;
  assign w_000_828 = r828;
  assign w_000_829 = r829;
  assign w_000_830 = r830;
  assign w_000_831 = r831;
  assign w_000_832 = r832;
  assign w_000_833 = r833;
  assign w_000_834 = r834;
  assign w_000_835 = r835;
  assign w_000_836 = r836;
  assign w_000_837 = r837;
  assign w_000_838 = r838;
  assign w_000_839 = r839;
  assign w_000_840 = r840;
  assign w_000_841 = r841;
  assign w_000_842 = r842;
  assign w_000_843 = r843;
  assign w_000_844 = r844;
  assign w_000_845 = r845;
  assign w_000_846 = r846;
  assign w_000_847 = r847;
  assign w_000_848 = r848;
  assign w_000_849 = r849;
  assign w_000_850 = r850;
  assign w_000_851 = r851;
  assign w_000_852 = r852;
  assign w_000_853 = r853;
  assign w_000_854 = r854;
  assign w_000_855 = r855;
  assign w_000_856 = r856;
  assign w_000_857 = r857;
  assign w_000_858 = r858;
  assign w_000_859 = r859;
  assign w_000_860 = r860;
  assign w_000_861 = r861;
  assign w_000_862 = r862;
  assign w_000_863 = r863;
  assign w_000_864 = r864;
  assign w_000_865 = r865;
  assign w_000_866 = r866;
  assign w_000_867 = r867;
  assign w_000_868 = r868;
  assign w_000_869 = r869;
  assign w_000_870 = r870;
  assign w_000_871 = r871;
  assign w_000_872 = r872;
  assign w_000_873 = r873;
  assign w_000_874 = r874;
  assign w_000_875 = r875;
  assign w_000_876 = r876;
  assign w_000_877 = r877;
  assign w_000_878 = r878;
  assign w_000_879 = r879;
  assign w_000_880 = r880;
  assign w_000_881 = r881;
  assign w_000_882 = r882;
  assign w_000_883 = r883;
  assign w_000_884 = r884;
  assign w_000_885 = r885;
  assign w_000_886 = r886;
  assign w_000_887 = r887;
  assign w_000_888 = r888;
  assign w_000_889 = r889;
  assign w_000_890 = r890;
  assign w_000_891 = r891;
  assign w_000_892 = r892;
  assign w_000_893 = r893;
  assign w_000_894 = r894;
  assign w_000_895 = r895;
  assign w_000_896 = r896;
  assign w_000_897 = r897;
  assign w_000_898 = r898;
  assign w_000_899 = r899;
  assign w_000_900 = r900;
  assign w_000_901 = r901;
  assign w_000_902 = r902;
  assign w_000_903 = r903;
  assign w_000_904 = r904;
  assign w_000_905 = r905;
  assign w_000_906 = r906;
  assign w_000_907 = r907;
  assign w_000_908 = r908;
  assign w_000_909 = r909;
  assign w_000_910 = r910;
  assign w_000_911 = r911;
  assign w_000_912 = r912;
  assign w_000_913 = r913;
  assign w_000_914 = r914;
  assign w_000_915 = r915;
  assign w_000_916 = r916;
  assign w_000_917 = r917;
  assign w_000_918 = r918;
  assign w_000_919 = r919;
  assign w_000_920 = r920;
  assign w_000_921 = r921;
  assign w_000_922 = r922;
  assign w_000_923 = r923;
  assign w_000_924 = r924;
  assign w_000_925 = r925;
  assign w_000_926 = r926;
  assign w_000_927 = r927;
  assign w_000_928 = r928;
  assign w_000_929 = r929;
  assign w_000_930 = r930;
  assign w_000_931 = r931;
  assign w_000_932 = r932;
  assign w_000_933 = r933;
  assign w_000_934 = r934;
  assign w_000_935 = r935;
  assign w_000_936 = r936;
  assign w_000_937 = r937;
  assign w_000_938 = r938;
  assign w_000_939 = r939;
  assign w_000_940 = r940;
  assign w_000_941 = r941;
  assign w_000_942 = r942;
  assign w_000_943 = r943;
  assign w_000_944 = r944;
  assign w_000_945 = r945;
  assign w_000_946 = r946;
  assign w_000_947 = r947;
  assign w_000_948 = r948;
  assign w_000_949 = r949;
  assign w_000_950 = r950;
  assign w_000_951 = r951;
  assign w_000_952 = r952;
  assign w_000_953 = r953;
  assign w_000_954 = r954;
  assign w_000_955 = r955;
  assign w_000_956 = r956;
  assign w_000_957 = r957;
  assign w_000_958 = r958;
  assign w_000_959 = r959;
  assign w_000_960 = r960;
  assign w_000_961 = r961;
  assign w_000_962 = r962;
  assign w_000_963 = r963;
  assign w_000_964 = r964;
  assign w_000_965 = r965;
  assign w_000_966 = r966;
  assign w_000_967 = r967;
  assign w_000_968 = r968;
  assign w_000_969 = r969;
  assign w_000_970 = r970;
  assign w_000_971 = r971;
  assign w_000_972 = r972;
  assign w_000_973 = r973;
  assign w_000_974 = r974;
  assign w_000_975 = r975;
  assign w_000_976 = r976;
  assign w_000_977 = r977;
  assign w_000_978 = r978;
  assign w_000_979 = r979;
  assign w_000_980 = r980;
  assign w_000_981 = r981;
  assign w_000_982 = r982;
  assign w_000_983 = r983;
  assign w_000_984 = r984;
  assign w_000_985 = r985;
  assign w_000_986 = r986;
  assign w_000_987 = r987;
  assign w_000_988 = r988;
  assign w_000_989 = r989;
  assign w_000_990 = r990;
  assign w_000_991 = r991;
  assign w_000_992 = r992;
  assign w_000_993 = r993;
  assign w_000_994 = r994;
  assign w_000_995 = r995;
  assign w_000_996 = r996;
  assign w_000_997 = r997;
  assign w_000_998 = r998;
  assign w_000_999 = r999;

  initial begin 
    r0 = 1'b0; 
    r1 = 1'b0; 
    r2 = 1'b0; 
    r3 = 1'b0; 
    r4 = 1'b0; 
    r5 = 1'b0; 
    r6 = 1'b0; 
    r7 = 1'b0; 
    r8 = 1'b0; 
    r9 = 1'b0; 
    r10 = 1'b0; 
    r11 = 1'b0; 
    r12 = 1'b0; 
    r13 = 1'b0; 
    r14 = 1'b0; 
    r15 = 1'b0; 
    r16 = 1'b0; 
    r17 = 1'b0; 
    r18 = 1'b0; 
    r19 = 1'b0; 
    r20 = 1'b0; 
    r21 = 1'b0; 
    r22 = 1'b0; 
    r23 = 1'b0; 
    r24 = 1'b0; 
    r25 = 1'b0; 
    r26 = 1'b0; 
    r27 = 1'b0; 
    r28 = 1'b0; 
    r29 = 1'b0; 
    r30 = 1'b0; 
    r31 = 1'b0; 
    r32 = 1'b0; 
    r33 = 1'b0; 
    r34 = 1'b0; 
    r35 = 1'b0; 
    r36 = 1'b0; 
    r37 = 1'b0; 
    r38 = 1'b0; 
    r39 = 1'b0; 
    r40 = 1'b0; 
    r41 = 1'b0; 
    r42 = 1'b0; 
    r43 = 1'b0; 
    r44 = 1'b0; 
    r45 = 1'b0; 
    r46 = 1'b0; 
    r47 = 1'b0; 
    r48 = 1'b0; 
    r49 = 1'b0; 
    r50 = 1'b0; 
    r51 = 1'b0; 
    r52 = 1'b0; 
    r53 = 1'b0; 
    r54 = 1'b0; 
    r55 = 1'b0; 
    r56 = 1'b0; 
    r57 = 1'b0; 
    r58 = 1'b0; 
    r59 = 1'b0; 
    r60 = 1'b0; 
    r61 = 1'b0; 
    r62 = 1'b0; 
    r63 = 1'b0; 
    r64 = 1'b0; 
    r65 = 1'b0; 
    r66 = 1'b0; 
    r67 = 1'b0; 
    r68 = 1'b0; 
    r69 = 1'b0; 
    r70 = 1'b0; 
    r71 = 1'b0; 
    r72 = 1'b0; 
    r73 = 1'b0; 
    r74 = 1'b0; 
    r75 = 1'b0; 
    r76 = 1'b0; 
    r77 = 1'b0; 
    r78 = 1'b0; 
    r79 = 1'b0; 
    r80 = 1'b0; 
    r81 = 1'b0; 
    r82 = 1'b0; 
    r83 = 1'b0; 
    r84 = 1'b0; 
    r85 = 1'b0; 
    r86 = 1'b0; 
    r87 = 1'b0; 
    r88 = 1'b0; 
    r89 = 1'b0; 
    r90 = 1'b0; 
    r91 = 1'b0; 
    r92 = 1'b0; 
    r93 = 1'b0; 
    r94 = 1'b0; 
    r95 = 1'b0; 
    r96 = 1'b0; 
    r97 = 1'b0; 
    r98 = 1'b0; 
    r99 = 1'b0; 
    r100 = 1'b0; 
    r101 = 1'b0; 
    r102 = 1'b0; 
    r103 = 1'b0; 
    r104 = 1'b0; 
    r105 = 1'b0; 
    r106 = 1'b0; 
    r107 = 1'b0; 
    r108 = 1'b0; 
    r109 = 1'b0; 
    r110 = 1'b0; 
    r111 = 1'b0; 
    r112 = 1'b0; 
    r113 = 1'b0; 
    r114 = 1'b0; 
    r115 = 1'b0; 
    r116 = 1'b0; 
    r117 = 1'b0; 
    r118 = 1'b0; 
    r119 = 1'b0; 
    r120 = 1'b0; 
    r121 = 1'b0; 
    r122 = 1'b0; 
    r123 = 1'b0; 
    r124 = 1'b0; 
    r125 = 1'b0; 
    r126 = 1'b0; 
    r127 = 1'b0; 
    r128 = 1'b0; 
    r129 = 1'b0; 
    r130 = 1'b0; 
    r131 = 1'b0; 
    r132 = 1'b0; 
    r133 = 1'b0; 
    r134 = 1'b0; 
    r135 = 1'b0; 
    r136 = 1'b0; 
    r137 = 1'b0; 
    r138 = 1'b0; 
    r139 = 1'b0; 
    r140 = 1'b0; 
    r141 = 1'b0; 
    r142 = 1'b0; 
    r143 = 1'b0; 
    r144 = 1'b0; 
    r145 = 1'b0; 
    r146 = 1'b0; 
    r147 = 1'b0; 
    r148 = 1'b0; 
    r149 = 1'b0; 
    r150 = 1'b0; 
    r151 = 1'b0; 
    r152 = 1'b0; 
    r153 = 1'b0; 
    r154 = 1'b0; 
    r155 = 1'b0; 
    r156 = 1'b0; 
    r157 = 1'b0; 
    r158 = 1'b0; 
    r159 = 1'b0; 
    r160 = 1'b0; 
    r161 = 1'b0; 
    r162 = 1'b0; 
    r163 = 1'b0; 
    r164 = 1'b0; 
    r165 = 1'b0; 
    r166 = 1'b0; 
    r167 = 1'b0; 
    r168 = 1'b0; 
    r169 = 1'b0; 
    r170 = 1'b0; 
    r171 = 1'b0; 
    r172 = 1'b0; 
    r173 = 1'b0; 
    r174 = 1'b0; 
    r175 = 1'b0; 
    r176 = 1'b0; 
    r177 = 1'b0; 
    r178 = 1'b0; 
    r179 = 1'b0; 
    r180 = 1'b0; 
    r181 = 1'b0; 
    r182 = 1'b0; 
    r183 = 1'b0; 
    r184 = 1'b0; 
    r185 = 1'b0; 
    r186 = 1'b0; 
    r187 = 1'b0; 
    r188 = 1'b0; 
    r189 = 1'b0; 
    r190 = 1'b0; 
    r191 = 1'b0; 
    r192 = 1'b0; 
    r193 = 1'b0; 
    r194 = 1'b0; 
    r195 = 1'b0; 
    r196 = 1'b0; 
    r197 = 1'b0; 
    r198 = 1'b0; 
    r199 = 1'b0; 
    r200 = 1'b0; 
    r201 = 1'b0; 
    r202 = 1'b0; 
    r203 = 1'b0; 
    r204 = 1'b0; 
    r205 = 1'b0; 
    r206 = 1'b0; 
    r207 = 1'b0; 
    r208 = 1'b0; 
    r209 = 1'b0; 
    r210 = 1'b0; 
    r211 = 1'b0; 
    r212 = 1'b0; 
    r213 = 1'b0; 
    r214 = 1'b0; 
    r215 = 1'b0; 
    r216 = 1'b0; 
    r217 = 1'b0; 
    r218 = 1'b0; 
    r219 = 1'b0; 
    r220 = 1'b0; 
    r221 = 1'b0; 
    r222 = 1'b0; 
    r223 = 1'b0; 
    r224 = 1'b0; 
    r225 = 1'b0; 
    r226 = 1'b0; 
    r227 = 1'b0; 
    r228 = 1'b0; 
    r229 = 1'b0; 
    r230 = 1'b0; 
    r231 = 1'b0; 
    r232 = 1'b0; 
    r233 = 1'b0; 
    r234 = 1'b0; 
    r235 = 1'b0; 
    r236 = 1'b0; 
    r237 = 1'b0; 
    r238 = 1'b0; 
    r239 = 1'b0; 
    r240 = 1'b0; 
    r241 = 1'b0; 
    r242 = 1'b0; 
    r243 = 1'b0; 
    r244 = 1'b0; 
    r245 = 1'b0; 
    r246 = 1'b0; 
    r247 = 1'b0; 
    r248 = 1'b0; 
    r249 = 1'b0; 
    r250 = 1'b0; 
    r251 = 1'b0; 
    r252 = 1'b0; 
    r253 = 1'b0; 
    r254 = 1'b0; 
    r255 = 1'b0; 
    r256 = 1'b0; 
    r257 = 1'b0; 
    r258 = 1'b0; 
    r259 = 1'b0; 
    r260 = 1'b0; 
    r261 = 1'b0; 
    r262 = 1'b0; 
    r263 = 1'b0; 
    r264 = 1'b0; 
    r265 = 1'b0; 
    r266 = 1'b0; 
    r267 = 1'b0; 
    r268 = 1'b0; 
    r269 = 1'b0; 
    r270 = 1'b0; 
    r271 = 1'b0; 
    r272 = 1'b0; 
    r273 = 1'b0; 
    r274 = 1'b0; 
    r275 = 1'b0; 
    r276 = 1'b0; 
    r277 = 1'b0; 
    r278 = 1'b0; 
    r279 = 1'b0; 
    r280 = 1'b0; 
    r281 = 1'b0; 
    r282 = 1'b0; 
    r283 = 1'b0; 
    r284 = 1'b0; 
    r285 = 1'b0; 
    r286 = 1'b0; 
    r287 = 1'b0; 
    r288 = 1'b0; 
    r289 = 1'b0; 
    r290 = 1'b0; 
    r291 = 1'b0; 
    r292 = 1'b0; 
    r293 = 1'b0; 
    r294 = 1'b0; 
    r295 = 1'b0; 
    r296 = 1'b0; 
    r297 = 1'b0; 
    r298 = 1'b0; 
    r299 = 1'b0; 
    r300 = 1'b0; 
    r301 = 1'b0; 
    r302 = 1'b0; 
    r303 = 1'b0; 
    r304 = 1'b0; 
    r305 = 1'b0; 
    r306 = 1'b0; 
    r307 = 1'b0; 
    r308 = 1'b0; 
    r309 = 1'b0; 
    r310 = 1'b0; 
    r311 = 1'b0; 
    r312 = 1'b0; 
    r313 = 1'b0; 
    r314 = 1'b0; 
    r315 = 1'b0; 
    r316 = 1'b0; 
    r317 = 1'b0; 
    r318 = 1'b0; 
    r319 = 1'b0; 
    r320 = 1'b0; 
    r321 = 1'b0; 
    r322 = 1'b0; 
    r323 = 1'b0; 
    r324 = 1'b0; 
    r325 = 1'b0; 
    r326 = 1'b0; 
    r327 = 1'b0; 
    r328 = 1'b0; 
    r329 = 1'b0; 
    r330 = 1'b0; 
    r331 = 1'b0; 
    r332 = 1'b0; 
    r333 = 1'b0; 
    r334 = 1'b0; 
    r335 = 1'b0; 
    r336 = 1'b0; 
    r337 = 1'b0; 
    r338 = 1'b0; 
    r339 = 1'b0; 
    r340 = 1'b0; 
    r341 = 1'b0; 
    r342 = 1'b0; 
    r343 = 1'b0; 
    r344 = 1'b0; 
    r345 = 1'b0; 
    r346 = 1'b0; 
    r347 = 1'b0; 
    r348 = 1'b0; 
    r349 = 1'b0; 
    r350 = 1'b0; 
    r351 = 1'b0; 
    r352 = 1'b0; 
    r353 = 1'b0; 
    r354 = 1'b0; 
    r355 = 1'b0; 
    r356 = 1'b0; 
    r357 = 1'b0; 
    r358 = 1'b0; 
    r359 = 1'b0; 
    r360 = 1'b0; 
    r361 = 1'b0; 
    r362 = 1'b0; 
    r363 = 1'b0; 
    r364 = 1'b0; 
    r365 = 1'b0; 
    r366 = 1'b0; 
    r367 = 1'b0; 
    r368 = 1'b0; 
    r369 = 1'b0; 
    r370 = 1'b0; 
    r371 = 1'b0; 
    r372 = 1'b0; 
    r373 = 1'b0; 
    r374 = 1'b0; 
    r375 = 1'b0; 
    r376 = 1'b0; 
    r377 = 1'b0; 
    r378 = 1'b0; 
    r379 = 1'b0; 
    r380 = 1'b0; 
    r381 = 1'b0; 
    r382 = 1'b0; 
    r383 = 1'b0; 
    r384 = 1'b0; 
    r385 = 1'b0; 
    r386 = 1'b0; 
    r387 = 1'b0; 
    r388 = 1'b0; 
    r389 = 1'b0; 
    r390 = 1'b0; 
    r391 = 1'b0; 
    r392 = 1'b0; 
    r393 = 1'b0; 
    r394 = 1'b0; 
    r395 = 1'b0; 
    r396 = 1'b0; 
    r397 = 1'b0; 
    r398 = 1'b0; 
    r399 = 1'b0; 
    r400 = 1'b0; 
    r401 = 1'b0; 
    r402 = 1'b0; 
    r403 = 1'b0; 
    r404 = 1'b0; 
    r405 = 1'b0; 
    r406 = 1'b0; 
    r407 = 1'b0; 
    r408 = 1'b0; 
    r409 = 1'b0; 
    r410 = 1'b0; 
    r411 = 1'b0; 
    r412 = 1'b0; 
    r413 = 1'b0; 
    r414 = 1'b0; 
    r415 = 1'b0; 
    r416 = 1'b0; 
    r417 = 1'b0; 
    r418 = 1'b0; 
    r419 = 1'b0; 
    r420 = 1'b0; 
    r421 = 1'b0; 
    r422 = 1'b0; 
    r423 = 1'b0; 
    r424 = 1'b0; 
    r425 = 1'b0; 
    r426 = 1'b0; 
    r427 = 1'b0; 
    r428 = 1'b0; 
    r429 = 1'b0; 
    r430 = 1'b0; 
    r431 = 1'b0; 
    r432 = 1'b0; 
    r433 = 1'b0; 
    r434 = 1'b0; 
    r435 = 1'b0; 
    r436 = 1'b0; 
    r437 = 1'b0; 
    r438 = 1'b0; 
    r439 = 1'b0; 
    r440 = 1'b0; 
    r441 = 1'b0; 
    r442 = 1'b0; 
    r443 = 1'b0; 
    r444 = 1'b0; 
    r445 = 1'b0; 
    r446 = 1'b0; 
    r447 = 1'b0; 
    r448 = 1'b0; 
    r449 = 1'b0; 
    r450 = 1'b0; 
    r451 = 1'b0; 
    r452 = 1'b0; 
    r453 = 1'b0; 
    r454 = 1'b0; 
    r455 = 1'b0; 
    r456 = 1'b0; 
    r457 = 1'b0; 
    r458 = 1'b0; 
    r459 = 1'b0; 
    r460 = 1'b0; 
    r461 = 1'b0; 
    r462 = 1'b0; 
    r463 = 1'b0; 
    r464 = 1'b0; 
    r465 = 1'b0; 
    r466 = 1'b0; 
    r467 = 1'b0; 
    r468 = 1'b0; 
    r469 = 1'b0; 
    r470 = 1'b0; 
    r471 = 1'b0; 
    r472 = 1'b0; 
    r473 = 1'b0; 
    r474 = 1'b0; 
    r475 = 1'b0; 
    r476 = 1'b0; 
    r477 = 1'b0; 
    r478 = 1'b0; 
    r479 = 1'b0; 
    r480 = 1'b0; 
    r481 = 1'b0; 
    r482 = 1'b0; 
    r483 = 1'b0; 
    r484 = 1'b0; 
    r485 = 1'b0; 
    r486 = 1'b0; 
    r487 = 1'b0; 
    r488 = 1'b0; 
    r489 = 1'b0; 
    r490 = 1'b0; 
    r491 = 1'b0; 
    r492 = 1'b0; 
    r493 = 1'b0; 
    r494 = 1'b0; 
    r495 = 1'b0; 
    r496 = 1'b0; 
    r497 = 1'b0; 
    r498 = 1'b0; 
    r499 = 1'b0; 
    r500 = 1'b0; 
    r501 = 1'b0; 
    r502 = 1'b0; 
    r503 = 1'b0; 
    r504 = 1'b0; 
    r505 = 1'b0; 
    r506 = 1'b0; 
    r507 = 1'b0; 
    r508 = 1'b0; 
    r509 = 1'b0; 
    r510 = 1'b0; 
    r511 = 1'b0; 
    r512 = 1'b0; 
    r513 = 1'b0; 
    r514 = 1'b0; 
    r515 = 1'b0; 
    r516 = 1'b0; 
    r517 = 1'b0; 
    r518 = 1'b0; 
    r519 = 1'b0; 
    r520 = 1'b0; 
    r521 = 1'b0; 
    r522 = 1'b0; 
    r523 = 1'b0; 
    r524 = 1'b0; 
    r525 = 1'b0; 
    r526 = 1'b0; 
    r527 = 1'b0; 
    r528 = 1'b0; 
    r529 = 1'b0; 
    r530 = 1'b0; 
    r531 = 1'b0; 
    r532 = 1'b0; 
    r533 = 1'b0; 
    r534 = 1'b0; 
    r535 = 1'b0; 
    r536 = 1'b0; 
    r537 = 1'b0; 
    r538 = 1'b0; 
    r539 = 1'b0; 
    r540 = 1'b0; 
    r541 = 1'b0; 
    r542 = 1'b0; 
    r543 = 1'b0; 
    r544 = 1'b0; 
    r545 = 1'b0; 
    r546 = 1'b0; 
    r547 = 1'b0; 
    r548 = 1'b0; 
    r549 = 1'b0; 
    r550 = 1'b0; 
    r551 = 1'b0; 
    r552 = 1'b0; 
    r553 = 1'b0; 
    r554 = 1'b0; 
    r555 = 1'b0; 
    r556 = 1'b0; 
    r557 = 1'b0; 
    r558 = 1'b0; 
    r559 = 1'b0; 
    r560 = 1'b0; 
    r561 = 1'b0; 
    r562 = 1'b0; 
    r563 = 1'b0; 
    r564 = 1'b0; 
    r565 = 1'b0; 
    r566 = 1'b0; 
    r567 = 1'b0; 
    r568 = 1'b0; 
    r569 = 1'b0; 
    r570 = 1'b0; 
    r571 = 1'b0; 
    r572 = 1'b0; 
    r573 = 1'b0; 
    r574 = 1'b0; 
    r575 = 1'b0; 
    r576 = 1'b0; 
    r577 = 1'b0; 
    r578 = 1'b0; 
    r579 = 1'b0; 
    r580 = 1'b0; 
    r581 = 1'b0; 
    r582 = 1'b0; 
    r583 = 1'b0; 
    r584 = 1'b0; 
    r585 = 1'b0; 
    r586 = 1'b0; 
    r587 = 1'b0; 
    r588 = 1'b0; 
    r589 = 1'b0; 
    r590 = 1'b0; 
    r591 = 1'b0; 
    r592 = 1'b0; 
    r593 = 1'b0; 
    r594 = 1'b0; 
    r595 = 1'b0; 
    r596 = 1'b0; 
    r597 = 1'b0; 
    r598 = 1'b0; 
    r599 = 1'b0; 
    r600 = 1'b0; 
    r601 = 1'b0; 
    r602 = 1'b0; 
    r603 = 1'b0; 
    r604 = 1'b0; 
    r605 = 1'b0; 
    r606 = 1'b0; 
    r607 = 1'b0; 
    r608 = 1'b0; 
    r609 = 1'b0; 
    r610 = 1'b0; 
    r611 = 1'b0; 
    r612 = 1'b0; 
    r613 = 1'b0; 
    r614 = 1'b0; 
    r615 = 1'b0; 
    r616 = 1'b0; 
    r617 = 1'b0; 
    r618 = 1'b0; 
    r619 = 1'b0; 
    r620 = 1'b0; 
    r621 = 1'b0; 
    r622 = 1'b0; 
    r623 = 1'b0; 
    r624 = 1'b0; 
    r625 = 1'b0; 
    r626 = 1'b0; 
    r627 = 1'b0; 
    r628 = 1'b0; 
    r629 = 1'b0; 
    r630 = 1'b0; 
    r631 = 1'b0; 
    r632 = 1'b0; 
    r633 = 1'b0; 
    r634 = 1'b0; 
    r635 = 1'b0; 
    r636 = 1'b0; 
    r637 = 1'b0; 
    r638 = 1'b0; 
    r639 = 1'b0; 
    r640 = 1'b0; 
    r641 = 1'b0; 
    r642 = 1'b0; 
    r643 = 1'b0; 
    r644 = 1'b0; 
    r645 = 1'b0; 
    r646 = 1'b0; 
    r647 = 1'b0; 
    r648 = 1'b0; 
    r649 = 1'b0; 
    r650 = 1'b0; 
    r651 = 1'b0; 
    r652 = 1'b0; 
    r653 = 1'b0; 
    r654 = 1'b0; 
    r655 = 1'b0; 
    r656 = 1'b0; 
    r657 = 1'b0; 
    r658 = 1'b0; 
    r659 = 1'b0; 
    r660 = 1'b0; 
    r661 = 1'b0; 
    r662 = 1'b0; 
    r663 = 1'b0; 
    r664 = 1'b0; 
    r665 = 1'b0; 
    r666 = 1'b0; 
    r667 = 1'b0; 
    r668 = 1'b0; 
    r669 = 1'b0; 
    r670 = 1'b0; 
    r671 = 1'b0; 
    r672 = 1'b0; 
    r673 = 1'b0; 
    r674 = 1'b0; 
    r675 = 1'b0; 
    r676 = 1'b0; 
    r677 = 1'b0; 
    r678 = 1'b0; 
    r679 = 1'b0; 
    r680 = 1'b0; 
    r681 = 1'b0; 
    r682 = 1'b0; 
    r683 = 1'b0; 
    r684 = 1'b0; 
    r685 = 1'b0; 
    r686 = 1'b0; 
    r687 = 1'b0; 
    r688 = 1'b0; 
    r689 = 1'b0; 
    r690 = 1'b0; 
    r691 = 1'b0; 
    r692 = 1'b0; 
    r693 = 1'b0; 
    r694 = 1'b0; 
    r695 = 1'b0; 
    r696 = 1'b0; 
    r697 = 1'b0; 
    r698 = 1'b0; 
    r699 = 1'b0; 
    r700 = 1'b0; 
    r701 = 1'b0; 
    r702 = 1'b0; 
    r703 = 1'b0; 
    r704 = 1'b0; 
    r705 = 1'b0; 
    r706 = 1'b0; 
    r707 = 1'b0; 
    r708 = 1'b0; 
    r709 = 1'b0; 
    r710 = 1'b0; 
    r711 = 1'b0; 
    r712 = 1'b0; 
    r713 = 1'b0; 
    r714 = 1'b0; 
    r715 = 1'b0; 
    r716 = 1'b0; 
    r717 = 1'b0; 
    r718 = 1'b0; 
    r719 = 1'b0; 
    r720 = 1'b0; 
    r721 = 1'b0; 
    r722 = 1'b0; 
    r723 = 1'b0; 
    r724 = 1'b0; 
    r725 = 1'b0; 
    r726 = 1'b0; 
    r727 = 1'b0; 
    r728 = 1'b0; 
    r729 = 1'b0; 
    r730 = 1'b0; 
    r731 = 1'b0; 
    r732 = 1'b0; 
    r733 = 1'b0; 
    r734 = 1'b0; 
    r735 = 1'b0; 
    r736 = 1'b0; 
    r737 = 1'b0; 
    r738 = 1'b0; 
    r739 = 1'b0; 
    r740 = 1'b0; 
    r741 = 1'b0; 
    r742 = 1'b0; 
    r743 = 1'b0; 
    r744 = 1'b0; 
    r745 = 1'b0; 
    r746 = 1'b0; 
    r747 = 1'b0; 
    r748 = 1'b0; 
    r749 = 1'b0; 
    r750 = 1'b0; 
    r751 = 1'b0; 
    r752 = 1'b0; 
    r753 = 1'b0; 
    r754 = 1'b0; 
    r755 = 1'b0; 
    r756 = 1'b0; 
    r757 = 1'b0; 
    r758 = 1'b0; 
    r759 = 1'b0; 
    r760 = 1'b0; 
    r761 = 1'b0; 
    r762 = 1'b0; 
    r763 = 1'b0; 
    r764 = 1'b0; 
    r765 = 1'b0; 
    r766 = 1'b0; 
    r767 = 1'b0; 
    r768 = 1'b0; 
    r769 = 1'b0; 
    r770 = 1'b0; 
    r771 = 1'b0; 
    r772 = 1'b0; 
    r773 = 1'b0; 
    r774 = 1'b0; 
    r775 = 1'b0; 
    r776 = 1'b0; 
    r777 = 1'b0; 
    r778 = 1'b0; 
    r779 = 1'b0; 
    r780 = 1'b0; 
    r781 = 1'b0; 
    r782 = 1'b0; 
    r783 = 1'b0; 
    r784 = 1'b0; 
    r785 = 1'b0; 
    r786 = 1'b0; 
    r787 = 1'b0; 
    r788 = 1'b0; 
    r789 = 1'b0; 
    r790 = 1'b0; 
    r791 = 1'b0; 
    r792 = 1'b0; 
    r793 = 1'b0; 
    r794 = 1'b0; 
    r795 = 1'b0; 
    r796 = 1'b0; 
    r797 = 1'b0; 
    r798 = 1'b0; 
    r799 = 1'b0; 
    r800 = 1'b0; 
    r801 = 1'b0; 
    r802 = 1'b0; 
    r803 = 1'b0; 
    r804 = 1'b0; 
    r805 = 1'b0; 
    r806 = 1'b0; 
    r807 = 1'b0; 
    r808 = 1'b0; 
    r809 = 1'b0; 
    r810 = 1'b0; 
    r811 = 1'b0; 
    r812 = 1'b0; 
    r813 = 1'b0; 
    r814 = 1'b0; 
    r815 = 1'b0; 
    r816 = 1'b0; 
    r817 = 1'b0; 
    r818 = 1'b0; 
    r819 = 1'b0; 
    r820 = 1'b0; 
    r821 = 1'b0; 
    r822 = 1'b0; 
    r823 = 1'b0; 
    r824 = 1'b0; 
    r825 = 1'b0; 
    r826 = 1'b0; 
    r827 = 1'b0; 
    r828 = 1'b0; 
    r829 = 1'b0; 
    r830 = 1'b0; 
    r831 = 1'b0; 
    r832 = 1'b0; 
    r833 = 1'b0; 
    r834 = 1'b0; 
    r835 = 1'b0; 
    r836 = 1'b0; 
    r837 = 1'b0; 
    r838 = 1'b0; 
    r839 = 1'b0; 
    r840 = 1'b0; 
    r841 = 1'b0; 
    r842 = 1'b0; 
    r843 = 1'b0; 
    r844 = 1'b0; 
    r845 = 1'b0; 
    r846 = 1'b0; 
    r847 = 1'b0; 
    r848 = 1'b0; 
    r849 = 1'b0; 
    r850 = 1'b0; 
    r851 = 1'b0; 
    r852 = 1'b0; 
    r853 = 1'b0; 
    r854 = 1'b0; 
    r855 = 1'b0; 
    r856 = 1'b0; 
    r857 = 1'b0; 
    r858 = 1'b0; 
    r859 = 1'b0; 
    r860 = 1'b0; 
    r861 = 1'b0; 
    r862 = 1'b0; 
    r863 = 1'b0; 
    r864 = 1'b0; 
    r865 = 1'b0; 
    r866 = 1'b0; 
    r867 = 1'b0; 
    r868 = 1'b0; 
    r869 = 1'b0; 
    r870 = 1'b0; 
    r871 = 1'b0; 
    r872 = 1'b0; 
    r873 = 1'b0; 
    r874 = 1'b0; 
    r875 = 1'b0; 
    r876 = 1'b0; 
    r877 = 1'b0; 
    r878 = 1'b0; 
    r879 = 1'b0; 
    r880 = 1'b0; 
    r881 = 1'b0; 
    r882 = 1'b0; 
    r883 = 1'b0; 
    r884 = 1'b0; 
    r885 = 1'b0; 
    r886 = 1'b0; 
    r887 = 1'b0; 
    r888 = 1'b0; 
    r889 = 1'b0; 
    r890 = 1'b0; 
    r891 = 1'b0; 
    r892 = 1'b0; 
    r893 = 1'b0; 
    r894 = 1'b0; 
    r895 = 1'b0; 
    r896 = 1'b0; 
    r897 = 1'b0; 
    r898 = 1'b0; 
    r899 = 1'b0; 
    r900 = 1'b0; 
    r901 = 1'b0; 
    r902 = 1'b0; 
    r903 = 1'b0; 
    r904 = 1'b0; 
    r905 = 1'b0; 
    r906 = 1'b0; 
    r907 = 1'b0; 
    r908 = 1'b0; 
    r909 = 1'b0; 
    r910 = 1'b0; 
    r911 = 1'b0; 
    r912 = 1'b0; 
    r913 = 1'b0; 
    r914 = 1'b0; 
    r915 = 1'b0; 
    r916 = 1'b0; 
    r917 = 1'b0; 
    r918 = 1'b0; 
    r919 = 1'b0; 
    r920 = 1'b0; 
    r921 = 1'b0; 
    r922 = 1'b0; 
    r923 = 1'b0; 
    r924 = 1'b0; 
    r925 = 1'b0; 
    r926 = 1'b0; 
    r927 = 1'b0; 
    r928 = 1'b0; 
    r929 = 1'b0; 
    r930 = 1'b0; 
    r931 = 1'b0; 
    r932 = 1'b0; 
    r933 = 1'b0; 
    r934 = 1'b0; 
    r935 = 1'b0; 
    r936 = 1'b0; 
    r937 = 1'b0; 
    r938 = 1'b0; 
    r939 = 1'b0; 
    r940 = 1'b0; 
    r941 = 1'b0; 
    r942 = 1'b0; 
    r943 = 1'b0; 
    r944 = 1'b0; 
    r945 = 1'b0; 
    r946 = 1'b0; 
    r947 = 1'b0; 
    r948 = 1'b0; 
    r949 = 1'b0; 
    r950 = 1'b0; 
    r951 = 1'b0; 
    r952 = 1'b0; 
    r953 = 1'b0; 
    r954 = 1'b0; 
    r955 = 1'b0; 
    r956 = 1'b0; 
    r957 = 1'b0; 
    r958 = 1'b0; 
    r959 = 1'b0; 
    r960 = 1'b0; 
    r961 = 1'b0; 
    r962 = 1'b0; 
    r963 = 1'b0; 
    r964 = 1'b0; 
    r965 = 1'b0; 
    r966 = 1'b0; 
    r967 = 1'b0; 
    r968 = 1'b0; 
    r969 = 1'b0; 
    r970 = 1'b0; 
    r971 = 1'b0; 
    r972 = 1'b0; 
    r973 = 1'b0; 
    r974 = 1'b0; 
    r975 = 1'b0; 
    r976 = 1'b0; 
    r977 = 1'b0; 
    r978 = 1'b0; 
    r979 = 1'b0; 
    r980 = 1'b0; 
    r981 = 1'b0; 
    r982 = 1'b0; 
    r983 = 1'b0; 
    r984 = 1'b0; 
    r985 = 1'b0; 
    r986 = 1'b0; 
    r987 = 1'b0; 
    r988 = 1'b0; 
    r989 = 1'b0; 
    r990 = 1'b0; 
    r991 = 1'b0; 
    r992 = 1'b0; 
    r993 = 1'b0; 
    r994 = 1'b0; 
    r995 = 1'b0; 
    r996 = 1'b0; 
    r997 = 1'b0; 
    r998 = 1'b0; 
    r999 = 1'b0; 
    $monitor("%t %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b  ", $time, w_000_000, w_000_001, w_000_002, w_000_003, w_000_004, w_000_005, w_000_006, w_000_007, w_000_008, w_000_009, w_000_010, w_000_011, w_000_012, w_000_013, w_000_014, w_000_015, w_000_016, w_000_017, w_000_018, w_000_019, w_000_020, w_000_021, w_000_022, w_000_023, w_000_024, w_000_025, w_000_026, w_000_027, w_000_028, w_000_029, w_000_030, w_000_031, w_000_032, w_000_033, w_000_034, w_000_035, w_000_036, w_000_037, w_000_038, w_000_039, w_000_040, w_000_041, w_000_042, w_000_043, w_000_044, w_000_045, w_000_046, w_000_047, w_000_048, w_000_049, w_000_050, w_000_051, w_000_052, w_000_053, w_000_054, w_000_055, w_000_056, w_000_057, w_000_058, w_000_059, w_000_060, w_000_061, w_000_062, w_000_063, w_000_064, w_000_065, w_000_066, w_000_067, w_000_068, w_000_069, w_000_070, w_000_071, w_000_072, w_000_073, w_000_074, w_000_075, w_000_076, w_000_077, w_000_078, w_000_079, w_000_080, w_000_081, w_000_082, w_000_083, w_000_084, w_000_085, w_000_086, w_000_087, w_000_088, w_000_089, w_000_090, w_000_091, w_000_092, w_000_093, w_000_094, w_000_095, w_000_096, w_000_097, w_000_098, w_000_099, w_000_100, w_000_101, w_000_102, w_000_103, w_000_104, w_000_105, w_000_106, w_000_107, w_000_108, w_000_109, w_000_110, w_000_111, w_000_112, w_000_113, w_000_114, w_000_115, w_000_116, w_000_117, w_000_118, w_000_119, w_000_120, w_000_121, w_000_122, w_000_123, w_000_124, w_000_125, w_000_126, w_000_127, w_000_128, w_000_129, w_000_130, w_000_131, w_000_132, w_000_133, w_000_134, w_000_135, w_000_136, w_000_137, w_000_138, w_000_139, w_000_140, w_000_141, w_000_142, w_000_143, w_000_144, w_000_145, w_000_146, w_000_147, w_000_148, w_000_149, w_000_150, w_000_151, w_000_152, w_000_153, w_000_154, w_000_155, w_000_156, w_000_157, w_000_158, w_000_159, w_000_160, w_000_161, w_000_162, w_000_163, w_000_164, w_000_165, w_000_166, w_000_167, w_000_168, w_000_169, w_000_170, w_000_171, w_000_172, w_000_173, w_000_174, w_000_175, w_000_176, w_000_177, w_000_178, w_000_179, w_000_180, w_000_181, w_000_182, w_000_183, w_000_184, w_000_185, w_000_186, w_000_187, w_000_188, w_000_189, w_000_190, w_000_191, w_000_192, w_000_193, w_000_194, w_000_195, w_000_196, w_000_197, w_000_198, w_000_199, w_000_200, w_000_201, w_000_202, w_000_203, w_000_204, w_000_205, w_000_206, w_000_207, w_000_208, w_000_209, w_000_210, w_000_211, w_000_212, w_000_213, w_000_214, w_000_215, w_000_216, w_000_217, w_000_218, w_000_219, w_000_220, w_000_221, w_000_222, w_000_223, w_000_224, w_000_225, w_000_226, w_000_227, w_000_228, w_000_229, w_000_230, w_000_231, w_000_232, w_000_233, w_000_234, w_000_235, w_000_236, w_000_237, w_000_238, w_000_239, w_000_240, w_000_241, w_000_242, w_000_243, w_000_244, w_000_245, w_000_246, w_000_247, w_000_248, w_000_249, w_000_250, w_000_251, w_000_252, w_000_253, w_000_254, w_000_255, w_000_256, w_000_257, w_000_258, w_000_259, w_000_260, w_000_261, w_000_262, w_000_263, w_000_264, w_000_265, w_000_266, w_000_267, w_000_268, w_000_269, w_000_270, w_000_271, w_000_272, w_000_273, w_000_274, w_000_275, w_000_276, w_000_277, w_000_278, w_000_279, w_000_280, w_000_281, w_000_282, w_000_283, w_000_284, w_000_285, w_000_286, w_000_287, w_000_288, w_000_289, w_000_290, w_000_291, w_000_292, w_000_293, w_000_294, w_000_295, w_000_296, w_000_297, w_000_298, w_000_299, w_000_300, w_000_301, w_000_302, w_000_303, w_000_304, w_000_305, w_000_306, w_000_307, w_000_308, w_000_309, w_000_310, w_000_311, w_000_312, w_000_313, w_000_314, w_000_315, w_000_316, w_000_317, w_000_318, w_000_319, w_000_320, w_000_321, w_000_322, w_000_323, w_000_324, w_000_325, w_000_326, w_000_327, w_000_328, w_000_329, w_000_330, w_000_331, w_000_332, w_000_333, w_000_334, w_000_335, w_000_336, w_000_337, w_000_338, w_000_339, w_000_340, w_000_341, w_000_342, w_000_343, w_000_344, w_000_345, w_000_346, w_000_347, w_000_348, w_000_349, w_000_350, w_000_351, w_000_352, w_000_353, w_000_354, w_000_355, w_000_356, w_000_357, w_000_358, w_000_359, w_000_360, w_000_361, w_000_362, w_000_363, w_000_364, w_000_365, w_000_366, w_000_367, w_000_368, w_000_369, w_000_370, w_000_371, w_000_372, w_000_373, w_000_374, w_000_375, w_000_376, w_000_377, w_000_378, w_000_379, w_000_380, w_000_381, w_000_382, w_000_383, w_000_384, w_000_385, w_000_386, w_000_387, w_000_388, w_000_389, w_000_390, w_000_391, w_000_392, w_000_393, w_000_394, w_000_395, w_000_396, w_000_397, w_000_398, w_000_399, w_000_400, w_000_401, w_000_402, w_000_403, w_000_404, w_000_405, w_000_406, w_000_407, w_000_408, w_000_409, w_000_410, w_000_411, w_000_412, w_000_413, w_000_414, w_000_415, w_000_416, w_000_417, w_000_418, w_000_419, w_000_420, w_000_421, w_000_422, w_000_423, w_000_424, w_000_425, w_000_426, w_000_427, w_000_428, w_000_429, w_000_430, w_000_431, w_000_432, w_000_433, w_000_434, w_000_435, w_000_436, w_000_437, w_000_438, w_000_439, w_000_440, w_000_441, w_000_442, w_000_443, w_000_444, w_000_445, w_000_446, w_000_447, w_000_448, w_000_449, w_000_450, w_000_451, w_000_452, w_000_453, w_000_454, w_000_455, w_000_456, w_000_457, w_000_458, w_000_459, w_000_460, w_000_461, w_000_462, w_000_463, w_000_464, w_000_465, w_000_466, w_000_467, w_000_468, w_000_469, w_000_470, w_000_471, w_000_472, w_000_473, w_000_474, w_000_475, w_000_476, w_000_477, w_000_478, w_000_479, w_000_480, w_000_481, w_000_482, w_000_483, w_000_484, w_000_485, w_000_486, w_000_487, w_000_488, w_000_489, w_000_490, w_000_491, w_000_492, w_000_493, w_000_494, w_000_495, w_000_496, w_000_497, w_000_498, w_000_499, w_000_500, w_000_501, w_000_502, w_000_503, w_000_504, w_000_505, w_000_506, w_000_507, w_000_508, w_000_509, w_000_510, w_000_511, w_000_512, w_000_513, w_000_514, w_000_515, w_000_516, w_000_517, w_000_518, w_000_519, w_000_520, w_000_521, w_000_522, w_000_523, w_000_524, w_000_525, w_000_526, w_000_527, w_000_528, w_000_529, w_000_530, w_000_531, w_000_532, w_000_533, w_000_534, w_000_535, w_000_536, w_000_537, w_000_538, w_000_539, w_000_540, w_000_541, w_000_542, w_000_543, w_000_544, w_000_545, w_000_546, w_000_547, w_000_548, w_000_549, w_000_550, w_000_551, w_000_552, w_000_553, w_000_554, w_000_555, w_000_556, w_000_557, w_000_558, w_000_559, w_000_560, w_000_561, w_000_562, w_000_563, w_000_564, w_000_565, w_000_566, w_000_567, w_000_568, w_000_569, w_000_570, w_000_571, w_000_572, w_000_573, w_000_574, w_000_575, w_000_576, w_000_577, w_000_578, w_000_579, w_000_580, w_000_581, w_000_582, w_000_583, w_000_584, w_000_585, w_000_586, w_000_587, w_000_588, w_000_589, w_000_590, w_000_591, w_000_592, w_000_593, w_000_594, w_000_595, w_000_596, w_000_597, w_000_598, w_000_599, w_000_600, w_000_601, w_000_602, w_000_603, w_000_604, w_000_605, w_000_606, w_000_607, w_000_608, w_000_609, w_000_610, w_000_611, w_000_612, w_000_613, w_000_614, w_000_615, w_000_616, w_000_617, w_000_618, w_000_619, w_000_620, w_000_621, w_000_622, w_000_623, w_000_624, w_000_625, w_000_626, w_000_627, w_000_628, w_000_629, w_000_630, w_000_631, w_000_632, w_000_633, w_000_634, w_000_635, w_000_636, w_000_637, w_000_638, w_000_639, w_000_640, w_000_641, w_000_642, w_000_643, w_000_644, w_000_645, w_000_646, w_000_647, w_000_648, w_000_649, w_000_650, w_000_651, w_000_652, w_000_653, w_000_654, w_000_655, w_000_656, w_000_657, w_000_658, w_000_659, w_000_660, w_000_661, w_000_662, w_000_663, w_000_664, w_000_665, w_000_666, w_000_667, w_000_668, w_000_669, w_000_670, w_000_671, w_000_672, w_000_673, w_000_674, w_000_675, w_000_676, w_000_677, w_000_678, w_000_679, w_000_680, w_000_681, w_000_682, w_000_683, w_000_684, w_000_685, w_000_686, w_000_687, w_000_688, w_000_689, w_000_690, w_000_691, w_000_692, w_000_693, w_000_694, w_000_695, w_000_696, w_000_697, w_000_698, w_000_699, w_000_700, w_000_701, w_000_702, w_000_703, w_000_704, w_000_705, w_000_706, w_000_707, w_000_708, w_000_709, w_000_710, w_000_711, w_000_712, w_000_713, w_000_714, w_000_715, w_000_716, w_000_717, w_000_718, w_000_719, w_000_720, w_000_721, w_000_722, w_000_723, w_000_724, w_000_725, w_000_726, w_000_727, w_000_728, w_000_729, w_000_730, w_000_731, w_000_732, w_000_733, w_000_734, w_000_735, w_000_736, w_000_737, w_000_738, w_000_739, w_000_740, w_000_741, w_000_742, w_000_743, w_000_744, w_000_745, w_000_746, w_000_747, w_000_748, w_000_749, w_000_750, w_000_751, w_000_752, w_000_753, w_000_754, w_000_755, w_000_756, w_000_757, w_000_758, w_000_759, w_000_760, w_000_761, w_000_762, w_000_763, w_000_764, w_000_765, w_000_766, w_000_767, w_000_768, w_000_769, w_000_770, w_000_771, w_000_772, w_000_773, w_000_774, w_000_775, w_000_776, w_000_777, w_000_778, w_000_779, w_000_780, w_000_781, w_000_782, w_000_783, w_000_784, w_000_785, w_000_786, w_000_787, w_000_788, w_000_789, w_000_790, w_000_791, w_000_792, w_000_793, w_000_794, w_000_795, w_000_796, w_000_797, w_000_798, w_000_799, w_000_800, w_000_801, w_000_802, w_000_803, w_000_804, w_000_805, w_000_806, w_000_807, w_000_808, w_000_809, w_000_810, w_000_811, w_000_812, w_000_813, w_000_814, w_000_815, w_000_816, w_000_817, w_000_818, w_000_819, w_000_820, w_000_821, w_000_822, w_000_823, w_000_824, w_000_825, w_000_826, w_000_827, w_000_828, w_000_829, w_000_830, w_000_831, w_000_832, w_000_833, w_000_834, w_000_835, w_000_836, w_000_837, w_000_838, w_000_839, w_000_840, w_000_841, w_000_842, w_000_843, w_000_844, w_000_845, w_000_846, w_000_847, w_000_848, w_000_849, w_000_850, w_000_851, w_000_852, w_000_853, w_000_854, w_000_855, w_000_856, w_000_857, w_000_858, w_000_859, w_000_860, w_000_861, w_000_862, w_000_863, w_000_864, w_000_865, w_000_866, w_000_867, w_000_868, w_000_869, w_000_870, w_000_871, w_000_872, w_000_873, w_000_874, w_000_875, w_000_876, w_000_877, w_000_878, w_000_879, w_000_880, w_000_881, w_000_882, w_000_883, w_000_884, w_000_885, w_000_886, w_000_887, w_000_888, w_000_889, w_000_890, w_000_891, w_000_892, w_000_893, w_000_894, w_000_895, w_000_896, w_000_897, w_000_898, w_000_899, w_000_900, w_000_901, w_000_902, w_000_903, w_000_904, w_000_905, w_000_906, w_000_907, w_000_908, w_000_909, w_000_910, w_000_911, w_000_912, w_000_913, w_000_914, w_000_915, w_000_916, w_000_917, w_000_918, w_000_919, w_000_920, w_000_921, w_000_922, w_000_923, w_000_924, w_000_925, w_000_926, w_000_927, w_000_928, w_000_929, w_000_930, w_000_931, w_000_932, w_000_933, w_000_934, w_000_935, w_000_936, w_000_937, w_000_938, w_000_939, w_000_940, w_000_941, w_000_942, w_000_943, w_000_944, w_000_945, w_000_946, w_000_947, w_000_948, w_000_949, w_000_950, w_000_951, w_000_952, w_000_953, w_000_954, w_000_955, w_000_956, w_000_957, w_000_958, w_000_959, w_000_960, w_000_961, w_000_962, w_000_963, w_000_964, w_000_965, w_000_966, w_000_967, w_000_968, w_000_969, w_000_970, w_000_971, w_000_972, w_000_973, w_000_974, w_000_975, w_000_976, w_000_977, w_000_978, w_000_979, w_000_980, w_000_981, w_000_982, w_000_983, w_000_984, w_000_985, w_000_986, w_000_987, w_000_988, w_000_989, w_000_990, w_000_991, w_000_992, w_000_993, w_000_994, w_000_995, w_000_996, w_000_997, w_000_998, w_000_999, w_1000_000, w_1000_001, w_1000_002, w_1000_003, w_1000_004, w_1000_005, w_1000_006, w_1000_007, w_1000_008, w_1000_009, w_1000_010, w_1000_011, w_1000_012, w_1000_013, w_1000_014, w_1000_015, w_1000_016, w_1000_017, w_1000_018, w_1000_019, w_1000_020, w_1000_021, w_1000_022, w_1000_023, w_1000_024, w_1000_025, w_1000_026, w_1000_027, w_1000_028, w_1000_029, w_1000_030, w_1000_031, w_1000_032, w_1000_033, w_1000_034, w_1000_035, w_1000_036, w_1000_037, w_1000_038, w_1000_039, w_1000_040, w_1000_041, w_1000_042, w_1000_043, w_1000_044, w_1000_045, w_1000_046, w_1000_047, w_1000_048, w_1000_049, w_1000_050, w_1000_051, w_1000_052, w_1000_053, w_1000_054, w_1000_055, w_1000_056, w_1000_057, w_1000_058, w_1000_059, w_1000_060, w_1000_061, w_1000_062, w_1000_063, w_1000_064, w_1000_065, w_1000_066, w_1000_067, w_1000_068, w_1000_069, w_1000_070, w_1000_071, w_1000_072, w_1000_073, w_1000_074, w_1000_075, w_1000_076, w_1000_077, w_1000_078, w_1000_079, w_1000_080, w_1000_081, w_1000_082, w_1000_083, w_1000_084, w_1000_085, w_1000_086, w_1000_087, w_1000_088, w_1000_089, w_1000_090, w_1000_091, w_1000_092, w_1000_093, w_1000_094, w_1000_095, w_1000_096, w_1000_097, w_1000_098, w_1000_099, w_1000_100, w_1000_101, w_1000_102, w_1000_103, w_1000_104, w_1000_105, w_1000_106, w_1000_107, w_1000_108, w_1000_109, w_1000_110, w_1000_111, w_1000_112, w_1000_113, w_1000_114, w_1000_115, w_1000_116, w_1000_117, w_1000_118, w_1000_119, w_1000_120, w_1000_121, w_1000_122, w_1000_123, w_1000_124, w_1000_125, w_1000_126, w_1000_127, w_1000_128, w_1000_129, w_1000_130, w_1000_131, w_1000_132, w_1000_133, w_1000_134, w_1000_135, w_1000_136, w_1000_137, w_1000_138, w_1000_139, w_1000_140, w_1000_141, w_1000_142, w_1000_143, w_1000_144, w_1000_145, w_1000_146, w_1000_147, w_1000_148, w_1000_149, w_1000_150, w_1000_151, w_1000_152, w_1000_153, w_1000_154, w_1000_155, w_1000_156, w_1000_157, w_1000_158, w_1000_159, w_1000_160, w_1000_161, w_1000_162, w_1000_163, w_1000_164, w_1000_165, w_1000_166, w_1000_167, w_1000_168, w_1000_169, w_1000_170, w_1000_171, w_1000_172, w_1000_173, w_1000_174, w_1000_175, w_1000_176, w_1000_177, w_1000_178, w_1000_179, w_1000_180, w_1000_181, w_1000_182, w_1000_183, w_1000_184, w_1000_185);
    #100;
    $finish;
  end
  always #1 r0 = ~r0;
  always #2 r1 = ~r1;
  always #4 r2 = ~r2;
  always #8 r3 = ~r3;
  always #16 r4 = ~r4;
  always #32 r5 = ~r5;
  always #64 r6 = ~r6;
  always #128 r7 = ~r7;
  always #256 r8 = ~r8;
  always #512 r9 = ~r9;
  always #1024 r10 = ~r10;
  always #2048 r11 = ~r11;
  always #4096 r12 = ~r12;
  always #8192 r13 = ~r13;
  always #16384 r14 = ~r14;
  always #32768 r15 = ~r15;
  always #65536 r16 = ~r16;
  always #131072 r17 = ~r17;
  always #262144 r18 = ~r18;
  always #524288 r19 = ~r19;
  always #1048576 r20 = ~r20;
  always #2097152 r21 = ~r21;
  always #4194304 r22 = ~r22;
  always #8388608 r23 = ~r23;
  always #16777216 r24 = ~r24;
  always #33554432 r25 = ~r25;
  always #67108864 r26 = ~r26;
  always #134217728 r27 = ~r27;
  always #268435456 r28 = ~r28;
  always #536870912 r29 = ~r29;
  always #1073741824 r30 = ~r30;
  always #2147483648 r31 = ~r31;
  always #4294967296 r32 = ~r32;
  always #8589934592 r33 = ~r33;
  always #17179869184 r34 = ~r34;
  always #34359738368 r35 = ~r35;
  always #68719476736 r36 = ~r36;
  always #137438953472 r37 = ~r37;
  always #274877906944 r38 = ~r38;
  always #549755813888 r39 = ~r39;
  always #1099511627776 r40 = ~r40;
  always #2199023255552 r41 = ~r41;
  always #4398046511104 r42 = ~r42;
  always #8796093022208 r43 = ~r43;
  always #17592186044416 r44 = ~r44;
  always #35184372088832 r45 = ~r45;
  always #70368744177664 r46 = ~r46;
  always #140737488355328 r47 = ~r47;
  always #281474976710656 r48 = ~r48;
  always #562949953421312 r49 = ~r49;
  always #1125899906842624 r50 = ~r50;
  always #2251799813685248 r51 = ~r51;
  always #4503599627370496 r52 = ~r52;
  always #9007199254740992 r53 = ~r53;
  always #18014398509481984 r54 = ~r54;
  always #36028797018963968 r55 = ~r55;
  always #72057594037927936 r56 = ~r56;
  always #144115188075855872 r57 = ~r57;
  always #288230376151711744 r58 = ~r58;
  always #576460752303423488 r59 = ~r59;
  always #1152921504606846976 r60 = ~r60;
  always #2305843009213693952 r61 = ~r61;
  always #4611686018427387904 r62 = ~r62;
  always #9223372036854775808 r63 = ~r63;
  always #1 r64 = ~r64;
  always #2 r65 = ~r65;
  always #4 r66 = ~r66;
  always #8 r67 = ~r67;
  always #16 r68 = ~r68;
  always #32 r69 = ~r69;
  always #64 r70 = ~r70;
  always #128 r71 = ~r71;
  always #256 r72 = ~r72;
  always #512 r73 = ~r73;
  always #1024 r74 = ~r74;
  always #2048 r75 = ~r75;
  always #4096 r76 = ~r76;
  always #8192 r77 = ~r77;
  always #16384 r78 = ~r78;
  always #32768 r79 = ~r79;
  always #65536 r80 = ~r80;
  always #131072 r81 = ~r81;
  always #262144 r82 = ~r82;
  always #524288 r83 = ~r83;
  always #1048576 r84 = ~r84;
  always #2097152 r85 = ~r85;
  always #4194304 r86 = ~r86;
  always #8388608 r87 = ~r87;
  always #16777216 r88 = ~r88;
  always #33554432 r89 = ~r89;
  always #67108864 r90 = ~r90;
  always #134217728 r91 = ~r91;
  always #268435456 r92 = ~r92;
  always #536870912 r93 = ~r93;
  always #1073741824 r94 = ~r94;
  always #2147483648 r95 = ~r95;
  always #4294967296 r96 = ~r96;
  always #8589934592 r97 = ~r97;
  always #17179869184 r98 = ~r98;
  always #34359738368 r99 = ~r99;
  always #68719476736 r100 = ~r100;
  always #137438953472 r101 = ~r101;
  always #274877906944 r102 = ~r102;
  always #549755813888 r103 = ~r103;
  always #1099511627776 r104 = ~r104;
  always #2199023255552 r105 = ~r105;
  always #4398046511104 r106 = ~r106;
  always #8796093022208 r107 = ~r107;
  always #17592186044416 r108 = ~r108;
  always #35184372088832 r109 = ~r109;
  always #70368744177664 r110 = ~r110;
  always #140737488355328 r111 = ~r111;
  always #281474976710656 r112 = ~r112;
  always #562949953421312 r113 = ~r113;
  always #1125899906842624 r114 = ~r114;
  always #2251799813685248 r115 = ~r115;
  always #4503599627370496 r116 = ~r116;
  always #9007199254740992 r117 = ~r117;
  always #18014398509481984 r118 = ~r118;
  always #36028797018963968 r119 = ~r119;
  always #72057594037927936 r120 = ~r120;
  always #144115188075855872 r121 = ~r121;
  always #288230376151711744 r122 = ~r122;
  always #576460752303423488 r123 = ~r123;
  always #1152921504606846976 r124 = ~r124;
  always #2305843009213693952 r125 = ~r125;
  always #4611686018427387904 r126 = ~r126;
  always #9223372036854775808 r127 = ~r127;
  always #1 r128 = ~r128;
  always #2 r129 = ~r129;
  always #4 r130 = ~r130;
  always #8 r131 = ~r131;
  always #16 r132 = ~r132;
  always #32 r133 = ~r133;
  always #64 r134 = ~r134;
  always #128 r135 = ~r135;
  always #256 r136 = ~r136;
  always #512 r137 = ~r137;
  always #1024 r138 = ~r138;
  always #2048 r139 = ~r139;
  always #4096 r140 = ~r140;
  always #8192 r141 = ~r141;
  always #16384 r142 = ~r142;
  always #32768 r143 = ~r143;
  always #65536 r144 = ~r144;
  always #131072 r145 = ~r145;
  always #262144 r146 = ~r146;
  always #524288 r147 = ~r147;
  always #1048576 r148 = ~r148;
  always #2097152 r149 = ~r149;
  always #4194304 r150 = ~r150;
  always #8388608 r151 = ~r151;
  always #16777216 r152 = ~r152;
  always #33554432 r153 = ~r153;
  always #67108864 r154 = ~r154;
  always #134217728 r155 = ~r155;
  always #268435456 r156 = ~r156;
  always #536870912 r157 = ~r157;
  always #1073741824 r158 = ~r158;
  always #2147483648 r159 = ~r159;
  always #4294967296 r160 = ~r160;
  always #8589934592 r161 = ~r161;
  always #17179869184 r162 = ~r162;
  always #34359738368 r163 = ~r163;
  always #68719476736 r164 = ~r164;
  always #137438953472 r165 = ~r165;
  always #274877906944 r166 = ~r166;
  always #549755813888 r167 = ~r167;
  always #1099511627776 r168 = ~r168;
  always #2199023255552 r169 = ~r169;
  always #4398046511104 r170 = ~r170;
  always #8796093022208 r171 = ~r171;
  always #17592186044416 r172 = ~r172;
  always #35184372088832 r173 = ~r173;
  always #70368744177664 r174 = ~r174;
  always #140737488355328 r175 = ~r175;
  always #281474976710656 r176 = ~r176;
  always #562949953421312 r177 = ~r177;
  always #1125899906842624 r178 = ~r178;
  always #2251799813685248 r179 = ~r179;
  always #4503599627370496 r180 = ~r180;
  always #9007199254740992 r181 = ~r181;
  always #18014398509481984 r182 = ~r182;
  always #36028797018963968 r183 = ~r183;
  always #72057594037927936 r184 = ~r184;
  always #144115188075855872 r185 = ~r185;
  always #288230376151711744 r186 = ~r186;
  always #576460752303423488 r187 = ~r187;
  always #1152921504606846976 r188 = ~r188;
  always #2305843009213693952 r189 = ~r189;
  always #4611686018427387904 r190 = ~r190;
  always #9223372036854775808 r191 = ~r191;
  always #1 r192 = ~r192;
  always #2 r193 = ~r193;
  always #4 r194 = ~r194;
  always #8 r195 = ~r195;
  always #16 r196 = ~r196;
  always #32 r197 = ~r197;
  always #64 r198 = ~r198;
  always #128 r199 = ~r199;
  always #256 r200 = ~r200;
  always #512 r201 = ~r201;
  always #1024 r202 = ~r202;
  always #2048 r203 = ~r203;
  always #4096 r204 = ~r204;
  always #8192 r205 = ~r205;
  always #16384 r206 = ~r206;
  always #32768 r207 = ~r207;
  always #65536 r208 = ~r208;
  always #131072 r209 = ~r209;
  always #262144 r210 = ~r210;
  always #524288 r211 = ~r211;
  always #1048576 r212 = ~r212;
  always #2097152 r213 = ~r213;
  always #4194304 r214 = ~r214;
  always #8388608 r215 = ~r215;
  always #16777216 r216 = ~r216;
  always #33554432 r217 = ~r217;
  always #67108864 r218 = ~r218;
  always #134217728 r219 = ~r219;
  always #268435456 r220 = ~r220;
  always #536870912 r221 = ~r221;
  always #1073741824 r222 = ~r222;
  always #2147483648 r223 = ~r223;
  always #4294967296 r224 = ~r224;
  always #8589934592 r225 = ~r225;
  always #17179869184 r226 = ~r226;
  always #34359738368 r227 = ~r227;
  always #68719476736 r228 = ~r228;
  always #137438953472 r229 = ~r229;
  always #274877906944 r230 = ~r230;
  always #549755813888 r231 = ~r231;
  always #1099511627776 r232 = ~r232;
  always #2199023255552 r233 = ~r233;
  always #4398046511104 r234 = ~r234;
  always #8796093022208 r235 = ~r235;
  always #17592186044416 r236 = ~r236;
  always #35184372088832 r237 = ~r237;
  always #70368744177664 r238 = ~r238;
  always #140737488355328 r239 = ~r239;
  always #281474976710656 r240 = ~r240;
  always #562949953421312 r241 = ~r241;
  always #1125899906842624 r242 = ~r242;
  always #2251799813685248 r243 = ~r243;
  always #4503599627370496 r244 = ~r244;
  always #9007199254740992 r245 = ~r245;
  always #18014398509481984 r246 = ~r246;
  always #36028797018963968 r247 = ~r247;
  always #72057594037927936 r248 = ~r248;
  always #144115188075855872 r249 = ~r249;
  always #288230376151711744 r250 = ~r250;
  always #576460752303423488 r251 = ~r251;
  always #1152921504606846976 r252 = ~r252;
  always #2305843009213693952 r253 = ~r253;
  always #4611686018427387904 r254 = ~r254;
  always #9223372036854775808 r255 = ~r255;
  always #1 r256 = ~r256;
  always #2 r257 = ~r257;
  always #4 r258 = ~r258;
  always #8 r259 = ~r259;
  always #16 r260 = ~r260;
  always #32 r261 = ~r261;
  always #64 r262 = ~r262;
  always #128 r263 = ~r263;
  always #256 r264 = ~r264;
  always #512 r265 = ~r265;
  always #1024 r266 = ~r266;
  always #2048 r267 = ~r267;
  always #4096 r268 = ~r268;
  always #8192 r269 = ~r269;
  always #16384 r270 = ~r270;
  always #32768 r271 = ~r271;
  always #65536 r272 = ~r272;
  always #131072 r273 = ~r273;
  always #262144 r274 = ~r274;
  always #524288 r275 = ~r275;
  always #1048576 r276 = ~r276;
  always #2097152 r277 = ~r277;
  always #4194304 r278 = ~r278;
  always #8388608 r279 = ~r279;
  always #16777216 r280 = ~r280;
  always #33554432 r281 = ~r281;
  always #67108864 r282 = ~r282;
  always #134217728 r283 = ~r283;
  always #268435456 r284 = ~r284;
  always #536870912 r285 = ~r285;
  always #1073741824 r286 = ~r286;
  always #2147483648 r287 = ~r287;
  always #4294967296 r288 = ~r288;
  always #8589934592 r289 = ~r289;
  always #17179869184 r290 = ~r290;
  always #34359738368 r291 = ~r291;
  always #68719476736 r292 = ~r292;
  always #137438953472 r293 = ~r293;
  always #274877906944 r294 = ~r294;
  always #549755813888 r295 = ~r295;
  always #1099511627776 r296 = ~r296;
  always #2199023255552 r297 = ~r297;
  always #4398046511104 r298 = ~r298;
  always #8796093022208 r299 = ~r299;
  always #17592186044416 r300 = ~r300;
  always #35184372088832 r301 = ~r301;
  always #70368744177664 r302 = ~r302;
  always #140737488355328 r303 = ~r303;
  always #281474976710656 r304 = ~r304;
  always #562949953421312 r305 = ~r305;
  always #1125899906842624 r306 = ~r306;
  always #2251799813685248 r307 = ~r307;
  always #4503599627370496 r308 = ~r308;
  always #9007199254740992 r309 = ~r309;
  always #18014398509481984 r310 = ~r310;
  always #36028797018963968 r311 = ~r311;
  always #72057594037927936 r312 = ~r312;
  always #144115188075855872 r313 = ~r313;
  always #288230376151711744 r314 = ~r314;
  always #576460752303423488 r315 = ~r315;
  always #1152921504606846976 r316 = ~r316;
  always #2305843009213693952 r317 = ~r317;
  always #4611686018427387904 r318 = ~r318;
  always #9223372036854775808 r319 = ~r319;
  always #1 r320 = ~r320;
  always #2 r321 = ~r321;
  always #4 r322 = ~r322;
  always #8 r323 = ~r323;
  always #16 r324 = ~r324;
  always #32 r325 = ~r325;
  always #64 r326 = ~r326;
  always #128 r327 = ~r327;
  always #256 r328 = ~r328;
  always #512 r329 = ~r329;
  always #1024 r330 = ~r330;
  always #2048 r331 = ~r331;
  always #4096 r332 = ~r332;
  always #8192 r333 = ~r333;
  always #16384 r334 = ~r334;
  always #32768 r335 = ~r335;
  always #65536 r336 = ~r336;
  always #131072 r337 = ~r337;
  always #262144 r338 = ~r338;
  always #524288 r339 = ~r339;
  always #1048576 r340 = ~r340;
  always #2097152 r341 = ~r341;
  always #4194304 r342 = ~r342;
  always #8388608 r343 = ~r343;
  always #16777216 r344 = ~r344;
  always #33554432 r345 = ~r345;
  always #67108864 r346 = ~r346;
  always #134217728 r347 = ~r347;
  always #268435456 r348 = ~r348;
  always #536870912 r349 = ~r349;
  always #1073741824 r350 = ~r350;
  always #2147483648 r351 = ~r351;
  always #4294967296 r352 = ~r352;
  always #8589934592 r353 = ~r353;
  always #17179869184 r354 = ~r354;
  always #34359738368 r355 = ~r355;
  always #68719476736 r356 = ~r356;
  always #137438953472 r357 = ~r357;
  always #274877906944 r358 = ~r358;
  always #549755813888 r359 = ~r359;
  always #1099511627776 r360 = ~r360;
  always #2199023255552 r361 = ~r361;
  always #4398046511104 r362 = ~r362;
  always #8796093022208 r363 = ~r363;
  always #17592186044416 r364 = ~r364;
  always #35184372088832 r365 = ~r365;
  always #70368744177664 r366 = ~r366;
  always #140737488355328 r367 = ~r367;
  always #281474976710656 r368 = ~r368;
  always #562949953421312 r369 = ~r369;
  always #1125899906842624 r370 = ~r370;
  always #2251799813685248 r371 = ~r371;
  always #4503599627370496 r372 = ~r372;
  always #9007199254740992 r373 = ~r373;
  always #18014398509481984 r374 = ~r374;
  always #36028797018963968 r375 = ~r375;
  always #72057594037927936 r376 = ~r376;
  always #144115188075855872 r377 = ~r377;
  always #288230376151711744 r378 = ~r378;
  always #576460752303423488 r379 = ~r379;
  always #1152921504606846976 r380 = ~r380;
  always #2305843009213693952 r381 = ~r381;
  always #4611686018427387904 r382 = ~r382;
  always #9223372036854775808 r383 = ~r383;
  always #1 r384 = ~r384;
  always #2 r385 = ~r385;
  always #4 r386 = ~r386;
  always #8 r387 = ~r387;
  always #16 r388 = ~r388;
  always #32 r389 = ~r389;
  always #64 r390 = ~r390;
  always #128 r391 = ~r391;
  always #256 r392 = ~r392;
  always #512 r393 = ~r393;
  always #1024 r394 = ~r394;
  always #2048 r395 = ~r395;
  always #4096 r396 = ~r396;
  always #8192 r397 = ~r397;
  always #16384 r398 = ~r398;
  always #32768 r399 = ~r399;
  always #65536 r400 = ~r400;
  always #131072 r401 = ~r401;
  always #262144 r402 = ~r402;
  always #524288 r403 = ~r403;
  always #1048576 r404 = ~r404;
  always #2097152 r405 = ~r405;
  always #4194304 r406 = ~r406;
  always #8388608 r407 = ~r407;
  always #16777216 r408 = ~r408;
  always #33554432 r409 = ~r409;
  always #67108864 r410 = ~r410;
  always #134217728 r411 = ~r411;
  always #268435456 r412 = ~r412;
  always #536870912 r413 = ~r413;
  always #1073741824 r414 = ~r414;
  always #2147483648 r415 = ~r415;
  always #4294967296 r416 = ~r416;
  always #8589934592 r417 = ~r417;
  always #17179869184 r418 = ~r418;
  always #34359738368 r419 = ~r419;
  always #68719476736 r420 = ~r420;
  always #137438953472 r421 = ~r421;
  always #274877906944 r422 = ~r422;
  always #549755813888 r423 = ~r423;
  always #1099511627776 r424 = ~r424;
  always #2199023255552 r425 = ~r425;
  always #4398046511104 r426 = ~r426;
  always #8796093022208 r427 = ~r427;
  always #17592186044416 r428 = ~r428;
  always #35184372088832 r429 = ~r429;
  always #70368744177664 r430 = ~r430;
  always #140737488355328 r431 = ~r431;
  always #281474976710656 r432 = ~r432;
  always #562949953421312 r433 = ~r433;
  always #1125899906842624 r434 = ~r434;
  always #2251799813685248 r435 = ~r435;
  always #4503599627370496 r436 = ~r436;
  always #9007199254740992 r437 = ~r437;
  always #18014398509481984 r438 = ~r438;
  always #36028797018963968 r439 = ~r439;
  always #72057594037927936 r440 = ~r440;
  always #144115188075855872 r441 = ~r441;
  always #288230376151711744 r442 = ~r442;
  always #576460752303423488 r443 = ~r443;
  always #1152921504606846976 r444 = ~r444;
  always #2305843009213693952 r445 = ~r445;
  always #4611686018427387904 r446 = ~r446;
  always #9223372036854775808 r447 = ~r447;
  always #1 r448 = ~r448;
  always #2 r449 = ~r449;
  always #4 r450 = ~r450;
  always #8 r451 = ~r451;
  always #16 r452 = ~r452;
  always #32 r453 = ~r453;
  always #64 r454 = ~r454;
  always #128 r455 = ~r455;
  always #256 r456 = ~r456;
  always #512 r457 = ~r457;
  always #1024 r458 = ~r458;
  always #2048 r459 = ~r459;
  always #4096 r460 = ~r460;
  always #8192 r461 = ~r461;
  always #16384 r462 = ~r462;
  always #32768 r463 = ~r463;
  always #65536 r464 = ~r464;
  always #131072 r465 = ~r465;
  always #262144 r466 = ~r466;
  always #524288 r467 = ~r467;
  always #1048576 r468 = ~r468;
  always #2097152 r469 = ~r469;
  always #4194304 r470 = ~r470;
  always #8388608 r471 = ~r471;
  always #16777216 r472 = ~r472;
  always #33554432 r473 = ~r473;
  always #67108864 r474 = ~r474;
  always #134217728 r475 = ~r475;
  always #268435456 r476 = ~r476;
  always #536870912 r477 = ~r477;
  always #1073741824 r478 = ~r478;
  always #2147483648 r479 = ~r479;
  always #4294967296 r480 = ~r480;
  always #8589934592 r481 = ~r481;
  always #17179869184 r482 = ~r482;
  always #34359738368 r483 = ~r483;
  always #68719476736 r484 = ~r484;
  always #137438953472 r485 = ~r485;
  always #274877906944 r486 = ~r486;
  always #549755813888 r487 = ~r487;
  always #1099511627776 r488 = ~r488;
  always #2199023255552 r489 = ~r489;
  always #4398046511104 r490 = ~r490;
  always #8796093022208 r491 = ~r491;
  always #17592186044416 r492 = ~r492;
  always #35184372088832 r493 = ~r493;
  always #70368744177664 r494 = ~r494;
  always #140737488355328 r495 = ~r495;
  always #281474976710656 r496 = ~r496;
  always #562949953421312 r497 = ~r497;
  always #1125899906842624 r498 = ~r498;
  always #2251799813685248 r499 = ~r499;
  always #4503599627370496 r500 = ~r500;
  always #9007199254740992 r501 = ~r501;
  always #18014398509481984 r502 = ~r502;
  always #36028797018963968 r503 = ~r503;
  always #72057594037927936 r504 = ~r504;
  always #144115188075855872 r505 = ~r505;
  always #288230376151711744 r506 = ~r506;
  always #576460752303423488 r507 = ~r507;
  always #1152921504606846976 r508 = ~r508;
  always #2305843009213693952 r509 = ~r509;
  always #4611686018427387904 r510 = ~r510;
  always #9223372036854775808 r511 = ~r511;
  always #1 r512 = ~r512;
  always #2 r513 = ~r513;
  always #4 r514 = ~r514;
  always #8 r515 = ~r515;
  always #16 r516 = ~r516;
  always #32 r517 = ~r517;
  always #64 r518 = ~r518;
  always #128 r519 = ~r519;
  always #256 r520 = ~r520;
  always #512 r521 = ~r521;
  always #1024 r522 = ~r522;
  always #2048 r523 = ~r523;
  always #4096 r524 = ~r524;
  always #8192 r525 = ~r525;
  always #16384 r526 = ~r526;
  always #32768 r527 = ~r527;
  always #65536 r528 = ~r528;
  always #131072 r529 = ~r529;
  always #262144 r530 = ~r530;
  always #524288 r531 = ~r531;
  always #1048576 r532 = ~r532;
  always #2097152 r533 = ~r533;
  always #4194304 r534 = ~r534;
  always #8388608 r535 = ~r535;
  always #16777216 r536 = ~r536;
  always #33554432 r537 = ~r537;
  always #67108864 r538 = ~r538;
  always #134217728 r539 = ~r539;
  always #268435456 r540 = ~r540;
  always #536870912 r541 = ~r541;
  always #1073741824 r542 = ~r542;
  always #2147483648 r543 = ~r543;
  always #4294967296 r544 = ~r544;
  always #8589934592 r545 = ~r545;
  always #17179869184 r546 = ~r546;
  always #34359738368 r547 = ~r547;
  always #68719476736 r548 = ~r548;
  always #137438953472 r549 = ~r549;
  always #274877906944 r550 = ~r550;
  always #549755813888 r551 = ~r551;
  always #1099511627776 r552 = ~r552;
  always #2199023255552 r553 = ~r553;
  always #4398046511104 r554 = ~r554;
  always #8796093022208 r555 = ~r555;
  always #17592186044416 r556 = ~r556;
  always #35184372088832 r557 = ~r557;
  always #70368744177664 r558 = ~r558;
  always #140737488355328 r559 = ~r559;
  always #281474976710656 r560 = ~r560;
  always #562949953421312 r561 = ~r561;
  always #1125899906842624 r562 = ~r562;
  always #2251799813685248 r563 = ~r563;
  always #4503599627370496 r564 = ~r564;
  always #9007199254740992 r565 = ~r565;
  always #18014398509481984 r566 = ~r566;
  always #36028797018963968 r567 = ~r567;
  always #72057594037927936 r568 = ~r568;
  always #144115188075855872 r569 = ~r569;
  always #288230376151711744 r570 = ~r570;
  always #576460752303423488 r571 = ~r571;
  always #1152921504606846976 r572 = ~r572;
  always #2305843009213693952 r573 = ~r573;
  always #4611686018427387904 r574 = ~r574;
  always #9223372036854775808 r575 = ~r575;
  always #1 r576 = ~r576;
  always #2 r577 = ~r577;
  always #4 r578 = ~r578;
  always #8 r579 = ~r579;
  always #16 r580 = ~r580;
  always #32 r581 = ~r581;
  always #64 r582 = ~r582;
  always #128 r583 = ~r583;
  always #256 r584 = ~r584;
  always #512 r585 = ~r585;
  always #1024 r586 = ~r586;
  always #2048 r587 = ~r587;
  always #4096 r588 = ~r588;
  always #8192 r589 = ~r589;
  always #16384 r590 = ~r590;
  always #32768 r591 = ~r591;
  always #65536 r592 = ~r592;
  always #131072 r593 = ~r593;
  always #262144 r594 = ~r594;
  always #524288 r595 = ~r595;
  always #1048576 r596 = ~r596;
  always #2097152 r597 = ~r597;
  always #4194304 r598 = ~r598;
  always #8388608 r599 = ~r599;
  always #16777216 r600 = ~r600;
  always #33554432 r601 = ~r601;
  always #67108864 r602 = ~r602;
  always #134217728 r603 = ~r603;
  always #268435456 r604 = ~r604;
  always #536870912 r605 = ~r605;
  always #1073741824 r606 = ~r606;
  always #2147483648 r607 = ~r607;
  always #4294967296 r608 = ~r608;
  always #8589934592 r609 = ~r609;
  always #17179869184 r610 = ~r610;
  always #34359738368 r611 = ~r611;
  always #68719476736 r612 = ~r612;
  always #137438953472 r613 = ~r613;
  always #274877906944 r614 = ~r614;
  always #549755813888 r615 = ~r615;
  always #1099511627776 r616 = ~r616;
  always #2199023255552 r617 = ~r617;
  always #4398046511104 r618 = ~r618;
  always #8796093022208 r619 = ~r619;
  always #17592186044416 r620 = ~r620;
  always #35184372088832 r621 = ~r621;
  always #70368744177664 r622 = ~r622;
  always #140737488355328 r623 = ~r623;
  always #281474976710656 r624 = ~r624;
  always #562949953421312 r625 = ~r625;
  always #1125899906842624 r626 = ~r626;
  always #2251799813685248 r627 = ~r627;
  always #4503599627370496 r628 = ~r628;
  always #9007199254740992 r629 = ~r629;
  always #18014398509481984 r630 = ~r630;
  always #36028797018963968 r631 = ~r631;
  always #72057594037927936 r632 = ~r632;
  always #144115188075855872 r633 = ~r633;
  always #288230376151711744 r634 = ~r634;
  always #576460752303423488 r635 = ~r635;
  always #1152921504606846976 r636 = ~r636;
  always #2305843009213693952 r637 = ~r637;
  always #4611686018427387904 r638 = ~r638;
  always #9223372036854775808 r639 = ~r639;
  always #1 r640 = ~r640;
  always #2 r641 = ~r641;
  always #4 r642 = ~r642;
  always #8 r643 = ~r643;
  always #16 r644 = ~r644;
  always #32 r645 = ~r645;
  always #64 r646 = ~r646;
  always #128 r647 = ~r647;
  always #256 r648 = ~r648;
  always #512 r649 = ~r649;
  always #1024 r650 = ~r650;
  always #2048 r651 = ~r651;
  always #4096 r652 = ~r652;
  always #8192 r653 = ~r653;
  always #16384 r654 = ~r654;
  always #32768 r655 = ~r655;
  always #65536 r656 = ~r656;
  always #131072 r657 = ~r657;
  always #262144 r658 = ~r658;
  always #524288 r659 = ~r659;
  always #1048576 r660 = ~r660;
  always #2097152 r661 = ~r661;
  always #4194304 r662 = ~r662;
  always #8388608 r663 = ~r663;
  always #16777216 r664 = ~r664;
  always #33554432 r665 = ~r665;
  always #67108864 r666 = ~r666;
  always #134217728 r667 = ~r667;
  always #268435456 r668 = ~r668;
  always #536870912 r669 = ~r669;
  always #1073741824 r670 = ~r670;
  always #2147483648 r671 = ~r671;
  always #4294967296 r672 = ~r672;
  always #8589934592 r673 = ~r673;
  always #17179869184 r674 = ~r674;
  always #34359738368 r675 = ~r675;
  always #68719476736 r676 = ~r676;
  always #137438953472 r677 = ~r677;
  always #274877906944 r678 = ~r678;
  always #549755813888 r679 = ~r679;
  always #1099511627776 r680 = ~r680;
  always #2199023255552 r681 = ~r681;
  always #4398046511104 r682 = ~r682;
  always #8796093022208 r683 = ~r683;
  always #17592186044416 r684 = ~r684;
  always #35184372088832 r685 = ~r685;
  always #70368744177664 r686 = ~r686;
  always #140737488355328 r687 = ~r687;
  always #281474976710656 r688 = ~r688;
  always #562949953421312 r689 = ~r689;
  always #1125899906842624 r690 = ~r690;
  always #2251799813685248 r691 = ~r691;
  always #4503599627370496 r692 = ~r692;
  always #9007199254740992 r693 = ~r693;
  always #18014398509481984 r694 = ~r694;
  always #36028797018963968 r695 = ~r695;
  always #72057594037927936 r696 = ~r696;
  always #144115188075855872 r697 = ~r697;
  always #288230376151711744 r698 = ~r698;
  always #576460752303423488 r699 = ~r699;
  always #1152921504606846976 r700 = ~r700;
  always #2305843009213693952 r701 = ~r701;
  always #4611686018427387904 r702 = ~r702;
  always #9223372036854775808 r703 = ~r703;
  always #1 r704 = ~r704;
  always #2 r705 = ~r705;
  always #4 r706 = ~r706;
  always #8 r707 = ~r707;
  always #16 r708 = ~r708;
  always #32 r709 = ~r709;
  always #64 r710 = ~r710;
  always #128 r711 = ~r711;
  always #256 r712 = ~r712;
  always #512 r713 = ~r713;
  always #1024 r714 = ~r714;
  always #2048 r715 = ~r715;
  always #4096 r716 = ~r716;
  always #8192 r717 = ~r717;
  always #16384 r718 = ~r718;
  always #32768 r719 = ~r719;
  always #65536 r720 = ~r720;
  always #131072 r721 = ~r721;
  always #262144 r722 = ~r722;
  always #524288 r723 = ~r723;
  always #1048576 r724 = ~r724;
  always #2097152 r725 = ~r725;
  always #4194304 r726 = ~r726;
  always #8388608 r727 = ~r727;
  always #16777216 r728 = ~r728;
  always #33554432 r729 = ~r729;
  always #67108864 r730 = ~r730;
  always #134217728 r731 = ~r731;
  always #268435456 r732 = ~r732;
  always #536870912 r733 = ~r733;
  always #1073741824 r734 = ~r734;
  always #2147483648 r735 = ~r735;
  always #4294967296 r736 = ~r736;
  always #8589934592 r737 = ~r737;
  always #17179869184 r738 = ~r738;
  always #34359738368 r739 = ~r739;
  always #68719476736 r740 = ~r740;
  always #137438953472 r741 = ~r741;
  always #274877906944 r742 = ~r742;
  always #549755813888 r743 = ~r743;
  always #1099511627776 r744 = ~r744;
  always #2199023255552 r745 = ~r745;
  always #4398046511104 r746 = ~r746;
  always #8796093022208 r747 = ~r747;
  always #17592186044416 r748 = ~r748;
  always #35184372088832 r749 = ~r749;
  always #70368744177664 r750 = ~r750;
  always #140737488355328 r751 = ~r751;
  always #281474976710656 r752 = ~r752;
  always #562949953421312 r753 = ~r753;
  always #1125899906842624 r754 = ~r754;
  always #2251799813685248 r755 = ~r755;
  always #4503599627370496 r756 = ~r756;
  always #9007199254740992 r757 = ~r757;
  always #18014398509481984 r758 = ~r758;
  always #36028797018963968 r759 = ~r759;
  always #72057594037927936 r760 = ~r760;
  always #144115188075855872 r761 = ~r761;
  always #288230376151711744 r762 = ~r762;
  always #576460752303423488 r763 = ~r763;
  always #1152921504606846976 r764 = ~r764;
  always #2305843009213693952 r765 = ~r765;
  always #4611686018427387904 r766 = ~r766;
  always #9223372036854775808 r767 = ~r767;
  always #1 r768 = ~r768;
  always #2 r769 = ~r769;
  always #4 r770 = ~r770;
  always #8 r771 = ~r771;
  always #16 r772 = ~r772;
  always #32 r773 = ~r773;
  always #64 r774 = ~r774;
  always #128 r775 = ~r775;
  always #256 r776 = ~r776;
  always #512 r777 = ~r777;
  always #1024 r778 = ~r778;
  always #2048 r779 = ~r779;
  always #4096 r780 = ~r780;
  always #8192 r781 = ~r781;
  always #16384 r782 = ~r782;
  always #32768 r783 = ~r783;
  always #65536 r784 = ~r784;
  always #131072 r785 = ~r785;
  always #262144 r786 = ~r786;
  always #524288 r787 = ~r787;
  always #1048576 r788 = ~r788;
  always #2097152 r789 = ~r789;
  always #4194304 r790 = ~r790;
  always #8388608 r791 = ~r791;
  always #16777216 r792 = ~r792;
  always #33554432 r793 = ~r793;
  always #67108864 r794 = ~r794;
  always #134217728 r795 = ~r795;
  always #268435456 r796 = ~r796;
  always #536870912 r797 = ~r797;
  always #1073741824 r798 = ~r798;
  always #2147483648 r799 = ~r799;
  always #4294967296 r800 = ~r800;
  always #8589934592 r801 = ~r801;
  always #17179869184 r802 = ~r802;
  always #34359738368 r803 = ~r803;
  always #68719476736 r804 = ~r804;
  always #137438953472 r805 = ~r805;
  always #274877906944 r806 = ~r806;
  always #549755813888 r807 = ~r807;
  always #1099511627776 r808 = ~r808;
  always #2199023255552 r809 = ~r809;
  always #4398046511104 r810 = ~r810;
  always #8796093022208 r811 = ~r811;
  always #17592186044416 r812 = ~r812;
  always #35184372088832 r813 = ~r813;
  always #70368744177664 r814 = ~r814;
  always #140737488355328 r815 = ~r815;
  always #281474976710656 r816 = ~r816;
  always #562949953421312 r817 = ~r817;
  always #1125899906842624 r818 = ~r818;
  always #2251799813685248 r819 = ~r819;
  always #4503599627370496 r820 = ~r820;
  always #9007199254740992 r821 = ~r821;
  always #18014398509481984 r822 = ~r822;
  always #36028797018963968 r823 = ~r823;
  always #72057594037927936 r824 = ~r824;
  always #144115188075855872 r825 = ~r825;
  always #288230376151711744 r826 = ~r826;
  always #576460752303423488 r827 = ~r827;
  always #1152921504606846976 r828 = ~r828;
  always #2305843009213693952 r829 = ~r829;
  always #4611686018427387904 r830 = ~r830;
  always #9223372036854775808 r831 = ~r831;
  always #1 r832 = ~r832;
  always #2 r833 = ~r833;
  always #4 r834 = ~r834;
  always #8 r835 = ~r835;
  always #16 r836 = ~r836;
  always #32 r837 = ~r837;
  always #64 r838 = ~r838;
  always #128 r839 = ~r839;
  always #256 r840 = ~r840;
  always #512 r841 = ~r841;
  always #1024 r842 = ~r842;
  always #2048 r843 = ~r843;
  always #4096 r844 = ~r844;
  always #8192 r845 = ~r845;
  always #16384 r846 = ~r846;
  always #32768 r847 = ~r847;
  always #65536 r848 = ~r848;
  always #131072 r849 = ~r849;
  always #262144 r850 = ~r850;
  always #524288 r851 = ~r851;
  always #1048576 r852 = ~r852;
  always #2097152 r853 = ~r853;
  always #4194304 r854 = ~r854;
  always #8388608 r855 = ~r855;
  always #16777216 r856 = ~r856;
  always #33554432 r857 = ~r857;
  always #67108864 r858 = ~r858;
  always #134217728 r859 = ~r859;
  always #268435456 r860 = ~r860;
  always #536870912 r861 = ~r861;
  always #1073741824 r862 = ~r862;
  always #2147483648 r863 = ~r863;
  always #4294967296 r864 = ~r864;
  always #8589934592 r865 = ~r865;
  always #17179869184 r866 = ~r866;
  always #34359738368 r867 = ~r867;
  always #68719476736 r868 = ~r868;
  always #137438953472 r869 = ~r869;
  always #274877906944 r870 = ~r870;
  always #549755813888 r871 = ~r871;
  always #1099511627776 r872 = ~r872;
  always #2199023255552 r873 = ~r873;
  always #4398046511104 r874 = ~r874;
  always #8796093022208 r875 = ~r875;
  always #17592186044416 r876 = ~r876;
  always #35184372088832 r877 = ~r877;
  always #70368744177664 r878 = ~r878;
  always #140737488355328 r879 = ~r879;
  always #281474976710656 r880 = ~r880;
  always #562949953421312 r881 = ~r881;
  always #1125899906842624 r882 = ~r882;
  always #2251799813685248 r883 = ~r883;
  always #4503599627370496 r884 = ~r884;
  always #9007199254740992 r885 = ~r885;
  always #18014398509481984 r886 = ~r886;
  always #36028797018963968 r887 = ~r887;
  always #72057594037927936 r888 = ~r888;
  always #144115188075855872 r889 = ~r889;
  always #288230376151711744 r890 = ~r890;
  always #576460752303423488 r891 = ~r891;
  always #1152921504606846976 r892 = ~r892;
  always #2305843009213693952 r893 = ~r893;
  always #4611686018427387904 r894 = ~r894;
  always #9223372036854775808 r895 = ~r895;
  always #1 r896 = ~r896;
  always #2 r897 = ~r897;
  always #4 r898 = ~r898;
  always #8 r899 = ~r899;
  always #16 r900 = ~r900;
  always #32 r901 = ~r901;
  always #64 r902 = ~r902;
  always #128 r903 = ~r903;
  always #256 r904 = ~r904;
  always #512 r905 = ~r905;
  always #1024 r906 = ~r906;
  always #2048 r907 = ~r907;
  always #4096 r908 = ~r908;
  always #8192 r909 = ~r909;
  always #16384 r910 = ~r910;
  always #32768 r911 = ~r911;
  always #65536 r912 = ~r912;
  always #131072 r913 = ~r913;
  always #262144 r914 = ~r914;
  always #524288 r915 = ~r915;
  always #1048576 r916 = ~r916;
  always #2097152 r917 = ~r917;
  always #4194304 r918 = ~r918;
  always #8388608 r919 = ~r919;
  always #16777216 r920 = ~r920;
  always #33554432 r921 = ~r921;
  always #67108864 r922 = ~r922;
  always #134217728 r923 = ~r923;
  always #268435456 r924 = ~r924;
  always #536870912 r925 = ~r925;
  always #1073741824 r926 = ~r926;
  always #2147483648 r927 = ~r927;
  always #4294967296 r928 = ~r928;
  always #8589934592 r929 = ~r929;
  always #17179869184 r930 = ~r930;
  always #34359738368 r931 = ~r931;
  always #68719476736 r932 = ~r932;
  always #137438953472 r933 = ~r933;
  always #274877906944 r934 = ~r934;
  always #549755813888 r935 = ~r935;
  always #1099511627776 r936 = ~r936;
  always #2199023255552 r937 = ~r937;
  always #4398046511104 r938 = ~r938;
  always #8796093022208 r939 = ~r939;
  always #17592186044416 r940 = ~r940;
  always #35184372088832 r941 = ~r941;
  always #70368744177664 r942 = ~r942;
  always #140737488355328 r943 = ~r943;
  always #281474976710656 r944 = ~r944;
  always #562949953421312 r945 = ~r945;
  always #1125899906842624 r946 = ~r946;
  always #2251799813685248 r947 = ~r947;
  always #4503599627370496 r948 = ~r948;
  always #9007199254740992 r949 = ~r949;
  always #18014398509481984 r950 = ~r950;
  always #36028797018963968 r951 = ~r951;
  always #72057594037927936 r952 = ~r952;
  always #144115188075855872 r953 = ~r953;
  always #288230376151711744 r954 = ~r954;
  always #576460752303423488 r955 = ~r955;
  always #1152921504606846976 r956 = ~r956;
  always #2305843009213693952 r957 = ~r957;
  always #4611686018427387904 r958 = ~r958;
  always #9223372036854775808 r959 = ~r959;
  always #1 r960 = ~r960;
  always #2 r961 = ~r961;
  always #4 r962 = ~r962;
  always #8 r963 = ~r963;
  always #16 r964 = ~r964;
  always #32 r965 = ~r965;
  always #64 r966 = ~r966;
  always #128 r967 = ~r967;
  always #256 r968 = ~r968;
  always #512 r969 = ~r969;
  always #1024 r970 = ~r970;
  always #2048 r971 = ~r971;
  always #4096 r972 = ~r972;
  always #8192 r973 = ~r973;
  always #16384 r974 = ~r974;
  always #32768 r975 = ~r975;
  always #65536 r976 = ~r976;
  always #131072 r977 = ~r977;
  always #262144 r978 = ~r978;
  always #524288 r979 = ~r979;
  always #1048576 r980 = ~r980;
  always #2097152 r981 = ~r981;
  always #4194304 r982 = ~r982;
  always #8388608 r983 = ~r983;
  always #16777216 r984 = ~r984;
  always #33554432 r985 = ~r985;
  always #67108864 r986 = ~r986;
  always #134217728 r987 = ~r987;
  always #268435456 r988 = ~r988;
  always #536870912 r989 = ~r989;
  always #1073741824 r990 = ~r990;
  always #2147483648 r991 = ~r991;
  always #4294967296 r992 = ~r992;
  always #8589934592 r993 = ~r993;
  always #17179869184 r994 = ~r994;
  always #34359738368 r995 = ~r995;
  always #68719476736 r996 = ~r996;
  always #137438953472 r997 = ~r997;
  always #274877906944 r998 = ~r998;
  always #549755813888 r999 = ~r999;
endmodule
*/
// ****** TestBench Module Defination End ******

/*
// ******* The results for this case *********
******* result_1.txt *********
1)
  Loop Signals: w_894_262, w_894_263, w_894_264, w_894_265, w_894_266, w_894_267, w_894_268, w_894_269, w_894_270, w_894_271, w_894_272, w_894_273, 
  Loop Gates: I894_261.port1, I894_262.port1, I894_263.port2, I894_264.port1, I894_265.port2, I894_266.port1, I894_267.port1, I894_268.port1, I894_269.port1, I894_270.port1, I894_271.port2, I894_272.port1, 

2)
  Loop Signals: w_894_270, w_894_277, w_894_278, w_894_279, w_894_280, w_894_281, w_894_282, w_894_283, w_894_284, w_894_285, w_894_287, 
  Loop Gates: I894_268.port2, I894_273.port1, I894_274.port1, I894_275.port1, I894_276.port1, I894_277.port1, I894_278.port2, I894_279.port2, I894_280.port2, I894_281.port1, I894_282.port2, 

3)
  Loop Signals: w_152_770, w_152_771, w_152_772, w_152_773, w_152_774, w_152_775, 
  Loop Gates: I152_769.port1, I152_770.port1, I152_771.port1, I152_772.port2, I152_773.port2, I152_774.port2, 

4)
  Loop Signals: w_152_770, w_152_779, w_152_780, w_152_781, w_152_782, w_152_783, w_152_784, w_152_786, 
  Loop Gates: I152_774.port1, I152_775.port1, I152_776.port2, I152_777.port1, I152_778.port1, I152_779.port2, I152_780.port1, I152_781.port2, 

5)
  Loop Signals: w_156_708, w_156_709, w_156_710, w_156_711, w_156_712, w_156_713, 
  Loop Gates: I156_707.port1, I156_708.port1, I156_709.port1, I156_710.port2, I156_711.port2, I156_712.port2, 

6)
  Loop Signals: w_450_116, w_450_117, w_450_118, w_450_119, w_450_120, w_450_121, w_450_122, w_450_123, 
  Loop Gates: I450_115.port2, I450_116.port1, I450_117.port1, I450_118.port1, I450_119.port2, I450_120.port2, I450_121.port1, I450_122.port1, 

7)
  Loop Signals: w_802_628, w_802_629, w_802_630, w_802_631, w_802_632, w_802_633, w_802_634, 
  Loop Gates: I802_627.port1, I802_628.port1, I802_629.port1, I802_630.port2, I802_631.port2, I802_632.port1, I802_633.port2, 

8)
  Loop Signals: w_474_430, w_474_431, w_474_432, w_474_433, w_474_434, 
  Loop Gates: I474_429.port2, I474_430.port1, I474_431.port1, I474_432.port2, I474_433.port2, 

9)
  Loop Signals: w_474_431, w_474_438, w_474_439, w_474_440, w_474_441, w_474_442, w_474_443, w_474_444, w_474_445, w_474_446, w_474_447, w_474_449, 
  Loop Gates: I474_429.port1, I474_434.port1, I474_435.port2, I474_436.port2, I474_437.port1, I474_438.port2, I474_439.port2, I474_440.port2, I474_441.port2, I474_442.port1, I474_443.port1, I474_444.port2, 

10)
  Loop Signals: w_847_002, w_847_003, w_847_004, w_847_005, w_847_006, 
  Loop Gates: I847_001.port2, I847_002.port2, I847_003.port1, I847_004.port2, I847_005.port1, 

11)
  Loop Signals: w_036_285, w_036_286, w_036_287, w_036_288, w_036_289, w_036_290, 
  Loop Gates: I036_284.port2, I036_285.port2, I036_286.port1, I036_287.port1, I036_288.port2, I036_289.port1, 

12)
  Loop Signals: w_737_555, w_737_556, w_737_557, w_737_558, w_737_559, w_737_560, w_737_561, 
  Loop Gates: I737_554.port1, I737_555.port2, I737_556.port1, I737_557.port2, I737_558.port2, I737_559.port1, I737_560.port1, 

13)
  Loop Signals: w_713_133, w_713_134, w_713_135, 
  Loop Gates: I713_132.port2, I713_133.port1, I713_134.port1, 

14)
  Loop Signals: w_713_134, w_713_139, w_713_140, w_713_141, w_713_142, w_713_143, w_713_144, w_713_145, w_713_146, w_713_147, w_713_148, w_713_149, w_713_151, 
  Loop Gates: I713_132.port1, I713_135.port1, I713_136.port1, I713_137.port1, I713_138.port1, I713_139.port2, I713_140.port2, I713_141.port1, I713_142.port2, I713_143.port1, I713_144.port2, I713_145.port1, I713_146.port2, 

15)
  Loop Signals: w_971_280, w_971_281, w_971_282, w_971_283, w_971_284, w_971_285, w_971_286, w_971_287, w_971_288, 
  Loop Gates: I971_279.port1, I971_280.port2, I971_281.port1, I971_282.port1, I971_283.port2, I971_284.port1, I971_285.port2, I971_286.port1, I971_287.port1, 

16)
  Loop Signals: w_318_063, w_318_064, w_318_065, w_318_066, w_318_067, w_318_068, w_318_069, w_318_070, w_318_071, w_318_072, 
  Loop Gates: I318_062.port1, I318_063.port1, I318_064.port2, I318_065.port1, I318_066.port1, I318_067.port2, I318_068.port2, I318_069.port1, I318_070.port1, I318_071.port1, 

17)
  Loop Signals: w_483_216, w_483_217, w_483_218, w_483_219, w_483_220, w_483_221, w_483_222, w_483_223, w_483_224, w_483_225, w_483_226, w_483_227, 
  Loop Gates: I483_215.port2, I483_216.port1, I483_217.port1, I483_218.port2, I483_219.port2, I483_220.port2, I483_221.port1, I483_222.port2, I483_223.port1, I483_224.port1, I483_225.port1, I483_226.port2, 

18)
  Loop Signals: w_935_969, w_935_970, w_935_971, w_935_972, w_935_973, 
  Loop Gates: I935_968.port2, I935_969.port1, I935_970.port2, I935_971.port2, I935_972.port1, 

19)
  Loop Signals: w_935_969, w_935_977, w_935_978, w_935_979, w_935_981, 
  Loop Gates: I935_972.port2, I935_973.port2, I935_974.port2, I935_975.port1, I935_976.port2, 

20)
  Loop Signals: w_188_535, w_188_536, w_188_537, w_188_538, w_188_539, 
  Loop Gates: I188_534.port1, I188_535.port2, I188_536.port2, I188_537.port1, I188_538.port2, 

21)
  Loop Signals: w_188_535, w_188_543, w_188_544, w_188_545, w_188_546, w_188_547, w_188_548, w_188_550, 
  Loop Gates: I188_538.port1, I188_539.port1, I188_540.port1, I188_541.port1, I188_542.port2, I188_543.port1, I188_544.port1, I188_545.port2, 

22)
  Loop Signals: w_240_814, w_240_815, w_240_816, w_240_817, w_240_818, w_240_819, w_240_820, w_240_821, 
  Loop Gates: I240_813.port1, I240_814.port1, I240_815.port2, I240_816.port2, I240_817.port2, I240_818.port2, I240_819.port1, I240_820.port1, 

23)
  Loop Signals: w_955_348, w_955_349, w_955_350, w_955_351, w_955_352, w_955_353, w_955_354, w_955_355, w_955_356, w_955_357, 
  Loop Gates: I955_347.port1, I955_348.port2, I955_349.port2, I955_350.port1, I955_351.port2, I955_352.port2, I955_353.port1, I955_354.port1, I955_355.port2, I955_356.port2, 

24)
  Loop Signals: w_905_810, w_905_811, w_905_812, 
  Loop Gates: I905_809.port1, I905_810.port2, I905_811.port1, 

25)
  Loop Signals: w_905_812, w_905_816, w_905_817, w_905_818, w_905_819, w_905_820, w_905_821, w_905_823, 
  Loop Gates: I905_810.port1, I905_812.port2, I905_813.port1, I905_814.port1, I905_815.port2, I905_816.port2, I905_817.port1, I905_818.port2, 

26)
  Loop Signals: w_968_916, w_968_917, w_968_918, w_968_919, w_968_920, w_968_921, w_968_922, w_968_923, w_968_924, w_968_925, w_968_926, w_968_927, 
  Loop Gates: I968_915.port2, I968_916.port1, I968_917.port1, I968_918.port1, I968_919.port2, I968_920.port2, I968_921.port1, I968_922.port1, I968_923.port2, I968_924.port1, I968_925.port1, I968_926.port1, 

27)
  Loop Signals: w_968_917, w_968_931, w_968_932, w_968_933, w_968_934, w_968_936, 
  Loop Gates: I968_915.port1, I968_927.port2, I968_928.port2, I968_929.port2, I968_930.port1, I968_931.port2, 

28)
  Loop Signals: w_035_651, w_035_652, w_035_653, w_035_654, w_035_655, w_035_656, w_035_657, w_035_658, w_035_659, w_035_660, 
  Loop Gates: I035_650.port1, I035_651.port2, I035_652.port1, I035_653.port2, I035_654.port1, I035_655.port2, I035_656.port1, I035_657.port1, I035_658.port2, I035_659.port2, 

29)
  Loop Signals: w_899_531, w_899_532, w_899_533, w_899_534, w_899_535, w_899_536, w_899_537, w_899_538, w_899_539, w_899_540, 
  Loop Gates: I899_530.port1, I899_531.port2, I899_532.port2, I899_533.port2, I899_534.port2, I899_535.port1, I899_536.port2, I899_537.port1, I899_538.port2, I899_539.port1, 

30)
  Loop Signals: w_416_776, w_416_777, w_416_778, w_416_779, w_416_780, w_416_781, 
  Loop Gates: I416_775.port1, I416_776.port2, I416_777.port2, I416_778.port1, I416_779.port2, I416_780.port1, 

31)
  Loop Signals: w_096_628, w_096_629, w_096_630, w_096_631, w_096_632, w_096_633, w_096_634, w_096_635, w_096_636, w_096_637, w_096_638, 
  Loop Gates: I096_627.port2, I096_628.port1, I096_629.port1, I096_630.port1, I096_631.port2, I096_632.port2, I096_633.port1, I096_634.port2, I096_635.port2, I096_636.port1, I096_637.port1, 

32)
  Loop Signals: w_096_631, w_096_642, w_096_643, w_096_644, w_096_645, w_096_646, w_096_647, w_096_648, w_096_649, w_096_650, w_096_651, w_096_653, 
  Loop Gates: I096_629.port2, I096_638.port1, I096_639.port1, I096_640.port2, I096_641.port2, I096_642.port1, I096_643.port1, I096_644.port1, I096_645.port1, I096_646.port2, I096_647.port1, I096_648.port2, 

33)
  Loop Signals: w_143_576, w_143_577, w_143_578, 
  Loop Gates: I143_575.port1, I143_576.port1, I143_577.port2, 

34)
  Loop Signals: w_316_852, w_316_853, w_316_854, w_316_855, w_316_856, w_316_857, w_316_858, w_316_859, w_316_860, w_316_861, w_316_862, 
  Loop Gates: I316_851.port2, I316_852.port1, I316_853.port1, I316_854.port1, I316_855.port1, I316_856.port1, I316_857.port1, I316_858.port1, I316_859.port1, I316_860.port1, I316_861.port2, 

35)
  Loop Signals: w_743_142, w_743_143, w_743_144, w_743_145, w_743_146, 
  Loop Gates: I743_141.port1, I743_142.port1, I743_143.port2, I743_144.port1, I743_145.port2, 

36)
  Loop Signals: w_719_615, w_719_616, w_719_617, w_719_618, w_719_619, w_719_620, w_719_621, w_719_622, w_719_623, 
  Loop Gates: I719_614.port2, I719_615.port1, I719_616.port1, I719_617.port1, I719_618.port1, I719_619.port2, I719_620.port2, I719_621.port1, I719_622.port2, 

37)
  Loop Signals: w_503_730, w_503_731, w_503_732, w_503_733, w_503_734, w_503_735, w_503_736, w_503_737, w_503_738, w_503_739, 
  Loop Gates: I503_729.port1, I503_730.port1, I503_731.port1, I503_732.port2, I503_733.port2, I503_734.port2, I503_735.port1, I503_736.port1, I503_737.port2, I503_738.port2, 

38)
  Loop Signals: w_503_739, w_503_743, w_503_744, w_503_745, w_503_746, w_503_747, w_503_748, w_503_749, w_503_750, w_503_751, w_503_752, w_503_754, 
  Loop Gates: I503_737.port1, I503_739.port1, I503_740.port2, I503_741.port1, I503_742.port2, I503_743.port2, I503_744.port2, I503_745.port1, I503_746.port1, I503_747.port1, I503_748.port1, I503_749.port2, 

39)
  Loop Signals: w_703_395, w_703_396, w_703_397, w_703_398, w_703_399, w_703_400, w_703_401, w_703_402, w_703_403, w_703_404, w_703_405, w_703_406, 
  Loop Gates: I703_394.port1, I703_395.port1, I703_396.port1, I703_397.port2, I703_398.port2, I703_399.port1, I703_400.port1, I703_401.port1, I703_402.port1, I703_403.port2, I703_404.port2, I703_405.port1, 

40)
  Loop Signals: w_292_705, w_292_706, w_292_707, w_292_708, w_292_709, w_292_710, w_292_711, w_292_712, w_292_713, w_292_714, 
  Loop Gates: I292_704.port2, I292_705.port2, I292_706.port1, I292_707.port1, I292_708.port1, I292_709.port1, I292_710.port1, I292_711.port2, I292_712.port1, I292_713.port1, 

41)
  Loop Signals: w_896_755, w_896_756, w_896_757, w_896_758, 
  Loop Gates: I896_754.port1, I896_755.port1, I896_756.port1, I896_757.port2, 

42)
  Loop Signals: w_878_748, w_878_749, w_878_750, w_878_751, w_878_752, w_878_753, w_878_754, w_878_755, 
  Loop Gates: I878_747.port1, I878_748.port1, I878_749.port2, I878_750.port1, I878_751.port2, I878_752.port1, I878_753.port2, I878_754.port2, 

43)
  Loop Signals: w_878_754, w_878_759, w_878_760, w_878_761, w_878_762, w_878_763, w_878_764, w_878_766, 
  Loop Gates: I878_752.port2, I878_755.port1, I878_756.port1, I878_757.port2, I878_758.port1, I878_759.port1, I878_760.port1, I878_761.port2, 

44)
  Loop Signals: w_400_790, w_400_791, w_400_792, w_400_793, w_400_794, w_400_795, w_400_796, w_400_797, w_400_798, 
  Loop Gates: I400_789.port2, I400_790.port1, I400_791.port1, I400_792.port1, I400_793.port2, I400_794.port2, I400_795.port1, I400_796.port1, I400_797.port1, 

45)
  Loop Signals: w_597_329, w_597_330, w_597_331, w_597_332, w_597_333, w_597_334, w_597_335, w_597_336, w_597_337, 
  Loop Gates: I597_328.port1, I597_329.port1, I597_330.port1, I597_331.port2, I597_332.port1, I597_333.port1, I597_334.port2, I597_335.port2, I597_336.port1, 

46)
  Loop Signals: w_597_330, w_597_341, w_597_342, w_597_343, w_597_344, w_597_345, w_597_346, w_597_347, w_597_348, w_597_349, w_597_351, 
  Loop Gates: I597_328.port2, I597_337.port1, I597_338.port2, I597_339.port1, I597_340.port1, I597_341.port2, I597_342.port2, I597_343.port1, I597_344.port1, I597_345.port1, I597_346.port2, 

47)
  Loop Signals: w_788_201, w_788_202, w_788_203, w_788_204, w_788_205, 
  Loop Gates: I788_200.port1, I788_201.port2, I788_202.port1, I788_203.port2, I788_204.port2, 

48)
  Loop Signals: w_788_204, w_788_209, w_788_210, w_788_211, w_788_212, w_788_213, w_788_214, w_788_215, w_788_216, w_788_217, w_788_219, 
  Loop Gates: I788_202.port2, I788_205.port2, I788_206.port1, I788_207.port2, I788_208.port1, I788_209.port2, I788_210.port2, I788_211.port1, I788_212.port1, I788_213.port1, I788_214.port2, 

49)
  Loop Signals: w_822_988, w_822_989, w_822_990, 
  Loop Gates: I822_987.port1, I822_988.port2, I822_989.port1, 

50)
  Loop Signals: w_720_811, w_720_812, w_720_813, w_720_814, w_720_815, w_720_816, 
  Loop Gates: I720_811.port1, I720_812.port1, I720_813.port1, I720_814.port1, I720_815.port2, I720_816.port1, 

******* result_2.txt *********
1)
  Loop Signals: w_894_262, w_894_263, w_894_264, w_894_265, w_894_266, w_894_267, w_894_268, w_894_269, w_894_270, w_894_271, w_894_272, w_894_273, 
  Loop Gates: I894_261.port1, I894_262.port1, I894_263.port2, I894_264.port1, I894_265.port2, I894_266.port1, I894_267.port1, I894_268.port1, I894_269.port1, I894_270.port1, I894_271.port2, I894_272.port1, 

2)
  Loop Signals: w_152_770, w_152_771, w_152_772, w_152_773, w_152_774, w_152_775, 
  Loop Gates: I152_769.port1, I152_770.port1, I152_771.port1, I152_772.port2, I152_773.port2, I152_774.port2, 

3)
  Loop Signals: w_152_770, w_152_779, w_152_780, w_152_781, w_152_782, w_152_783, w_152_784, w_152_786, 
  Loop Gates: I152_774.port1, I152_775.port1, I152_776.port2, I152_777.port1, I152_778.port1, I152_779.port2, I152_780.port1, I152_781.port2, 

4)
  Loop Signals: w_156_708, w_156_709, w_156_710, w_156_711, w_156_712, w_156_713, 
  Loop Gates: I156_707.port1, I156_708.port1, I156_709.port1, I156_710.port2, I156_711.port2, I156_712.port2, 

5)
  Loop Signals: w_474_431, w_474_438, w_474_439, w_474_440, w_474_441, w_474_442, w_474_443, w_474_444, w_474_445, w_474_446, w_474_447, w_474_449, 
  Loop Gates: I474_429.port1, I474_434.port1, I474_435.port2, I474_436.port2, I474_437.port1, I474_438.port2, I474_439.port2, I474_440.port2, I474_441.port2, I474_442.port1, I474_443.port1, I474_444.port2, 

6)
  Loop Signals: w_737_555, w_737_556, w_737_557, w_737_558, w_737_559, w_737_560, w_737_561, 
  Loop Gates: I737_554.port1, I737_555.port2, I737_556.port1, I737_557.port2, I737_558.port2, I737_559.port1, I737_560.port1, 

7)
  Loop Signals: w_713_134, w_713_139, w_713_140, w_713_141, w_713_142, w_713_143, w_713_144, w_713_145, w_713_146, w_713_147, w_713_148, w_713_149, w_713_151, 
  Loop Gates: I713_132.port1, I713_135.port1, I713_136.port1, I713_137.port1, I713_138.port1, I713_139.port2, I713_140.port2, I713_141.port1, I713_142.port2, I713_143.port1, I713_144.port2, I713_145.port1, I713_146.port2, 

8)
  Loop Signals: w_971_280, w_971_281, w_971_282, w_971_283, w_971_284, w_971_285, w_971_286, w_971_287, w_971_288, 
  Loop Gates: I971_279.port1, I971_280.port2, I971_281.port1, I971_282.port1, I971_283.port2, I971_284.port1, I971_285.port2, I971_286.port1, I971_287.port1, 

9)
  Loop Signals: w_935_969, w_935_977, w_935_978, w_935_979, w_935_981, 
  Loop Gates: I935_972.port2, I935_973.port2, I935_974.port2, I935_975.port1, I935_976.port2, 

10)
  Loop Signals: w_188_535, w_188_536, w_188_537, w_188_538, w_188_539, 
  Loop Gates: I188_534.port1, I188_535.port2, I188_536.port2, I188_537.port1, I188_538.port2, 

11)
  Loop Signals: w_188_535, w_188_543, w_188_544, w_188_545, w_188_546, w_188_547, w_188_548, w_188_550, 
  Loop Gates: I188_538.port1, I188_539.port1, I188_540.port1, I188_541.port1, I188_542.port2, I188_543.port1, I188_544.port1, I188_545.port2, 

12)
  Loop Signals: w_240_814, w_240_815, w_240_816, w_240_817, w_240_818, w_240_819, w_240_820, w_240_821, 
  Loop Gates: I240_813.port1, I240_814.port1, I240_815.port2, I240_816.port2, I240_817.port2, I240_818.port2, I240_819.port1, I240_820.port1, 

13)
  Loop Signals: w_905_810, w_905_811, w_905_812, 
  Loop Gates: I905_809.port1, I905_810.port2, I905_811.port1, 

14)
  Loop Signals: w_899_531, w_899_532, w_899_533, w_899_534, w_899_535, w_899_536, w_899_537, w_899_538, w_899_539, w_899_540, 
  Loop Gates: I899_530.port1, I899_531.port2, I899_532.port2, I899_533.port2, I899_534.port2, I899_535.port1, I899_536.port2, I899_537.port1, I899_538.port2, I899_539.port1, 

15)
  Loop Signals: w_416_776, w_416_777, w_416_778, w_416_779, w_416_780, w_416_781, 
  Loop Gates: I416_775.port1, I416_776.port2, I416_777.port2, I416_778.port1, I416_779.port2, I416_780.port1, 

16)
  Loop Signals: w_143_576, w_143_577, w_143_578, 
  Loop Gates: I143_575.port1, I143_576.port1, I143_577.port2, 

17)
  Loop Signals: w_719_615, w_719_616, w_719_617, w_719_618, w_719_619, w_719_620, w_719_621, w_719_622, w_719_623, 
  Loop Gates: I719_614.port2, I719_615.port1, I719_616.port1, I719_617.port1, I719_618.port1, I719_619.port2, I719_620.port2, I719_621.port1, I719_622.port2, 

18)
  Loop Signals: w_292_705, w_292_706, w_292_707, w_292_708, w_292_709, w_292_710, w_292_711, w_292_712, w_292_713, w_292_714, 
  Loop Gates: I292_704.port2, I292_705.port2, I292_706.port1, I292_707.port1, I292_708.port1, I292_709.port1, I292_710.port1, I292_711.port2, I292_712.port1, I292_713.port1, 

19)
  Loop Signals: w_400_790, w_400_791, w_400_792, w_400_793, w_400_794, w_400_795, w_400_796, w_400_797, w_400_798, 
  Loop Gates: I400_789.port2, I400_790.port1, I400_791.port1, I400_792.port1, I400_793.port2, I400_794.port2, I400_795.port1, I400_796.port1, I400_797.port1, 

20)
  Loop Signals: w_597_330, w_597_341, w_597_342, w_597_343, w_597_344, w_597_345, w_597_346, w_597_347, w_597_348, w_597_349, w_597_351, 
  Loop Gates: I597_328.port2, I597_337.port1, I597_338.port2, I597_339.port1, I597_340.port1, I597_341.port2, I597_342.port2, I597_343.port1, I597_344.port1, I597_345.port1, I597_346.port2, 

21)
  Loop Signals: w_822_988, w_822_989, w_822_990, 
  Loop Gates: I822_987.port1, I822_988.port2, I822_989.port1, 

22)
  Loop Signals: w_720_811, w_720_812, w_720_813, w_720_814, w_720_815, w_720_816, 
  Loop Gates: I720_811.port1, I720_812.port1, I720_813.port1, I720_814.port1, I720_815.port2, I720_816.port1, 

******* result_3.txt *********
1)
  Loop Signals: w_894_270, w_894_277, w_894_278, w_894_279, w_894_280, w_894_281, w_894_282, w_894_283, w_894_284, w_894_285, w_894_287, 
  Loop Gates: I894_268.port2, I894_273.port1, I894_274.port1, I894_275.port1, I894_276.port1, I894_277.port1, I894_278.port2, I894_279.port2, I894_280.port2, I894_281.port1, I894_282.port2, 
  Loop Conditions: I894_268.port2=1, I894_274.port2=1, I894_277.port2=0, I894_278.port1=0, I894_279.port1=0, I894_280.port1=1, I894_282.port2=1, 
  (Signal Values: w_068_024=0, w_095_040=0, w_280_023=1, w_449_078=0, w_511_108=1, w_894_285=1, w_894_287=1, )

2)
  Loop Signals: w_450_116, w_450_117, w_450_118, w_450_119, w_450_120, w_450_121, w_450_122, w_450_123, 
  Loop Gates: I450_115.port2, I450_116.port1, I450_117.port1, I450_118.port1, I450_119.port2, I450_120.port2, I450_121.port1, I450_122.port1, 
  Loop Conditions: I450_115.port1=1, I450_116.port2=1, I450_119.port1=0, I450_120.port1=1, I450_121.port2=1, I450_122.port2=1, 
  (Signal Values: w_158_546=1, w_183_110=0, w_246_274=1, w_369_081=1, w_373_024=1, w_389_092=1, )

3)
  Loop Signals: w_802_628, w_802_629, w_802_630, w_802_631, w_802_632, w_802_633, w_802_634, 
  Loop Gates: I802_627.port1, I802_628.port1, I802_629.port1, I802_630.port2, I802_631.port2, I802_632.port1, I802_633.port2, 
  Loop Conditions: I802_628.port2=1, I802_629.port2=1, I802_630.port1=1, I802_631.port1=1, I802_632.port2=1, I802_633.port1=1, 
  (Signal Values: w_042_065=1, w_256_124=1, w_344_001=1, w_402_188=1, w_423_151=1, w_564_518=1, )

4)
  Loop Signals: w_474_430, w_474_431, w_474_432, w_474_433, w_474_434, 
  Loop Gates: I474_429.port2, I474_430.port1, I474_431.port1, I474_432.port2, I474_433.port2, 
  Loop Conditions: I474_429.port2=1, I474_430.port2=1, I474_431.port2=1, I474_432.port1=1, I474_433.port1=0, 
  (Signal Values: w_133_416=0, w_283_373=1, w_325_265=1, w_344_000=1, w_474_430=1, )

5)
  Loop Signals: w_847_002, w_847_003, w_847_004, w_847_005, w_847_006, 
  Loop Gates: I847_001.port2, I847_002.port2, I847_003.port1, I847_004.port2, I847_005.port1, 
  Loop Conditions: I847_001.port1=1, I847_002.port1=1, I847_003.port2=1, I847_004.port1=1, I847_005.port2=1, 
  (Signal Values: w_004_033=1, w_076_422=1, w_197_778=1, w_202_012=1, w_826_130=1, )

6)
  Loop Signals: w_036_285, w_036_286, w_036_287, w_036_288, w_036_289, w_036_290, 
  Loop Gates: I036_284.port2, I036_285.port2, I036_286.port1, I036_287.port1, I036_288.port2, I036_289.port1, 
  Loop Conditions: I036_284.port1=1, I036_285.port1=1, I036_286.port2=1, I036_287.port2=1, I036_288.port1=0, I036_289.port2=1, 
  (Signal Values: w_001_264=1, w_004_009=1, w_016_370=0, w_026_361=1, w_028_281=1, w_035_274=1, )

7)
  Loop Signals: w_713_133, w_713_134, w_713_135, 
  Loop Gates: I713_132.port2, I713_133.port1, I713_134.port1, 
  Loop Conditions: I713_132.port2=1, I713_134.port2=0, 
  (Signal Values: w_578_266=0, w_713_133=1, )

8)
  Loop Signals: w_318_063, w_318_064, w_318_065, w_318_066, w_318_067, w_318_068, w_318_069, w_318_070, w_318_071, w_318_072, 
  Loop Gates: I318_062.port1, I318_063.port1, I318_064.port2, I318_065.port1, I318_066.port1, I318_067.port2, I318_068.port2, I318_069.port1, I318_070.port1, I318_071.port1, 
  Loop Conditions: I318_062.port2=0, I318_064.port1=1, I318_067.port1=1, I318_068.port1=1, I318_069.port2=1, 
  (Signal Values: w_004_009=1, w_026_387=1, w_119_119=1, w_138_183=1, w_260_510=0, )

9)
  Loop Signals: w_483_216, w_483_217, w_483_218, w_483_219, w_483_220, w_483_221, w_483_222, w_483_223, w_483_224, w_483_225, w_483_226, w_483_227, 
  Loop Gates: I483_215.port2, I483_216.port1, I483_217.port1, I483_218.port2, I483_219.port2, I483_220.port2, I483_221.port1, I483_222.port2, I483_223.port1, I483_224.port1, I483_225.port1, I483_226.port2, 
  Loop Conditions: I483_215.port1=0, I483_216.port2=0, I483_217.port2=1, I483_218.port1=1, I483_219.port1=0, I483_220.port1=1, I483_221.port2=1, I483_222.port1=1, I483_223.port2=0, I483_224.port2=1, I483_225.port2=1, I483_226.port1=1, 
  (Signal Values: w_019_353=1, w_034_113=0, w_053_404=1, w_137_579=0, w_146_106=1, w_223_023=1, w_260_812=0, w_269_031=1, w_270_103=1, w_293_625=1, w_442_003=0, w_444_007=1, )

10)
  Loop Signals: w_935_969, w_935_970, w_935_971, w_935_972, w_935_973, 
  Loop Gates: I935_968.port2, I935_969.port1, I935_970.port2, I935_971.port2, I935_972.port1, 
  Loop Conditions: I935_968.port1=1, I935_969.port2=1, I935_970.port1=1, I935_971.port1=1, I935_972.port2=0, 
  (Signal Values: w_498_527=1, w_567_775=1, w_610_178=1, w_804_005=1, w_935_981=0, )

11)
  Loop Signals: w_955_348, w_955_349, w_955_350, w_955_351, w_955_352, w_955_353, w_955_354, w_955_355, w_955_356, w_955_357, 
  Loop Gates: I955_347.port1, I955_348.port2, I955_349.port2, I955_350.port1, I955_351.port2, I955_352.port2, I955_353.port1, I955_354.port1, I955_355.port2, I955_356.port2, 
  Loop Conditions: I955_347.port2=1, I955_348.port1=1, I955_349.port1=0, I955_351.port1=1, I955_352.port1=1, I955_355.port1=1, I955_356.port1=0, 
  (Signal Values: w_132_166=1, w_287_109=1, w_289_855=1, w_450_081=0, w_509_040=0, w_628_163=1, w_689_291=1, )

12)
  Loop Signals: w_905_812, w_905_816, w_905_817, w_905_818, w_905_819, w_905_820, w_905_821, w_905_823, 
  Loop Gates: I905_810.port1, I905_812.port2, I905_813.port1, I905_814.port1, I905_815.port2, I905_816.port2, I905_817.port1, I905_818.port2, 
  Loop Conditions: I905_810.port2=1, I905_812.port1=1, I905_813.port2=1, I905_814.port2=0, I905_815.port1=1, I905_816.port1=1, I905_818.port2=1, 
  (Signal Values: w_156_622=1, w_205_113=0, w_377_284=1, w_721_271=1, w_842_229=1, w_905_811=1, w_905_821=1, )

13)
  Loop Signals: w_968_916, w_968_917, w_968_918, w_968_919, w_968_920, w_968_921, w_968_922, w_968_923, w_968_924, w_968_925, w_968_926, w_968_927, 
  Loop Gates: I968_915.port2, I968_916.port1, I968_917.port1, I968_918.port1, I968_919.port2, I968_920.port2, I968_921.port1, I968_922.port1, I968_923.port2, I968_924.port1, I968_925.port1, I968_926.port1, 
  Loop Conditions: I968_915.port2=1, I968_916.port2=0, I968_918.port2=1, I968_919.port1=0, I968_920.port1=1, I968_921.port2=0, I968_922.port2=0, I968_923.port1=1, 
  (Signal Values: w_076_142=1, w_097_495=0, w_146_314=1, w_238_080=1, w_280_016=0, w_560_550=0, w_691_066=0, w_968_916=1, )

14)
  Loop Signals: w_968_917, w_968_931, w_968_932, w_968_933, w_968_934, w_968_936, 
  Loop Gates: I968_915.port1, I968_927.port2, I968_928.port2, I968_929.port2, I968_930.port1, I968_931.port2, 
  Loop Conditions: I968_915.port2=1, I968_927.port1=1, I968_928.port1=1, I968_929.port1=1, I968_931.port2=1, 
  (Signal Values: w_292_413=1, w_556_244=1, w_644_363=1, w_968_916=1, w_968_934=1, )

15)
  Loop Signals: w_035_651, w_035_652, w_035_653, w_035_654, w_035_655, w_035_656, w_035_657, w_035_658, w_035_659, w_035_660, 
  Loop Gates: I035_650.port1, I035_651.port2, I035_652.port1, I035_653.port2, I035_654.port1, I035_655.port2, I035_656.port1, I035_657.port1, I035_658.port2, I035_659.port2, 
  Loop Conditions: I035_651.port1=0, I035_652.port2=1, I035_653.port1=1, I035_654.port2=1, I035_655.port1=1, I035_656.port2=1, I035_658.port1=1, I035_659.port1=0, 
  (Signal Values: w_001_666=1, w_002_110=1, w_007_437=0, w_008_613=0, w_008_746=1, w_016_370=1, w_017_002=1, w_030_166=1, )

16)
  Loop Signals: w_096_628, w_096_629, w_096_630, w_096_631, w_096_632, w_096_633, w_096_634, w_096_635, w_096_636, w_096_637, w_096_638, 
  Loop Gates: I096_627.port2, I096_628.port1, I096_629.port1, I096_630.port1, I096_631.port2, I096_632.port2, I096_633.port1, I096_634.port2, I096_635.port2, I096_636.port1, I096_637.port1, 
  Loop Conditions: I096_627.port1=1, I096_628.port2=1, I096_629.port2=1, I096_630.port2=1, I096_631.port1=1, I096_632.port1=1, I096_633.port2=0, I096_634.port1=1, I096_635.port1=1, I096_637.port2=1, 
  (Signal Values: w_003_107=1, w_010_492=1, w_014_474=1, w_025_532=1, w_043_028=1, w_051_123=0, w_082_323=1, w_086_060=1, w_093_600=1, w_096_653=1, )

17)
  Loop Signals: w_096_631, w_096_642, w_096_643, w_096_644, w_096_645, w_096_646, w_096_647, w_096_648, w_096_649, w_096_650, w_096_651, w_096_653, 
  Loop Gates: I096_629.port2, I096_638.port1, I096_639.port1, I096_640.port2, I096_641.port2, I096_642.port1, I096_643.port1, I096_644.port1, I096_645.port1, I096_646.port2, I096_647.port1, I096_648.port2, 
  Loop Conditions: I096_629.port2=1, I096_638.port2=0, I096_640.port1=1, I096_641.port1=0, I096_643.port2=1, I096_644.port2=1, I096_646.port1=1, I096_648.port2=1, 
  (Signal Values: w_005_259=0, w_017_011=1, w_020_013=0, w_026_309=1, w_046_539=1, w_075_189=1, w_096_651=1, w_096_653=1, )

18)
  Loop Signals: w_316_852, w_316_853, w_316_854, w_316_855, w_316_856, w_316_857, w_316_858, w_316_859, w_316_860, w_316_861, w_316_862, 
  Loop Gates: I316_851.port2, I316_852.port1, I316_853.port1, I316_854.port1, I316_855.port1, I316_856.port1, I316_857.port1, I316_858.port1, I316_859.port1, I316_860.port1, I316_861.port2, 
  Loop Conditions: I316_851.port1=1, I316_852.port2=1, I316_854.port2=0, I316_855.port2=0, I316_857.port2=1, I316_858.port2=1, I316_861.port1=1, 
  (Signal Values: w_049_250=0, w_060_242=1, w_117_290=1, w_145_091=0, w_158_198=1, w_191_036=1, w_314_388=1, )

19)
  Loop Signals: w_743_142, w_743_143, w_743_144, w_743_145, w_743_146, 
  Loop Gates: I743_141.port1, I743_142.port1, I743_143.port2, I743_144.port1, I743_145.port2, 
  Loop Conditions: I743_142.port2=0, I743_143.port1=1, I743_144.port2=0, I743_145.port1=0, 
  (Signal Values: w_138_690=0, w_143_279=1, w_430_279=0, w_510_377=0, )

20)
  Loop Signals: w_503_730, w_503_731, w_503_732, w_503_733, w_503_734, w_503_735, w_503_736, w_503_737, w_503_738, w_503_739, 
  Loop Gates: I503_729.port1, I503_730.port1, I503_731.port1, I503_732.port2, I503_733.port2, I503_734.port2, I503_735.port1, I503_736.port1, I503_737.port2, I503_738.port2, 
  Loop Conditions: I503_729.port2=1, I503_732.port1=0, I503_733.port1=0, I503_734.port1=0, I503_735.port2=0, I503_736.port2=1, I503_737.port2=0, I503_738.port1=1, 
  (Signal Values: w_025_146=0, w_097_329=0, w_133_177=0, w_257_044=1, w_406_437=1, w_410_093=0, w_497_072=1, w_503_738=0, )

21)
  Loop Signals: w_503_739, w_503_743, w_503_744, w_503_745, w_503_746, w_503_747, w_503_748, w_503_749, w_503_750, w_503_751, w_503_752, w_503_754, 
  Loop Gates: I503_737.port1, I503_739.port1, I503_740.port2, I503_741.port1, I503_742.port2, I503_743.port2, I503_744.port2, I503_745.port1, I503_746.port1, I503_747.port1, I503_748.port1, I503_749.port2, 
  Loop Conditions: I503_737.port2=0, I503_739.port2=1, I503_740.port1=1, I503_742.port1=1, I503_743.port1=1, I503_744.port1=1, I503_745.port2=1, I503_749.port2=1, 
  (Signal Values: w_059_272=1, w_099_070=1, w_107_072=1, w_381_632=1, w_394_118=1, w_493_023=1, w_503_738=0, w_503_752=1, )

22)
  Loop Signals: w_703_395, w_703_396, w_703_397, w_703_398, w_703_399, w_703_400, w_703_401, w_703_402, w_703_403, w_703_404, w_703_405, w_703_406, 
  Loop Gates: I703_394.port1, I703_395.port1, I703_396.port1, I703_397.port2, I703_398.port2, I703_399.port1, I703_400.port1, I703_401.port1, I703_402.port1, I703_403.port2, I703_404.port2, I703_405.port1, 
  Loop Conditions: I703_394.port2=1, I703_395.port2=1, I703_396.port2=0, I703_397.port1=1, I703_398.port1=1, I703_400.port2=1, I703_403.port1=1, I703_404.port1=1, I703_405.port2=1, 
  (Signal Values: w_058_128=1, w_091_002=1, w_169_034=1, w_428_765=1, w_480_285=1, w_500_173=1, w_518_369=1, w_611_013=0, w_686_000=1, )

23)
  Loop Signals: w_896_755, w_896_756, w_896_757, w_896_758, 
  Loop Gates: I896_754.port1, I896_755.port1, I896_756.port1, I896_757.port2, 
  Loop Conditions: I896_754.port2=1, I896_756.port2=1, I896_757.port1=1, 
  (Signal Values: w_149_392=1, w_182_210=1, w_300_036=1, )

24)
  Loop Signals: w_878_748, w_878_749, w_878_750, w_878_751, w_878_752, w_878_753, w_878_754, w_878_755, 
  Loop Gates: I878_747.port1, I878_748.port1, I878_749.port2, I878_750.port1, I878_751.port2, I878_752.port1, I878_753.port2, I878_754.port2, 
  Loop Conditions: I878_748.port2=0, I878_749.port1=1, I878_751.port1=1, I878_752.port2=0, I878_753.port1=0, I878_754.port1=1, 
  (Signal Values: w_033_352=1, w_451_379=1, w_520_251=1, w_539_036=0, w_635_153=0, w_878_766=0, )

25)
  Loop Signals: w_878_754, w_878_759, w_878_760, w_878_761, w_878_762, w_878_763, w_878_764, w_878_766, 
  Loop Gates: I878_752.port2, I878_755.port1, I878_756.port1, I878_757.port2, I878_758.port1, I878_759.port1, I878_760.port1, I878_761.port2, 
  Loop Conditions: I878_752.port2=0, I878_756.port2=1, I878_757.port1=1, I878_758.port2=1, I878_759.port2=0, I878_761.port2=1, 
  (Signal Values: w_155_027=0, w_396_533=1, w_527_041=1, w_658_148=1, w_878_764=1, w_878_766=0, )

26)
  Loop Signals: w_597_329, w_597_330, w_597_331, w_597_332, w_597_333, w_597_334, w_597_335, w_597_336, w_597_337, 
  Loop Gates: I597_328.port1, I597_329.port1, I597_330.port1, I597_331.port2, I597_332.port1, I597_333.port1, I597_334.port2, I597_335.port2, I597_336.port1, 
  Loop Conditions: I597_328.port2=0, I597_329.port2=1, I597_331.port1=1, I597_332.port2=0, I597_334.port1=0, I597_335.port1=0, I597_336.port2=1, 
  (Signal Values: w_003_003=0, w_227_199=0, w_362_019=1, w_435_090=1, w_468_004=0, w_543_064=1, w_597_351=0, )

27)
  Loop Signals: w_788_201, w_788_202, w_788_203, w_788_204, w_788_205, 
  Loop Gates: I788_200.port1, I788_201.port2, I788_202.port1, I788_203.port2, I788_204.port2, 
  Loop Conditions: I788_200.port2=0, I788_201.port1=0, I788_202.port2=0, I788_203.port1=1, I788_204.port1=1, 
  (Signal Values: w_357_147=0, w_705_598=1, w_706_150=1, w_751_361=0, w_788_219=0, )

28)
  Loop Signals: w_788_204, w_788_209, w_788_210, w_788_211, w_788_212, w_788_213, w_788_214, w_788_215, w_788_216, w_788_217, w_788_219, 
  Loop Gates: I788_202.port2, I788_205.port2, I788_206.port1, I788_207.port2, I788_208.port1, I788_209.port2, I788_210.port2, I788_211.port1, I788_212.port1, I788_213.port1, I788_214.port2, 
  Loop Conditions: I788_202.port2=0, I788_205.port1=1, I788_206.port2=1, I788_207.port1=1, I788_208.port2=1, I788_209.port1=1, I788_210.port1=0, I788_211.port2=1, I788_212.port2=0, I788_214.port2=1, 
  (Signal Values: w_066_210=1, w_125_190=1, w_138_191=1, w_194_453=1, w_209_171=0, w_730_090=1, w_759_380=0, w_764_052=1, w_788_217=1, w_788_219=0, )

******* result_4.txt *********
1)
  Loop Breaker: I894_268.port0-w_894_270-Register-w_894_270'-I894_281.port1 

2)
  Loop Breaker: I450_115.port0-w_450_117-Register-w_450_117'-I450_116.port1 

3)
  Loop Breaker: I802_627.port0-w_802_629-Register-w_802_629'-I802_628.port1 

4)
  Loop Breaker: I474_429.port0-w_474_431-Register-w_474_431'-I474_430.port1 

5)
  Loop Breaker: I847_001.port0-w_847_003-Register-w_847_003'-I847_002.port2 

6)
  Loop Breaker: I036_284.port0-w_036_286-Register-w_036_286'-I036_285.port2 

7)
  Loop Breaker: I713_132.port0-w_713_134-Register-w_713_134'-I713_133.port1 

8)
  Loop Breaker: I318_062.port0-w_318_064-Register-w_318_064'-I318_063.port1 

9)
  Loop Breaker: I483_215.port0-w_483_217-Register-w_483_217'-I483_216.port1 

10)
  Loop Breaker: I935_972.port0-w_935_969-Register-w_935_969'-I935_968.port2 

11)
  Loop Breaker: I955_347.port0-w_955_349-Register-w_955_349'-I955_348.port2 

12)
  Loop Breaker: I905_810.port0-w_905_812-Register-w_905_812'-I905_817.port1 

13)
  Loop Breaker: I968_915.port0-w_968_917-Register-w_968_917'-I968_916.port1 

14)
  Loop Breaker: I968_915.port0-w_968_917-Register-w_968_917'-I968_930.port1 

15)
  Loop Breaker: I035_650.port0-w_035_652-Register-w_035_652'-I035_651.port2 

16)
  Loop Breaker: I096_629.port0-w_096_631-Register-w_096_631'-I096_630.port1 

17)
  Loop Breaker: I096_629.port0-w_096_631-Register-w_096_631'-I096_647.port1 

18)
  Loop Breaker: I316_851.port0-w_316_853-Register-w_316_853'-I316_852.port1 

19)
  Loop Breaker: I743_141.port0-w_743_143-Register-w_743_143'-I743_142.port1 

20)
  Loop Breaker: I503_737.port0-w_503_739-Register-w_503_739'-I503_738.port2 

21)
  Loop Breaker: I503_737.port0-w_503_739-Register-w_503_739'-I503_748.port1 

22)
  Loop Breaker: I703_394.port0-w_703_396-Register-w_703_396'-I703_395.port1 

23)
  Loop Breaker: I896_754.port0-w_896_756-Register-w_896_756'-I896_755.port1 

24)
  Loop Breaker: I878_752.port0-w_878_754-Register-w_878_754'-I878_753.port2 

25)
  Loop Breaker: I878_752.port0-w_878_754-Register-w_878_754'-I878_760.port1 

26)
  Loop Breaker: I597_328.port0-w_597_330-Register-w_597_330'-I597_329.port1 

27)
  Loop Breaker: I788_202.port0-w_788_204-Register-w_788_204'-I788_203.port2 

28)
  Loop Breaker: I788_202.port0-w_788_204-Register-w_788_204'-I788_213.port1 

// ******* The results for this case End *********
*/

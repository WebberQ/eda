// Gate Level Verilog Code Generated!
// GateLvl:100 GateNum:100 GateInputNum:2
// ****** Basic Gate Module Defination ******
module or2(out, in1, in2);
  output out;
  input in1, in2;
  wire in1, in2, out;
  assign out = in1 || in2;
endmodule

module and2(out, in1, in2);
  output out;
  input in1, in2;
  wire in1, in2, out;
  assign out = in1 && in2;
endmodule

module not1(out, in);
  output out;
  input in;
  wire in,out;
  assign out = ~in;
endmodule

module nand2(out, in1, in2);
  output out;
  input in1, in2;
  wire in1, in2, out;
  assign out = ~(in1 && in2);
endmodule
// ****** Basic Gate Module Defination End ******

// ****** Combined Logic Module Defination ******
module combLogic( w_000_000, w_000_001, w_000_002, w_000_003, w_000_004, w_000_005, w_000_006, w_000_007, w_000_008, w_000_009, w_000_010, w_000_011, w_000_012, w_000_013, w_000_014, w_000_015, w_000_016, w_000_018, w_000_019, w_000_020, w_000_021, w_000_022, w_000_023, w_000_024, w_000_025, w_000_026, w_000_027, w_000_028, w_000_029, w_000_030, w_000_031, w_000_032, w_000_033, w_000_034, w_000_035, w_000_036, w_000_037, w_000_038, w_000_039, w_000_040, w_000_041, w_000_042, w_000_043, w_000_044, w_000_045, w_000_046, w_000_047, w_000_048, w_000_049, w_000_050, w_000_051, w_000_052, w_000_053, w_000_054, w_000_055, w_000_056, w_000_057, w_000_058, w_000_059, w_000_060, w_000_061, w_000_062, w_000_064, w_000_065, w_000_066, w_000_067, w_000_068, w_000_069, w_000_070, w_000_071, w_000_072, w_000_073, w_000_074, w_000_076, w_000_077, w_000_078, w_000_079, w_000_082, w_000_083, w_000_084, w_000_085, w_000_086, w_000_087, w_000_088, w_000_089, w_000_090, w_000_091, w_000_092, w_000_096, w_100_000, w_100_001, w_100_002, w_100_003, w_100_004, w_100_005, w_100_006, w_100_007, w_100_008, w_100_009, w_100_010, w_100_011, w_100_012, w_100_013, w_100_014, w_100_015, w_100_016, w_100_017, w_100_018, w_100_019, w_100_020, w_100_021, w_100_022, w_100_023, w_100_024, w_100_025, w_100_026, w_100_027, w_100_028, w_100_029, w_100_030, w_100_031, w_100_032, w_100_033, w_100_034, w_100_035, w_100_036, w_100_037, w_100_038, w_100_039 );
  inout w_000_000, w_000_001, w_000_002, w_000_003, w_000_004, w_000_005, w_000_006, w_000_007, w_000_008, w_000_009, w_000_010, w_000_011, w_000_012, w_000_013, w_000_014, w_000_015, w_000_016, w_000_018, w_000_019, w_000_020, w_000_021, w_000_022, w_000_023, w_000_024, w_000_025, w_000_026, w_000_027, w_000_028, w_000_029, w_000_030, w_000_031, w_000_032, w_000_033, w_000_034, w_000_035, w_000_036, w_000_037, w_000_038, w_000_039, w_000_040, w_000_041, w_000_042, w_000_043, w_000_044, w_000_045, w_000_046, w_000_047, w_000_048, w_000_049, w_000_050, w_000_051, w_000_052, w_000_053, w_000_054, w_000_055, w_000_056, w_000_057, w_000_058, w_000_059, w_000_060, w_000_061, w_000_062, w_000_064, w_000_065, w_000_066, w_000_067, w_000_068, w_000_069, w_000_070, w_000_071, w_000_072, w_000_073, w_000_074, w_000_076, w_000_077, w_000_078, w_000_079, w_000_082, w_000_083, w_000_084, w_000_085, w_000_086, w_000_087, w_000_088, w_000_089, w_000_090, w_000_091, w_000_092, w_000_096;
  output w_100_000, w_100_001, w_100_002, w_100_003, w_100_004, w_100_005, w_100_006, w_100_007, w_100_008, w_100_009, w_100_010, w_100_011, w_100_012, w_100_013, w_100_014, w_100_015, w_100_016, w_100_017, w_100_018, w_100_019, w_100_020, w_100_021, w_100_022, w_100_023, w_100_024, w_100_025, w_100_026, w_100_027, w_100_028, w_100_029, w_100_030, w_100_031, w_100_032, w_100_033, w_100_034, w_100_035, w_100_036, w_100_037, w_100_038, w_100_039;
  wire w_000_000, w_000_001, w_000_002, w_000_003, w_000_004, w_000_005, w_000_006, w_000_007, w_000_008, w_000_009, w_000_010, w_000_011, w_000_012, w_000_013, w_000_014, w_000_015, w_000_016, w_000_018, w_000_019, w_000_020, w_000_021, w_000_022, w_000_023, w_000_024, w_000_025, w_000_026, w_000_027, w_000_028, w_000_029, w_000_030, w_000_031, w_000_032, w_000_033, w_000_034, w_000_035, w_000_036, w_000_037, w_000_038, w_000_039, w_000_040, w_000_041, w_000_042, w_000_043, w_000_044, w_000_045, w_000_046, w_000_047, w_000_048, w_000_049, w_000_050, w_000_051, w_000_052, w_000_053, w_000_054, w_000_055, w_000_056, w_000_057, w_000_058, w_000_059, w_000_060, w_000_061, w_000_062, w_000_064, w_000_065, w_000_066, w_000_067, w_000_068, w_000_069, w_000_070, w_000_071, w_000_072, w_000_073, w_000_074, w_000_076, w_000_077, w_000_078, w_000_079, w_000_082, w_000_083, w_000_084, w_000_085, w_000_086, w_000_087, w_000_088, w_000_089, w_000_090, w_000_091, w_000_092, w_000_096;
  wire w_001_000, w_001_001, w_001_002, w_001_003, w_001_004, w_001_005, w_001_006, w_001_007, w_001_008, w_001_009, w_001_011, w_001_012, w_001_013, w_001_014, w_001_015, w_001_016, w_001_017, w_001_018, w_001_019, w_001_020, w_001_021, w_001_022, w_001_023, w_001_024, w_001_025, w_001_026, w_001_027, w_001_028, w_001_029, w_001_030, w_001_031;
  wire w_002_000, w_002_001, w_002_002, w_002_004, w_002_005, w_002_009, w_002_011, w_002_013, w_002_014, w_002_015, w_002_016, w_002_017, w_002_020, w_002_022, w_002_023, w_002_024, w_002_026, w_002_027, w_002_028, w_002_029, w_002_030, w_002_031, w_002_032, w_002_034, w_002_035, w_002_036, w_002_037, w_002_038, w_002_039, w_002_040, w_002_043, w_002_044, w_002_047, w_002_048, w_002_050, w_002_054, w_002_055, w_002_058, w_002_059, w_002_060, w_002_062, w_002_063, w_002_065, w_002_066, w_002_067, w_002_068, w_002_071, w_002_072, w_002_073, w_002_074, w_002_075, w_002_076, w_002_077, w_002_078, w_002_079, w_002_081, w_002_087, w_002_089, w_002_090, w_002_091, w_002_093, w_002_098;
  wire w_003_000, w_003_001, w_003_002, w_003_003, w_003_004, w_003_005, w_003_006, w_003_007, w_003_008, w_003_009, w_003_010, w_003_011, w_003_012, w_003_013, w_003_014, w_003_015, w_003_016, w_003_017, w_003_018, w_003_019, w_003_020, w_003_021, w_003_022, w_003_023;
  wire w_004_000, w_004_001, w_004_002, w_004_003, w_004_005, w_004_006, w_004_007, w_004_008, w_004_009, w_004_010, w_004_012, w_004_014, w_004_015, w_004_016, w_004_017, w_004_019, w_004_020, w_004_022, w_004_023, w_004_024, w_004_025, w_004_026, w_004_027, w_004_028, w_004_031, w_004_032, w_004_033, w_004_036, w_004_037, w_004_038, w_004_040;
  wire w_005_000, w_005_002, w_005_003, w_005_004, w_005_005, w_005_007, w_005_009, w_005_010, w_005_011, w_005_012, w_005_013, w_005_014, w_005_015, w_005_016, w_005_018;
  wire w_006_000;
  wire w_007_000, w_007_001, w_007_002, w_007_003, w_007_004, w_007_005, w_007_006, w_007_007;
  wire w_008_000, w_008_001, w_008_002, w_008_003, w_008_005, w_008_008, w_008_009, w_008_010, w_008_012, w_008_015, w_008_017, w_008_020, w_008_021, w_008_025, w_008_027, w_008_028, w_008_029, w_008_033, w_008_038, w_008_042, w_008_043, w_008_046, w_008_052, w_008_055, w_008_060, w_008_061, w_008_063, w_008_065, w_008_067, w_008_069, w_008_075, w_008_076, w_008_079, w_008_080, w_008_084;
  wire w_009_000, w_009_001, w_009_002, w_009_003, w_009_004, w_009_005, w_009_006, w_009_007, w_009_008, w_009_009, w_009_010, w_009_011, w_009_012, w_009_013;
  wire w_010_000, w_010_002, w_010_004, w_010_005, w_010_007, w_010_010, w_010_011, w_010_020, w_010_022, w_010_023, w_010_024, w_010_025, w_010_027, w_010_028, w_010_030, w_010_032, w_010_038, w_010_042, w_010_043, w_010_050, w_010_054, w_010_056, w_010_058, w_010_060, w_010_062, w_010_063;
  wire w_011_000, w_011_004, w_011_006, w_011_008, w_011_010, w_011_016, w_011_018, w_011_019, w_011_022, w_011_023, w_011_024, w_011_025, w_011_026, w_011_029, w_011_031, w_011_035, w_011_036, w_011_043, w_011_047, w_011_050, w_011_057, w_011_064, w_011_071, w_011_073, w_011_077;
  wire w_012_000, w_012_002, w_012_003, w_012_004, w_012_005, w_012_006, w_012_009, w_012_011, w_012_019, w_012_023, w_012_026, w_012_027, w_012_028, w_012_029, w_012_030, w_012_031, w_012_032, w_012_037, w_012_038, w_012_044, w_012_045, w_012_046, w_012_052, w_012_053, w_012_054, w_012_055, w_012_059, w_012_060, w_012_061, w_012_062, w_012_063, w_012_064, w_012_065, w_012_067;
  wire w_013_000;
  wire w_014_000, w_014_001, w_014_003, w_014_004, w_014_006, w_014_008, w_014_009, w_014_011, w_014_012, w_014_013, w_014_018, w_014_021, w_014_022, w_014_023, w_014_024, w_014_025, w_014_027;
  wire w_015_000, w_015_002, w_015_009, w_015_011, w_015_012, w_015_013, w_015_014, w_015_017, w_015_021, w_015_022, w_015_023, w_015_025, w_015_028, w_015_032, w_015_033;
  wire w_016_000, w_016_001, w_016_002, w_016_003, w_016_004, w_016_005, w_016_006;
  wire w_017_001, w_017_002, w_017_003, w_017_004, w_017_008, w_017_012, w_017_013, w_017_016, w_017_017, w_017_020, w_017_021, w_017_022, w_017_027, w_017_030, w_017_032, w_017_034, w_017_049, w_017_062, w_017_068;
  wire w_018_001, w_018_003, w_018_004, w_018_005, w_018_007, w_018_008, w_018_012, w_018_013, w_018_014, w_018_015, w_018_016, w_018_019, w_018_021, w_018_023, w_018_028, w_018_030, w_018_032, w_018_033;
  wire w_019_000, w_019_002, w_019_003, w_019_004, w_019_006, w_019_007, w_019_008, w_019_009, w_019_010, w_019_019, w_019_021, w_019_023, w_019_024;
  wire w_020_000, w_020_002, w_020_003, w_020_004, w_020_005, w_020_006, w_020_007, w_020_009, w_020_011, w_020_012, w_020_013, w_020_014, w_020_015, w_020_016, w_020_017, w_020_018, w_020_019, w_020_020;
  wire w_021_000, w_021_003, w_021_008, w_021_013, w_021_017, w_021_020, w_021_025, w_021_028, w_021_030, w_021_035, w_021_037, w_021_042, w_021_043, w_021_049, w_021_052;
  wire w_022_001, w_022_008, w_022_009, w_022_015, w_022_016, w_022_023, w_022_048, w_022_055;
  wire w_023_005, w_023_009, w_023_028, w_023_029, w_023_041, w_023_042, w_023_043, w_023_049, w_023_050, w_023_062, w_023_067, w_023_069, w_023_070, w_023_071, w_023_072, w_023_073, w_023_074, w_023_075, w_023_079, w_023_080, w_023_081, w_023_082, w_023_083, w_023_084, w_023_085, w_023_086, w_023_087, w_023_088, w_023_089, w_023_090, w_023_092;
  wire w_024_002, w_024_003, w_024_008, w_024_013, w_024_017, w_024_019, w_024_020, w_024_022, w_024_024, w_024_033, w_024_035, w_024_059;
  wire w_025_005, w_025_006, w_025_012, w_025_014, w_025_019, w_025_024, w_025_052, w_025_053, w_025_055, w_025_057;
  wire w_026_025, w_026_031, w_026_038, w_026_044, w_026_045, w_026_052, w_026_058, w_026_065, w_026_072, w_026_079, w_026_087, w_026_090, w_026_093;
  wire w_027_006, w_027_017, w_027_020, w_027_021, w_027_022, w_027_023, w_027_026, w_027_029, w_027_033, w_027_043, w_027_045;
  wire w_028_000, w_028_005, w_028_006, w_028_009, w_028_011, w_028_012, w_028_013, w_028_014, w_028_015, w_028_017, w_028_018;
  wire w_029_009, w_029_067, w_029_075, w_029_078;
  wire w_030_006, w_030_010, w_030_027, w_030_059, w_030_067, w_030_073;
  wire w_031_007, w_031_009, w_031_019, w_031_022, w_031_024, w_031_025, w_031_040, w_031_050, w_031_065;
  wire w_032_000, w_032_001, w_032_002, w_032_004, w_032_005, w_032_006, w_032_007, w_032_008, w_032_009, w_032_013, w_032_014, w_032_015, w_032_016, w_032_018;
  wire w_033_013, w_033_018, w_033_023, w_033_038, w_033_050, w_033_057, w_033_066;
  wire w_034_012, w_034_042, w_034_051, w_034_054, w_034_080;
  wire w_035_000, w_035_004, w_035_005, w_035_006, w_035_007;
  wire w_036_003, w_036_051, w_036_070;
  wire w_037_038, w_037_054, w_037_058, w_037_062, w_037_067, w_037_077;
  wire w_038_003, w_038_012, w_038_020, w_038_023, w_038_029, w_038_038;
  wire w_039_002, w_039_004, w_039_008, w_039_029, w_039_032, w_039_036;
  wire w_040_000, w_040_003, w_040_005, w_040_006;
  wire w_041_002, w_041_007, w_041_010, w_041_014, w_041_017, w_041_025, w_041_030, w_041_033, w_041_035;
  wire w_042_000, w_042_020, w_042_030, w_042_035;
  wire w_043_000, w_043_003, w_043_008, w_043_016, w_043_020, w_043_023, w_043_040, w_043_045, w_043_058, w_043_063;
  wire w_044_001, w_044_008, w_044_010, w_044_014, w_044_015, w_044_016, w_044_022, w_044_043, w_044_050;
  wire w_045_006, w_045_045;
  wire w_046_003, w_046_004, w_046_013, w_046_035, w_046_037, w_046_038, w_046_039, w_046_043, w_046_044, w_046_045, w_046_046, w_046_047, w_046_048, w_046_050;
  wire w_047_005, w_047_029, w_047_088, w_047_089, w_047_090, w_047_091, w_047_092, w_047_093, w_047_094, w_047_095, w_047_096, w_047_097, w_047_099, w_047_101, w_047_102, w_047_103, w_047_105;
  wire w_048_024, w_048_035, w_048_036, w_048_040;
  wire w_049_001, w_049_002, w_049_005;
  wire w_050_001, w_050_009;
  wire w_051_000, w_051_008;
  wire w_052_009, w_052_011, w_052_041, w_052_043, w_052_044, w_052_045, w_052_046, w_052_047, w_052_048;
  wire w_053_002, w_053_004, w_053_016, w_053_019, w_053_023, w_053_062;
  wire w_054_003, w_054_004, w_054_011, w_054_013, w_054_018, w_054_020;
  wire w_055_009, w_055_017, w_055_049;
  wire w_056_000, w_056_003, w_056_042;
  wire w_057_008, w_057_009, w_057_012;
  wire w_058_005, w_058_014, w_058_054, w_058_061;
  wire w_059_032;
  wire w_060_002, w_060_011;
  wire w_061_005, w_061_045;
  wire w_062_000, w_062_001, w_062_002, w_062_004, w_062_005, w_062_006, w_062_007, w_062_008, w_062_009, w_062_010, w_062_011, w_062_012;
  wire w_063_023, w_063_028;
  wire w_064_040;
  wire w_065_024, w_065_059;
  wire w_066_013;
  wire w_068_006, w_068_007;
  wire w_069_006, w_069_009, w_069_043, w_069_068;
  wire w_070_006, w_070_043, w_070_080, w_070_081, w_070_082;
  wire w_071_013, w_071_030, w_071_080;
  wire w_072_027;
  wire w_073_020;
  wire w_076_031, w_076_065;
  wire w_077_008;
  wire w_078_027, w_078_055;
  wire w_079_006;
  wire w_080_019, w_080_020;
  wire w_082_001;
  wire w_083_005;
  wire w_084_002, w_084_005, w_084_006, w_084_007, w_084_008, w_084_009, w_084_010, w_084_011, w_084_012, w_084_016, w_084_017, w_084_018, w_084_019, w_084_020, w_084_021, w_084_022, w_084_023, w_084_024, w_084_025, w_084_026, w_084_027, w_084_029;
  wire w_085_032, w_085_086;
  wire w_088_010, w_088_017;
  wire w_089_016, w_089_054;
  wire w_091_023;
  wire w_092_059;
  wire w_093_010, w_093_030;
  wire w_094_028, w_094_033;
  wire w_095_000, w_095_001, w_095_002;
  wire w_096_039;
  wire w_097_046, w_097_047, w_097_048, w_097_049, w_097_050;
  wire w_098_002;
  wire w_100_000, w_100_001, w_100_002, w_100_003, w_100_004, w_100_005, w_100_006, w_100_007, w_100_008, w_100_009, w_100_010, w_100_011, w_100_012, w_100_013, w_100_014, w_100_015, w_100_016, w_100_017, w_100_018, w_100_019, w_100_020, w_100_021, w_100_022, w_100_023, w_100_024, w_100_025, w_100_026, w_100_027, w_100_028, w_100_029, w_100_030, w_100_031, w_100_032, w_100_033, w_100_034, w_100_035, w_100_036, w_100_037, w_100_038, w_100_039;
  not1 I001_000(w_001_000, w_000_000);
  nand2 I001_001(w_001_001, w_000_001, w_000_002);
  not1 I001_002(w_001_002, w_000_003);
  or2  I001_003(w_001_003, w_000_004, w_000_005);
  nand2 I001_004(w_001_004, w_000_006, w_000_007);
  nand2 I001_005(w_001_005, w_000_008, w_000_009);
  not1 I001_006(w_001_006, w_000_010);
  and2 I001_007(w_001_007, w_000_011, w_000_012);
  nand2 I001_008(w_001_008, w_000_013, w_000_014);
  not1 I001_009(w_001_009, w_000_015);
  or2  I001_011(w_001_011, w_000_002, w_000_018);
  not1 I001_012(w_001_012, w_000_019);
  nand2 I001_013(w_001_013, w_000_020, w_000_021);
  nand2 I001_014(w_001_014, w_000_022, w_000_023);
  or2  I001_015(w_001_015, w_000_021, w_000_019);
  and2 I001_016(w_001_016, w_000_024, w_000_025);
  and2 I001_017(w_001_017, w_000_015, w_000_026);
  or2  I001_018(w_001_018, w_000_026, w_000_027);
  and2 I001_019(w_001_019, w_000_028, w_000_029);
  not1 I001_020(w_001_020, w_000_030);
  and2 I001_021(w_001_021, w_000_031, w_000_005);
  or2  I001_022(w_001_022, w_000_032, w_000_027);
  and2 I001_023(w_001_023, w_000_005, w_000_033);
  or2  I001_024(w_001_024, w_000_013, w_000_034);
  and2 I001_025(w_001_025, w_000_035, w_000_036);
  or2  I001_026(w_001_026, w_000_014, w_000_037);
  not1 I001_027(w_001_027, w_000_038);
  nand2 I001_028(w_001_028, w_000_039, w_000_040);
  and2 I001_029(w_001_029, w_000_041, w_000_042);
  and2 I001_030(w_001_030, w_000_043, w_000_003);
  nand2 I001_031(w_001_031, w_000_044, w_000_045);
  and2 I002_000(w_002_000, w_000_046, w_001_012);
  not1 I002_001(w_002_001, w_000_047);
  nand2 I002_002(w_002_002, w_001_006, w_000_048);
  and2 I002_004(w_002_004, w_000_049, w_001_016);
  not1 I002_005(w_002_005, w_001_001);
  or2  I002_009(w_002_009, w_001_022, w_001_006);
  and2 I002_011(w_002_011, w_001_003, w_001_006);
  and2 I002_013(w_002_013, w_001_018, w_001_014);
  nand2 I002_014(w_002_014, w_001_023, w_001_024);
  and2 I002_015(w_002_015, w_000_041, w_000_051);
  and2 I002_016(w_002_016, w_000_052, w_000_014);
  nand2 I002_017(w_002_017, w_000_043, w_001_027);
  or2  I002_020(w_002_020, w_000_054, w_001_005);
  nand2 I002_022(w_002_022, w_000_029, w_000_004);
  nand2 I002_023(w_002_023, w_001_013, w_000_006);
  and2 I002_024(w_002_024, w_000_018, w_000_055);
  nand2 I002_026(w_002_026, w_000_056, w_000_057);
  and2 I002_027(w_002_027, w_001_012, w_000_005);
  nand2 I002_028(w_002_028, w_000_058, w_001_018);
  not1 I002_029(w_002_029, w_000_059);
  nand2 I002_030(w_002_030, w_001_004, w_000_011);
  not1 I002_031(w_002_031, w_000_060);
  nand2 I002_032(w_002_032, w_000_061, w_000_022);
  not1 I002_034(w_002_034, w_000_005);
  and2 I002_035(w_002_035, w_000_044, w_000_022);
  or2  I002_036(w_002_036, w_000_016, w_000_058);
  and2 I002_037(w_002_037, w_001_030, w_000_000);
  and2 I002_038(w_002_038, w_000_062, w_001_018);
  and2 I002_039(w_002_039, w_001_009, w_001_017);
  not1 I002_040(w_002_040, w_001_030);
  not1 I002_043(w_002_043, w_000_064);
  and2 I002_044(w_002_044, w_000_065, w_000_042);
  and2 I002_047(w_002_047, w_000_059, w_001_004);
  not1 I002_048(w_002_048, w_000_067);
  and2 I002_050(w_002_050, w_001_023, w_001_003);
  or2  I002_054(w_002_054, w_000_068, w_000_069);
  and2 I002_055(w_002_055, w_000_070, w_000_025);
  not1 I002_058(w_002_058, w_000_072);
  or2  I002_059(w_002_059, w_001_019, w_000_032);
  nand2 I002_060(w_002_060, w_000_004, w_001_005);
  not1 I002_062(w_002_062, w_001_020);
  or2  I002_063(w_002_063, w_001_021, w_001_004);
  and2 I002_065(w_002_065, w_000_002, w_000_073);
  or2  I002_066(w_002_066, w_000_068, w_000_074);
  and2 I002_067(w_002_067, w_000_058, w_000_036);
  and2 I002_068(w_002_068, w_001_016, w_001_001);
  and2 I002_071(w_002_071, w_000_076, w_001_017);
  not1 I002_072(w_002_072, w_001_001);
  nand2 I002_073(w_002_073, w_001_021, w_000_077);
  or2  I002_074(w_002_074, w_000_078, w_001_024);
  or2  I002_075(w_002_075, w_001_004, w_000_014);
  or2  I002_076(w_002_076, w_000_004, w_000_027);
  not1 I002_077(w_002_077, w_000_056);
  not1 I002_078(w_002_078, w_000_079);
  nand2 I002_079(w_002_079, w_001_007, w_000_028);
  nand2 I002_081(w_002_081, w_001_003, w_000_039);
  not1 I002_087(w_002_087, w_000_041);
  and2 I002_089(w_002_089, w_001_023, w_001_017);
  or2  I002_090(w_002_090, w_000_025, w_000_067);
  or2  I002_091(w_002_091, w_000_083, w_000_024);
  and2 I002_093(w_002_093, w_000_000, w_000_026);
  nand2 I002_098(w_002_098, w_000_084, w_000_055);
  or2  I003_000(w_003_000, w_002_055, w_002_020);
  or2  I003_001(w_003_001, w_000_085, w_001_002);
  not1 I003_002(w_003_002, w_001_024);
  or2  I003_003(w_003_003, w_000_060, w_001_005);
  or2  I003_004(w_003_004, w_001_017, w_000_045);
  nand2 I003_005(w_003_005, w_001_026, w_002_037);
  or2  I003_006(w_003_006, w_001_007, w_000_057);
  not1 I003_007(w_003_007, w_000_029);
  and2 I003_008(w_003_008, w_001_018, w_001_025);
  and2 I003_009(w_003_009, w_000_033, w_001_017);
  or2  I003_010(w_003_010, w_000_070, w_001_017);
  nand2 I003_011(w_003_011, w_002_063, w_001_030);
  or2  I003_012(w_003_012, w_001_031, w_001_018);
  not1 I003_013(w_003_013, w_002_091);
  or2  I003_014(w_003_014, w_000_021, w_002_074);
  nand2 I003_015(w_003_015, w_001_019, w_000_021);
  or2  I003_016(w_003_016, w_002_054, w_002_098);
  or2  I003_017(w_003_017, w_001_016, w_001_002);
  nand2 I003_018(w_003_018, w_000_086, w_001_006);
  and2 I003_019(w_003_019, w_000_021, w_000_062);
  and2 I003_020(w_003_020, w_000_077, w_001_004);
  and2 I003_021(w_003_021, w_000_083, w_002_059);
  or2  I003_022(w_003_022, w_001_003, w_000_027);
  not1 I003_023(w_003_023, w_002_060);
  or2  I004_000(w_004_000, w_003_001, w_000_011);
  or2  I004_001(w_004_001, w_002_091, w_003_007);
  not1 I004_002(w_004_002, w_001_004);
  or2  I004_003(w_004_003, w_002_005, w_002_022);
  or2  I004_005(w_004_005, w_002_026, w_001_022);
  or2  I004_006(w_004_006, w_003_002, w_002_013);
  nand2 I004_007(w_004_007, w_001_030, w_003_016);
  nand2 I004_008(w_004_008, w_002_032, w_002_017);
  not1 I004_009(w_004_009, w_003_013);
  nand2 I004_010(w_004_010, w_001_011, w_001_028);
  and2 I004_012(w_004_012, w_003_007, w_002_058);
  or2  I004_014(w_004_014, w_001_021, w_001_009);
  and2 I004_015(w_004_015, w_003_005, w_002_068);
  nand2 I004_016(w_004_016, w_001_006, w_003_015);
  or2  I004_017(w_004_017, w_000_067, w_002_063);
  and2 I004_019(w_004_019, w_003_022, w_002_011);
  not1 I004_020(w_004_020, w_000_087);
  nand2 I004_022(w_004_022, w_002_040, w_003_000);
  not1 I004_023(w_004_023, w_002_063);
  nand2 I004_024(w_004_024, w_002_030, w_001_014);
  nand2 I004_025(w_004_025, w_002_047, w_000_082);
  nand2 I004_026(w_004_026, w_000_004, w_002_043);
  not1 I004_027(w_004_027, w_002_040);
  not1 I004_028(w_004_028, w_003_014);
  not1 I004_031(w_004_031, w_003_021);
  or2  I004_032(w_004_032, w_001_015, w_003_004);
  or2  I004_033(w_004_033, w_002_001, w_003_005);
  and2 I004_035(w_004_037, w_004_036, w_003_023);
  or2  I004_036(w_004_038, w_004_037, w_003_017);
  or2  I004_037(w_004_036, w_004_038, w_001_014);
  and2 I005_000(w_005_000, w_004_008, w_004_028);
  nand2 I005_001(w_005_003, w_004_028, w_005_002);
  or2  I005_002(w_005_004, w_005_003, w_005_018);
  not1 I005_003(w_005_005, w_005_004);
  nand2 I005_004(w_005_002, w_004_005, w_005_005);
  and2 I005_005(w_005_010, w_005_009, w_003_020);
  nand2 I005_006(w_005_011, w_001_020, w_005_010);
  and2 I005_007(w_005_012, w_003_008, w_005_011);
  not1 I005_008(w_005_013, w_005_012);
  and2 I005_009(w_005_014, w_005_013, w_003_001);
  nand2 I005_010(w_005_015, w_005_014, w_004_023);
  or2  I005_011(w_005_016, w_002_016, w_005_015);
  not1 I005_012(w_005_009, w_005_004);
  and2 I005_013(w_005_018, w_004_010, w_005_016);
  and2 I005_014(w_004_040, w_000_089, w_004_036);
  and2 I006_000(w_006_000, w_000_015, w_000_071);
  and2 I006_001(w_005_007, w_004_040, w_005_002);
  nand2 I007_000(w_007_000, w_004_010, w_004_024);
  or2  I007_001(w_007_001, w_002_000, w_002_009);
  or2  I007_002(w_007_002, w_004_014, w_000_088);
  not1 I007_003(w_007_003, w_002_047);
  nand2 I007_004(w_007_004, w_004_031, w_005_000);
  or2  I007_005(w_007_005, w_002_050, w_001_026);
  not1 I007_006(w_007_006, w_002_031);
  or2  I007_007(w_007_007, w_005_007, w_001_017);
  and2 I008_000(w_008_000, w_001_018, w_005_000);
  nand2 I008_001(w_008_001, w_000_025, w_004_022);
  and2 I008_002(w_008_002, w_007_001, w_000_034);
  or2  I008_003(w_008_003, w_002_015, w_001_008);
  and2 I008_005(w_008_005, w_002_077, w_005_000);
  or2  I008_008(w_008_008, w_002_090, w_007_006);
  and2 I008_009(w_008_009, w_004_020, w_004_025);
  and2 I008_010(w_008_010, w_007_001, w_002_036);
  not1 I008_012(w_008_012, w_005_000);
  not1 I008_015(w_008_015, w_001_001);
  or2  I008_017(w_008_017, w_006_000, w_007_002);
  or2  I008_020(w_008_020, w_003_009, w_006_000);
  or2  I008_021(w_008_021, w_001_003, w_000_090);
  and2 I008_025(w_008_025, w_006_000, w_000_025);
  or2  I008_027(w_008_027, w_005_000, w_007_002);
  or2  I008_028(w_008_028, w_007_005, w_005_000);
  or2  I008_029(w_008_029, w_002_072, w_005_000);
  and2 I008_033(w_008_033, w_005_000, w_003_004);
  and2 I008_038(w_008_038, w_001_000, w_002_004);
  nand2 I008_042(w_008_042, w_007_005, w_007_004);
  or2  I008_043(w_008_043, w_001_026, w_001_009);
  or2  I008_046(w_008_046, w_003_007, w_001_004);
  or2  I008_052(w_008_052, w_006_000, w_000_083);
  and2 I008_055(w_008_055, w_000_029, w_006_000);
  or2  I008_060(w_008_060, w_004_005, w_006_000);
  nand2 I008_061(w_008_061, w_002_060, w_002_024);
  and2 I008_063(w_008_063, w_006_000, w_005_000);
  nand2 I008_065(w_008_065, w_006_000, w_001_026);
  nand2 I008_067(w_008_067, w_005_000, w_004_008);
  not1 I008_069(w_008_069, w_001_000);
  nand2 I008_075(w_008_075, w_005_000, w_007_002);
  not1 I008_076(w_008_076, w_004_024);
  nand2 I008_079(w_008_079, w_006_000, w_003_011);
  nand2 I008_080(w_008_080, w_005_000, w_002_087);
  and2 I008_084(w_008_084, w_005_000, w_003_013);
  not1 I009_000(w_009_000, w_006_000);
  or2  I009_001(w_009_001, w_002_087, w_003_003);
  or2  I009_002(w_009_002, w_005_000, w_002_048);
  not1 I009_003(w_009_003, w_005_000);
  nand2 I009_004(w_009_004, w_002_017, w_005_000);
  and2 I009_005(w_009_005, w_003_018, w_003_006);
  nand2 I009_006(w_009_006, w_008_033, w_008_017);
  and2 I009_007(w_009_007, w_005_000, w_001_013);
  nand2 I009_008(w_009_008, w_005_000, w_008_069);
  nand2 I009_009(w_009_009, w_002_076, w_002_071);
  and2 I009_010(w_009_010, w_004_008, w_002_091);
  or2  I009_011(w_009_011, w_000_066, w_006_000);
  not1 I009_012(w_009_012, w_001_024);
  or2  I009_013(w_009_013, w_007_006, w_006_000);
  and2 I010_000(w_010_000, w_005_000, w_002_039);
  not1 I010_002(w_010_002, w_003_007);
  nand2 I010_004(w_010_004, w_008_025, w_005_000);
  or2  I010_005(w_010_005, w_002_026, w_004_023);
  not1 I010_007(w_010_007, w_009_011);
  not1 I010_010(w_010_010, w_007_006);
  or2  I010_011(w_010_011, w_007_003, w_000_050);
  or2  I010_020(w_010_020, w_009_007, w_007_007);
  or2  I010_022(w_010_022, w_008_027, w_004_019);
  nand2 I010_023(w_010_023, w_001_023, w_008_002);
  nand2 I010_024(w_010_024, w_003_014, w_008_009);
  and2 I010_025(w_010_025, w_000_092, w_006_000);
  or2  I010_027(w_010_027, w_009_000, w_006_000);
  or2  I010_028(w_010_028, w_002_078, w_003_018);
  not1 I010_030(w_010_030, w_002_059);
  nand2 I010_032(w_010_032, w_005_000, w_007_002);
  or2  I010_038(w_010_038, w_009_006, w_006_000);
  or2  I010_042(w_010_042, w_008_076, w_007_005);
  not1 I010_043(w_010_043, w_000_062);
  not1 I010_050(w_010_050, w_002_034);
  or2  I010_054(w_010_054, w_007_005, w_002_081);
  or2  I010_056(w_010_056, w_004_028, w_005_000);
  and2 I010_058(w_010_058, w_003_018, w_001_000);
  not1 I010_060(w_010_060, w_003_009);
  not1 I010_062(w_010_062, w_002_044);
  nand2 I010_063(w_010_063, w_003_014, w_001_019);
  nand2 I011_000(w_011_000, w_007_005, w_004_014);
  and2 I011_004(w_011_004, w_001_007, w_007_002);
  or2  I011_006(w_011_006, w_008_067, w_000_035);
  or2  I011_008(w_011_008, w_008_005, w_001_015);
  and2 I011_010(w_011_010, w_008_055, w_000_066);
  and2 I011_016(w_011_016, w_004_016, w_010_023);
  nand2 I011_018(w_011_018, w_007_007, w_010_062);
  and2 I011_019(w_011_019, w_006_000, w_004_033);
  or2  I011_022(w_011_022, w_006_000, w_008_080);
  and2 I011_023(w_011_023, w_007_007, w_009_012);
  not1 I011_024(w_011_024, w_003_011);
  or2  I011_025(w_011_025, w_002_073, w_008_038);
  nand2 I011_026(w_011_026, w_010_058, w_003_022);
  and2 I011_029(w_011_029, w_008_052, w_000_004);
  or2  I011_031(w_011_031, w_004_001, w_002_060);
  and2 I011_035(w_011_035, w_009_002, w_009_013);
  not1 I011_036(w_011_036, w_009_003);
  or2  I011_043(w_011_043, w_001_005, w_002_028);
  and2 I011_047(w_011_047, w_000_090, w_005_000);
  nand2 I011_050(w_011_050, w_010_020, w_002_038);
  and2 I011_057(w_011_057, w_010_030, w_003_001);
  nand2 I011_064(w_011_064, w_000_054, w_006_000);
  not1 I011_071(w_011_071, w_009_009);
  not1 I011_073(w_011_073, w_001_004);
  or2  I011_077(w_011_077, w_006_000, w_008_008);
  not1 I012_000(w_012_000, w_003_002);
  not1 I012_002(w_012_002, w_003_013);
  and2 I012_003(w_012_003, w_010_004, w_007_007);
  nand2 I012_004(w_012_004, w_007_003, w_000_020);
  or2  I012_005(w_012_005, w_008_003, w_005_000);
  not1 I012_006(w_012_006, w_001_014);
  nand2 I012_009(w_012_009, w_001_026, w_011_035);
  not1 I012_011(w_012_011, w_000_049);
  not1 I012_019(w_012_019, w_008_079);
  not1 I012_023(w_012_023, w_008_065);
  not1 I012_026(w_012_026, w_008_063);
  not1 I012_027(w_012_027, w_002_027);
  not1 I012_028(w_012_028, w_008_033);
  not1 I012_029(w_012_029, w_006_000);
  or2  I012_030(w_012_030, w_007_003, w_003_023);
  or2  I012_031(w_012_031, w_005_000, w_010_060);
  or2  I012_032(w_012_032, w_007_004, w_003_019);
  not1 I012_037(w_012_037, w_001_004);
  and2 I012_038(w_012_038, w_006_000, w_001_014);
  and2 I012_044(w_012_044, w_003_012, w_004_012);
  nand2 I012_045(w_012_045, w_005_000, w_011_010);
  or2  I012_046(w_012_046, w_002_066, w_003_015);
  not1 I012_051(w_012_053, w_012_052);
  not1 I012_052(w_012_054, w_012_053);
  and2 I012_053(w_012_055, w_012_054, w_012_067);
  not1 I012_054(w_012_052, w_012_055);
  not1 I012_055(w_012_060, w_012_059);
  not1 I012_056(w_012_061, w_012_060);
  and2 I012_057(w_012_062, w_012_061, w_008_028);
  nand2 I012_058(w_012_063, w_012_062, w_003_007);
  not1 I012_059(w_012_064, w_012_063);
  and2 I012_060(w_012_065, w_012_064, w_004_019);
  not1 I012_061(w_012_059, w_012_055);
  and2 I012_062(w_012_067, w_001_017, w_012_065);
  and2 I013_000(w_013_000, w_005_000, w_003_018);
  or2  I014_000(w_014_000, w_004_001, w_006_000);
  nand2 I014_001(w_014_001, w_002_055, w_009_005);
  and2 I014_003(w_014_003, w_001_004, w_004_010);
  and2 I014_004(w_014_004, w_006_000, w_009_010);
  or2  I014_006(w_014_006, w_003_023, w_011_000);
  nand2 I014_008(w_014_008, w_008_029, w_008_001);
  not1 I014_009(w_014_009, w_012_045);
  not1 I014_011(w_014_011, w_008_005);
  or2  I014_012(w_014_012, w_000_030, w_011_047);
  nand2 I014_013(w_014_013, w_010_000, w_002_029);
  nand2 I014_018(w_014_018, w_003_001, w_011_010);
  and2 I014_021(w_014_021, w_007_000, w_002_062);
  nand2 I014_022(w_014_022, w_007_002, w_003_023);
  or2  I014_023(w_014_023, w_004_026, w_000_072);
  nand2 I014_024(w_014_024, w_013_000, w_001_030);
  not1 I014_025(w_014_025, w_012_006);
  not1 I014_027(w_014_027, w_006_000);
  or2  I015_000(w_015_000, w_014_025, w_002_065);
  nand2 I015_002(w_015_002, w_010_010, w_010_024);
  or2  I015_009(w_015_009, w_004_016, w_008_060);
  nand2 I015_011(w_015_011, w_000_070, w_001_013);
  nand2 I015_012(w_015_012, w_014_000, w_007_006);
  or2  I015_013(w_015_013, w_005_000, w_013_000);
  or2  I015_014(w_015_014, w_002_089, w_012_002);
  and2 I015_017(w_015_017, w_012_032, w_012_045);
  or2  I015_021(w_015_021, w_013_000, w_003_017);
  not1 I015_022(w_015_022, w_008_080);
  and2 I015_023(w_015_023, w_001_006, w_004_000);
  and2 I015_025(w_015_025, w_007_001, w_000_025);
  and2 I015_028(w_015_028, w_008_061, w_000_038);
  nand2 I015_032(w_015_032, w_003_013, w_000_096);
  and2 I015_033(w_015_033, w_011_018, w_001_013);
  nand2 I016_000(w_016_000, w_014_006, w_008_010);
  not1 I016_001(w_016_001, w_009_004);
  and2 I016_002(w_016_002, w_011_006, w_003_003);
  and2 I016_003(w_016_003, w_009_005, w_002_039);
  and2 I016_004(w_016_004, w_014_022, w_008_043);
  not1 I016_005(w_016_005, w_012_019);
  and2 I016_006(w_016_006, w_010_011, w_009_011);
  or2  I017_001(w_017_001, w_015_009, w_010_030);
  and2 I017_002(w_017_002, w_012_000, w_008_020);
  not1 I017_003(w_017_003, w_012_005);
  or2  I017_004(w_017_004, w_014_000, w_004_015);
  not1 I017_008(w_017_008, w_003_002);
  nand2 I017_012(w_017_012, w_010_005, w_010_011);
  or2  I017_013(w_017_013, w_001_003, w_005_000);
  nand2 I017_016(w_017_016, w_014_009, w_012_004);
  nand2 I017_017(w_017_017, w_016_002, w_014_004);
  and2 I017_020(w_017_020, w_015_012, w_016_002);
  or2  I017_021(w_017_021, w_000_086, w_004_006);
  or2  I017_022(w_017_022, w_004_002, w_016_003);
  and2 I017_027(w_017_027, w_001_003, w_000_034);
  or2  I017_030(w_017_030, w_002_048, w_008_000);
  or2  I017_032(w_017_032, w_006_000, w_008_021);
  or2  I017_034(w_017_034, w_009_006, w_015_002);
  or2  I017_049(w_017_049, w_009_011, w_012_029);
  not1 I017_062(w_017_062, w_012_023);
  not1 I017_068(w_017_068, w_002_067);
  or2  I018_001(w_018_001, w_005_000, w_007_001);
  and2 I018_003(w_018_003, w_007_007, w_008_001);
  and2 I018_004(w_018_004, w_009_012, w_000_032);
  nand2 I018_005(w_018_005, w_014_011, w_012_037);
  or2  I018_007(w_018_007, w_013_000, w_006_000);
  nand2 I018_008(w_018_008, w_011_073, w_011_057);
  nand2 I018_012(w_018_012, w_016_000, w_012_026);
  or2  I018_013(w_018_013, w_002_071, w_016_003);
  nand2 I018_014(w_018_014, w_002_087, w_002_079);
  or2  I018_015(w_018_015, w_013_000, w_012_009);
  and2 I018_016(w_018_016, w_000_066, w_011_029);
  not1 I018_019(w_018_019, w_009_001);
  or2  I018_021(w_018_021, w_008_042, w_011_000);
  or2  I018_023(w_018_023, w_008_038, w_016_003);
  nand2 I018_028(w_018_028, w_010_054, w_009_000);
  and2 I018_030(w_018_030, w_012_032, w_015_022);
  nand2 I018_032(w_018_032, w_009_012, w_003_023);
  not1 I018_033(w_018_033, w_013_000);
  or2  I019_000(w_019_000, w_017_022, w_007_007);
  or2  I019_002(w_019_002, w_011_026, w_001_001);
  nand2 I019_003(w_019_003, w_017_020, w_003_008);
  not1 I019_004(w_019_004, w_016_002);
  and2 I019_006(w_019_006, w_007_001, w_003_003);
  or2  I019_007(w_019_007, w_011_023, w_013_000);
  not1 I019_008(w_019_008, w_003_009);
  and2 I019_009(w_019_009, w_014_003, w_013_000);
  not1 I019_010(w_019_010, w_008_000);
  nand2 I019_019(w_019_019, w_008_015, w_018_001);
  or2  I019_021(w_019_021, w_009_008, w_018_021);
  and2 I019_023(w_019_023, w_001_025, w_012_027);
  nand2 I019_024(w_019_024, w_010_056, w_004_012);
  nand2 I020_000(w_020_000, w_003_005, w_016_000);
  and2 I020_002(w_020_002, w_006_000, w_004_002);
  not1 I020_003(w_020_003, w_015_011);
  not1 I020_004(w_020_004, w_004_024);
  nand2 I020_005(w_020_005, w_009_009, w_013_000);
  or2  I020_006(w_020_006, w_002_035, w_017_003);
  not1 I020_007(w_020_007, w_000_001);
  nand2 I020_009(w_020_009, w_015_033, w_007_003);
  nand2 I020_010(w_020_012, w_019_002, w_020_011);
  or2  I020_011(w_020_013, w_020_012, w_019_007);
  not1 I020_012(w_020_014, w_020_013);
  and2 I020_013(w_020_015, w_016_000, w_020_014);
  and2 I020_014(w_020_016, w_008_075, w_020_015);
  not1 I020_015(w_020_017, w_020_016);
  and2 I020_016(w_020_018, w_016_004, w_020_017);
  or2  I020_017(w_020_019, w_008_001, w_020_018);
  or2  I020_018(w_020_020, w_007_007, w_020_019);
  or2  I020_019(w_020_011, w_019_019, w_020_020);
  not1 I021_000(w_021_000, w_003_017);
  nand2 I021_003(w_021_003, w_011_016, w_018_015);
  or2  I021_008(w_021_008, w_001_006, w_007_001);
  and2 I021_013(w_021_013, w_015_014, w_008_001);
  or2  I021_017(w_021_017, w_006_000, w_008_046);
  nand2 I021_020(w_021_020, w_015_023, w_003_006);
  and2 I021_025(w_021_025, w_006_000, w_005_000);
  or2  I021_028(w_021_028, w_011_077, w_020_000);
  not1 I021_030(w_021_030, w_003_010);
  and2 I021_035(w_021_035, w_017_068, w_019_006);
  or2  I021_037(w_021_037, w_009_012, w_016_000);
  not1 I021_042(w_021_042, w_016_005);
  and2 I021_043(w_021_043, w_007_006, w_006_000);
  nand2 I021_049(w_021_049, w_010_002, w_018_007);
  not1 I021_052(w_021_052, w_020_009);
  not1 I022_001(w_022_001, w_017_049);
  and2 I022_008(w_022_008, w_005_000, w_003_000);
  or2  I022_009(w_022_009, w_014_011, w_012_046);
  nand2 I022_015(w_022_015, w_017_002, w_000_091);
  and2 I022_016(w_022_016, w_012_030, w_015_009);
  not1 I022_023(w_022_023, w_018_030);
  not1 I022_048(w_022_048, w_010_028);
  or2  I022_055(w_022_055, w_018_005, w_008_012);
  not1 I023_005(w_023_005, w_013_000);
  nand2 I023_009(w_023_009, w_012_045, w_019_023);
  or2  I023_028(w_023_028, w_021_000, w_014_013);
  not1 I023_029(w_023_029, w_004_003);
  not1 I023_041(w_023_041, w_013_000);
  or2  I023_042(w_023_042, w_000_086, w_020_005);
  or2  I023_043(w_023_043, w_010_007, w_020_002);
  nand2 I023_049(w_023_049, w_009_003, w_018_005);
  and2 I023_050(w_023_050, w_022_001, w_000_088);
  or2  I023_062(w_023_062, w_007_004, w_017_021);
  or2  I023_067(w_023_067, w_004_026, w_007_004);
  nand2 I023_068(w_023_070, w_009_007, w_023_069);
  not1 I023_069(w_023_071, w_023_070);
  nand2 I023_070(w_023_072, w_023_071, w_023_092);
  nand2 I023_071(w_023_073, w_023_072, w_001_015);
  not1 I023_072(w_023_074, w_023_073);
  and2 I023_073(w_023_075, w_023_074, w_001_005);
  not1 I023_074(w_023_069, w_023_075);
  not1 I023_075(w_023_080, w_023_079);
  nand2 I023_076(w_023_081, w_005_007, w_023_080);
  and2 I023_077(w_023_082, w_014_024, w_023_081);
  or2  I023_078(w_023_083, w_023_082, w_012_065);
  or2  I023_079(w_023_084, w_001_031, w_023_083);
  or2  I023_080(w_023_085, w_002_066, w_023_084);
  nand2 I023_081(w_023_086, w_001_003, w_023_085);
  or2  I023_082(w_023_087, w_023_086, w_010_063);
  and2 I023_083(w_023_088, w_016_004, w_023_087);
  nand2 I023_084(w_023_089, w_023_088, w_006_000);
  not1 I023_085(w_023_090, w_023_089);
  not1 I023_086(w_023_079, w_023_072);
  and2 I023_087(w_023_092, w_012_003, w_023_090);
  and2 I024_002(w_024_002, w_020_004, w_003_018);
  not1 I024_003(w_024_003, w_003_003);
  and2 I024_008(w_024_008, w_003_019, w_019_019);
  not1 I024_013(w_024_013, w_004_014);
  and2 I024_017(w_024_017, w_023_005, w_014_000);
  or2  I024_019(w_024_019, w_006_000, w_015_032);
  nand2 I024_020(w_024_020, w_019_009, w_001_029);
  not1 I024_022(w_024_022, w_000_058);
  and2 I024_024(w_024_024, w_017_013, w_008_027);
  not1 I024_033(w_024_033, w_016_001);
  or2  I024_035(w_024_035, w_007_005, w_000_082);
  or2  I024_059(w_024_059, w_003_021, w_020_006);
  not1 I025_005(w_025_005, w_012_003);
  nand2 I025_006(w_025_006, w_019_024, w_001_018);
  or2  I025_012(w_025_012, w_017_027, w_005_000);
  or2  I025_014(w_025_014, w_018_014, w_003_016);
  not1 I025_019(w_025_019, w_015_023);
  or2  I025_024(w_025_024, w_021_020, w_016_005);
  nand2 I025_052(w_025_052, w_021_013, w_021_025);
  or2  I025_053(w_025_053, w_014_027, w_011_071);
  nand2 I025_055(w_025_055, w_007_004, w_014_021);
  nand2 I025_057(w_025_057, w_001_000, w_015_021);
  nand2 I026_025(w_026_025, w_006_000, w_005_000);
  or2  I026_031(w_026_031, w_005_000, w_012_038);
  or2  I026_038(w_026_038, w_016_000, w_023_067);
  nand2 I026_044(w_026_044, w_010_043, w_016_003);
  nand2 I026_045(w_026_045, w_018_004, w_025_012);
  and2 I026_052(w_026_052, w_006_000, w_013_000);
  nand2 I026_058(w_026_058, w_024_013, w_023_062);
  and2 I026_065(w_026_065, w_006_000, w_017_001);
  nand2 I026_072(w_026_072, w_019_000, w_021_017);
  or2  I026_079(w_026_079, w_022_009, w_002_017);
  nand2 I026_087(w_026_087, w_018_021, w_018_033);
  nand2 I026_090(w_026_090, w_001_018, w_011_004);
  or2  I026_093(w_026_093, w_014_012, w_003_014);
  not1 I027_006(w_027_006, w_018_005);
  and2 I027_017(w_027_017, w_015_013, w_002_079);
  nand2 I027_020(w_027_020, w_014_000, w_011_008);
  nand2 I027_021(w_027_021, w_007_001, w_004_032);
  nand2 I027_022(w_027_022, w_005_000, w_012_011);
  and2 I027_023(w_027_023, w_013_000, w_026_038);
  and2 I027_026(w_027_026, w_018_032, w_026_065);
  not1 I027_029(w_027_029, w_008_029);
  nand2 I027_033(w_027_033, w_006_000, w_010_042);
  and2 I027_043(w_027_043, w_011_023, w_000_039);
  nand2 I027_045(w_027_045, w_026_090, w_015_017);
  nand2 I028_000(w_028_000, w_000_050, w_021_030);
  and2 I028_005(w_028_005, w_019_024, w_027_022);
  nand2 I028_006(w_028_006, w_023_028, w_018_016);
  not1 I028_009(w_028_009, w_007_005);
  and2 I028_011(w_028_011, w_023_009, w_006_000);
  and2 I028_012(w_028_012, w_027_017, w_004_005);
  not1 I028_013(w_028_013, w_011_031);
  nand2 I028_014(w_028_014, w_014_018, w_011_024);
  not1 I028_015(w_028_015, w_014_003);
  and2 I028_017(w_028_017, w_006_000, w_001_008);
  and2 I028_018(w_028_018, w_001_020, w_024_002);
  and2 I029_009(w_029_009, w_000_053, w_020_003);
  or2  I029_067(w_029_067, w_023_043, w_009_006);
  nand2 I029_075(w_029_075, w_021_008, w_028_013);
  nand2 I029_078(w_029_078, w_010_050, w_028_017);
  or2  I030_006(w_030_006, w_027_026, w_004_001);
  or2  I030_010(w_030_010, w_003_012, w_002_002);
  or2  I030_027(w_030_027, w_010_038, w_003_009);
  not1 I030_059(w_030_059, w_011_019);
  nand2 I030_067(w_030_067, w_018_005, w_024_003);
  nand2 I030_073(w_030_073, w_002_059, w_028_006);
  not1 I031_007(w_031_007, w_004_009);
  or2  I031_009(w_031_009, w_026_079, w_014_023);
  and2 I031_019(w_031_019, w_017_062, w_018_012);
  nand2 I031_022(w_031_022, w_025_024, w_000_030);
  nand2 I031_024(w_031_024, w_026_044, w_004_002);
  nand2 I031_025(w_031_025, w_028_000, w_011_022);
  not1 I031_040(w_031_040, w_011_036);
  or2  I031_050(w_031_050, w_010_032, w_002_001);
  nand2 I031_065(w_031_065, w_028_015, w_020_007);
  or2  I032_000(w_032_000, w_006_000, w_004_007);
  and2 I032_001(w_032_001, w_010_025, w_019_010);
  or2  I032_002(w_032_002, w_000_016, w_017_012);
  or2  I032_003(w_032_005, w_010_027, w_032_004);
  not1 I032_004(w_032_006, w_032_005);
  nand2 I032_005(w_032_007, w_032_006, w_032_018);
  and2 I032_006(w_032_008, w_027_022, w_032_007);
  and2 I032_007(w_032_009, w_032_008, w_031_065);
  and2 I032_008(w_032_004, w_032_009, w_024_035);
  and2 I032_009(w_032_014, w_032_013, w_028_012);
  or2  I032_010(w_032_015, w_032_014, w_009_011);
  and2 I032_011(w_032_016, w_032_015, w_001_024);
  not1 I032_012(w_032_013, w_032_007);
  and2 I032_013(w_032_018, w_028_012, w_032_016);
  not1 I033_013(w_033_013, w_015_028);
  and2 I033_018(w_033_018, w_010_024, w_024_033);
  nand2 I033_023(w_033_023, w_013_000, w_003_004);
  or2  I033_038(w_033_038, w_011_064, w_026_072);
  not1 I033_050(w_033_050, w_018_023);
  not1 I033_057(w_033_057, w_026_052);
  not1 I033_066(w_033_066, w_000_046);
  nand2 I034_012(w_034_012, w_025_055, w_028_018);
  not1 I034_042(w_034_042, w_005_000);
  or2  I034_051(w_034_051, w_025_019, w_009_009);
  not1 I034_054(w_034_054, w_032_001);
  nand2 I034_080(w_034_080, w_018_021, w_005_000);
  and2 I035_000(w_035_000, w_017_008, w_020_000);
  or2  I035_004(w_035_004, w_001_014, w_012_045);
  and2 I035_005(w_035_005, w_026_025, w_001_007);
  or2  I035_006(w_035_006, w_027_029, w_024_020);
  or2  I035_007(w_035_007, w_009_002, w_017_027);
  or2  I036_003(w_036_003, w_028_005, w_025_014);
  nand2 I036_051(w_036_051, w_012_044, w_026_093);
  not1 I036_070(w_036_070, w_003_015);
  and2 I037_038(w_037_038, w_004_027, w_023_049);
  not1 I037_054(w_037_054, w_034_080);
  not1 I037_058(w_037_058, w_016_004);
  nand2 I037_062(w_037_062, w_030_067, w_008_052);
  or2  I037_067(w_037_067, w_020_000, w_019_023);
  and2 I037_077(w_037_077, w_005_000, w_019_002);
  not1 I038_003(w_038_003, w_012_031);
  not1 I038_012(w_038_012, w_034_042);
  not1 I038_020(w_038_020, w_005_000);
  nand2 I038_023(w_038_023, w_021_042, w_022_008);
  nand2 I038_029(w_038_029, w_032_000, w_029_067);
  and2 I038_038(w_038_038, w_015_025, w_004_028);
  and2 I039_002(w_039_002, w_014_018, w_012_028);
  not1 I039_004(w_039_004, w_004_008);
  and2 I039_008(w_039_008, w_031_065, w_007_005);
  and2 I039_029(w_039_029, w_031_025, w_021_043);
  and2 I039_032(w_039_032, w_019_024, w_021_035);
  and2 I039_036(w_039_036, w_032_000, w_006_000);
  or2  I040_000(w_040_000, w_018_001, w_010_005);
  and2 I040_003(w_040_003, w_032_001, w_016_006);
  not1 I040_005(w_040_005, w_027_021);
  nand2 I040_006(w_040_006, w_000_088, w_032_001);
  nand2 I041_002(w_041_002, w_009_002, w_035_004);
  or2  I041_007(w_041_007, w_023_050, w_010_020);
  nand2 I041_010(w_041_010, w_040_006, w_025_006);
  not1 I041_014(w_041_014, w_018_008);
  or2  I041_017(w_041_017, w_014_001, w_015_017);
  nand2 I041_025(w_041_025, w_009_002, w_004_010);
  or2  I041_030(w_041_030, w_033_038, w_005_000);
  nand2 I041_033(w_041_033, w_036_003, w_024_017);
  nand2 I041_035(w_041_035, w_008_076, w_002_023);
  nand2 I042_000(w_042_000, w_002_014, w_025_057);
  or2  I042_020(w_042_020, w_009_005, w_010_022);
  and2 I042_030(w_042_030, w_018_021, w_004_017);
  nand2 I042_035(w_042_035, w_001_001, w_031_019);
  nand2 I043_000(w_043_000, w_040_003, w_031_024);
  and2 I043_003(w_043_003, w_026_045, w_026_087);
  and2 I043_008(w_043_008, w_038_023, w_000_092);
  and2 I043_016(w_043_016, w_022_055, w_037_077);
  not1 I043_020(w_043_020, w_014_023);
  and2 I043_023(w_043_023, w_030_073, w_003_003);
  not1 I043_040(w_043_040, w_009_013);
  not1 I043_045(w_043_045, w_024_019);
  not1 I043_058(w_043_058, w_009_009);
  not1 I043_063(w_043_063, w_011_043);
  nand2 I044_001(w_044_001, w_018_019, w_022_016);
  or2  I044_008(w_044_008, w_032_000, w_024_024);
  and2 I044_010(w_044_010, w_032_002, w_025_005);
  or2  I044_014(w_044_014, w_019_008, w_002_075);
  not1 I044_015(w_044_015, w_032_001);
  and2 I044_016(w_044_016, w_038_020, w_000_046);
  or2  I044_022(w_044_022, w_043_000, w_001_001);
  or2  I044_043(w_044_043, w_023_029, w_028_012);
  and2 I044_050(w_044_050, w_021_028, w_008_084);
  and2 I045_006(w_045_006, w_041_014, w_023_042);
  and2 I045_045(w_045_045, w_003_006, w_025_019);
  nand2 I046_003(w_046_003, w_002_014, w_043_045);
  not1 I046_004(w_046_004, w_019_003);
  not1 I046_013(w_046_013, w_034_054);
  and2 I046_035(w_046_035, w_029_075, w_038_003);
  not1 I046_036(w_046_038, w_046_037);
  and2 I046_037(w_046_039, w_046_038, w_011_050);
  and2 I046_038(w_046_037, w_046_050, w_046_039);
  not1 I046_039(w_046_044, w_046_043);
  nand2 I046_040(w_046_045, w_021_049, w_046_044);
  not1 I046_041(w_046_046, w_046_045);
  or2  I046_042(w_046_047, w_046_046, w_044_043);
  and2 I046_043(w_046_048, w_046_047, w_043_003);
  not1 I046_044(w_046_043, w_046_037);
  and2 I046_045(w_046_050, w_044_022, w_046_048);
  nand2 I047_005(w_047_005, w_001_031, w_014_003);
  and2 I047_029(w_047_029, w_034_051, w_036_051);
  nand2 I047_088(w_047_089, w_017_062, w_047_088);
  nand2 I047_089(w_047_090, w_047_089, w_017_004);
  or2  I047_090(w_047_091, w_047_090, w_039_008);
  nand2 I047_091(w_047_092, w_047_091, w_040_005);
  and2 I047_092(w_047_093, w_047_092, w_031_040);
  and2 I047_093(w_047_094, w_033_057, w_047_093);
  or2  I047_094(w_047_095, w_047_105, w_047_094);
  nand2 I047_095(w_047_096, w_025_053, w_047_095);
  nand2 I047_096(w_047_097, w_047_096, w_042_035);
  nand2 I047_097(w_047_088, w_047_097, w_046_039);
  and2 I047_098(w_047_102, w_047_101, w_012_064);
  nand2 I047_099(w_047_103, w_028_013, w_047_102);
  not1 I047_100(w_047_101, w_047_095);
  and2 I047_101(w_047_105, w_032_004, w_047_103);
  or2  I048_024(w_048_024, w_033_018, w_045_045);
  and2 I048_035(w_048_035, w_007_003, w_013_000);
  nand2 I048_036(w_048_036, w_040_006, w_027_033);
  not1 I048_040(w_048_040, w_037_058);
  and2 I048_043(w_047_099, w_030_006, w_047_088);
  nand2 I049_001(w_049_001, w_046_035, w_030_027);
  or2  I049_002(w_049_002, w_020_002, w_041_025);
  or2  I049_005(w_049_005, w_047_099, w_042_000);
  not1 I050_001(w_050_001, w_041_033);
  and2 I050_009(w_050_009, w_044_014, w_031_007);
  and2 I051_000(w_051_000, w_021_037, w_031_009);
  nand2 I051_008(w_051_008, w_027_043, w_033_023);
  nand2 I052_009(w_052_009, w_001_029, w_013_000);
  or2  I052_011(w_052_011, w_042_020, w_046_013);
  not1 I052_041(w_052_041, w_038_029);
  not1 I052_042(w_052_044, w_052_043);
  nand2 I052_043(w_052_045, w_039_032, w_052_044);
  and2 I052_044(w_052_046, w_052_045, w_007_000);
  and2 I052_045(w_052_047, w_044_050, w_052_046);
  nand2 I052_046(w_052_048, w_052_047, w_033_066);
  not1 I052_047(w_052_043, w_052_048);
  or2  I053_002(w_053_002, w_052_041, w_014_006);
  or2  I053_004(w_053_004, w_000_069, w_025_052);
  nand2 I053_016(w_053_016, w_041_007, w_043_063);
  not1 I053_019(w_053_019, w_052_009);
  nand2 I053_023(w_053_023, w_024_022, w_026_025);
  and2 I053_062(w_053_062, w_019_004, w_048_024);
  and2 I054_003(w_054_003, w_000_083, w_018_019);
  not1 I054_004(w_054_004, w_020_002);
  or2  I054_011(w_054_011, w_020_006, w_018_013);
  and2 I054_013(w_054_013, w_002_038, w_050_009);
  nand2 I054_018(w_054_018, w_040_005, w_053_023);
  and2 I054_020(w_054_020, w_044_015, w_006_000);
  and2 I055_009(w_055_009, w_041_014, w_020_009);
  nand2 I055_017(w_055_017, w_002_040, w_014_008);
  and2 I055_049(w_055_049, w_053_002, w_009_012);
  not1 I056_000(w_056_000, w_044_016);
  and2 I056_003(w_056_003, w_026_031, w_054_020);
  not1 I056_042(w_056_042, w_033_050);
  not1 I057_008(w_057_008, w_041_035);
  and2 I057_009(w_057_009, w_055_049, w_043_058);
  or2  I057_012(w_057_012, w_000_010, w_017_016);
  nand2 I058_005(w_058_005, w_022_023, w_034_012);
  not1 I058_014(w_058_014, w_033_066);
  or2  I058_054(w_058_054, w_049_005, w_049_002);
  and2 I058_061(w_058_061, w_042_030, w_018_003);
  nand2 I059_032(w_059_032, w_043_008, w_017_021);
  or2  I060_002(w_060_002, w_056_042, w_032_002);
  not1 I060_011(w_060_011, w_051_000);
  nand2 I061_005(w_061_005, w_054_003, w_048_036);
  not1 I061_045(w_061_045, w_021_003);
  and2 I062_000(w_062_000, w_011_016, w_019_008);
  nand2 I062_001(w_062_001, w_024_002, w_033_013);
  and2 I062_002(w_062_002, w_050_001, w_061_005);
  and2 I062_003(w_062_005, w_062_004, w_028_015);
  not1 I062_004(w_062_006, w_062_005);
  nand2 I062_005(w_062_007, w_028_009, w_062_006);
  or2  I062_006(w_062_008, w_041_030, w_062_007);
  and2 I062_007(w_062_009, w_062_008, w_059_032);
  or2  I062_008(w_062_010, w_056_000, w_062_009);
  or2  I062_009(w_062_011, w_062_010, w_009_002);
  and2 I062_010(w_062_012, w_031_022, w_062_011);
  not1 I062_011(w_062_004, w_062_012);
  and2 I063_023(w_063_023, w_026_058, w_062_000);
  and2 I063_028(w_063_028, w_043_023, w_053_004);
  nand2 I064_040(w_064_040, w_046_004, w_053_016);
  nand2 I065_024(w_065_024, w_008_000, w_054_011);
  not1 I065_059(w_065_059, w_020_006);
  nand2 I066_013(w_066_013, w_009_001, w_023_041);
  not1 I068_006(w_068_006, w_050_009);
  nand2 I068_007(w_068_007, w_044_010, w_026_038);
  not1 I069_006(w_069_006, w_017_017);
  and2 I069_009(w_069_009, w_043_040, w_054_018);
  or2  I069_043(w_069_043, w_055_017, w_015_000);
  nand2 I069_068(w_069_068, w_037_067, w_029_078);
  not1 I070_006(w_070_006, w_038_038);
  and2 I070_043(w_070_043, w_027_045, w_041_014);
  not1 I070_079(w_070_081, w_070_080);
  not1 I070_080(w_070_082, w_070_081);
  and2 I070_081(w_070_080, w_041_010, w_070_082);
  or2  I071_013(w_071_013, w_008_005, w_044_008);
  or2  I071_030(w_071_030, w_019_021, w_039_029);
  and2 I071_080(w_071_080, w_009_006, w_002_093);
  not1 I072_027(w_072_027, w_009_007);
  and2 I073_020(w_073_020, w_003_016, w_053_019);
  not1 I076_031(w_076_031, w_050_001);
  not1 I076_065(w_076_065, w_052_011);
  or2  I077_008(w_077_008, w_032_000, w_068_007);
  or2  I078_027(w_078_027, w_060_002, w_016_004);
  not1 I078_055(w_078_055, w_077_008);
  not1 I079_006(w_079_006, w_027_023);
  or2  I080_019(w_080_019, w_017_034, w_036_070);
  not1 I080_020(w_080_020, w_057_012);
  and2 I082_001(w_082_001, w_022_015, w_003_018);
  or2  I083_005(w_083_005, w_021_052, w_010_043);
  not1 I084_002(w_084_002, w_030_010);
  not1 I084_004(w_084_006, w_084_005);
  or2  I084_005(w_084_007, w_084_006, w_084_029);
  not1 I084_006(w_084_008, w_084_007);
  not1 I084_007(w_084_009, w_084_008);
  nand2 I084_008(w_084_010, w_084_009, w_011_025);
  nand2 I084_009(w_084_011, w_084_010, w_057_009);
  and2 I084_010(w_084_012, w_084_011, w_069_043);
  or2  I084_011(w_084_005, w_084_012, w_016_000);
  or2  I084_012(w_084_017, w_084_016, w_064_040);
  and2 I084_013(w_084_018, w_084_017, w_065_059);
  nand2 I084_014(w_084_019, w_005_016, w_084_018);
  and2 I084_015(w_084_020, w_058_061, w_084_019);
  and2 I084_016(w_084_021, w_039_004, w_084_020);
  and2 I084_017(w_084_022, w_084_021, w_017_030);
  nand2 I084_018(w_084_023, w_084_022, w_023_086);
  and2 I084_019(w_084_024, w_084_023, w_024_003);
  and2 I084_020(w_084_025, w_018_032, w_084_024);
  and2 I084_021(w_084_026, w_063_023, w_084_025);
  and2 I084_022(w_084_027, w_084_026, w_037_054);
  not1 I084_023(w_084_016, w_084_007);
  and2 I084_024(w_084_029, w_001_029, w_084_027);
  not1 I085_032(w_085_032, w_022_048);
  not1 I085_086(w_085_086, w_043_020);
  or2  I088_010(w_088_010, w_028_005, w_085_032);
  or2  I088_017(w_088_017, w_051_008, w_030_059);
  and2 I089_016(w_089_016, w_044_001, w_080_020);
  and2 I089_054(w_089_054, w_027_006, w_078_027);
  not1 I091_023(w_091_023, w_071_030);
  not1 I092_059(w_092_059, w_046_003);
  nand2 I093_010(w_093_010, w_083_005, w_055_009);
  nand2 I093_030(w_093_030, w_024_008, w_002_016);
  and2 I094_028(w_094_028, w_057_008, w_046_013);
  nand2 I094_033(w_094_033, w_003_021, w_066_013);
  nand2 I095_000(w_095_000, w_006_000, w_041_002);
  not1 I095_001(w_095_001, w_027_020);
  and2 I095_002(w_095_002, w_038_012, w_080_019);
  and2 I096_039(w_096_039, w_054_013, w_094_028);
  and2 I097_045(w_097_047, w_097_046, w_068_006);
  nand2 I097_046(w_097_048, w_097_047, w_092_059);
  or2  I097_047(w_097_049, w_097_048, w_047_029);
  or2  I097_048(w_097_050, w_097_049, w_071_013);
  or2  I097_049(w_097_046, w_097_050, w_072_027);
  not1 I098_002(w_098_002, w_035_006);
  not1 I100_000(w_100_000, w_065_024);
  nand2 I100_001(w_100_001, w_062_001, w_054_004);
  nand2 I100_002(w_100_002, w_035_007, w_007_000);
  or2  I100_003(w_100_003, w_088_017, w_058_014);
  and2 I100_004(w_100_004, w_039_036, w_095_002);
  not1 I100_005(w_100_005, w_062_000);
  not1 I100_006(w_100_006, w_073_020);
  and2 I100_007(w_100_007, w_032_002, w_029_009);
  not1 I100_008(w_100_008, w_043_016);
  and2 I100_009(w_100_009, w_089_016, w_035_000);
  nand2 I100_010(w_100_010, w_095_001, w_063_028);
  nand2 I100_011(w_100_011, w_014_008, w_031_050);
  and2 I100_012(w_100_012, w_028_011, w_098_002);
  not1 I100_013(w_100_013, w_071_080);
  nand2 I100_014(w_100_014, w_056_003, w_076_065);
  or2  I100_015(w_100_015, w_020_003, w_049_001);
  or2  I100_016(w_100_016, w_084_002, w_076_031);
  nand2 I100_017(w_100_017, w_039_002, w_047_005);
  and2 I100_018(w_100_018, w_078_055, w_032_001);
  and2 I100_019(w_100_019, w_082_001, w_058_054);
  or2  I100_020(w_100_020, w_053_062, w_040_005);
  nand2 I100_021(w_100_021, w_089_054, w_060_011);
  nand2 I100_022(w_100_022, w_062_002, w_037_038);
  not1 I100_023(w_100_023, w_093_030);
  not1 I100_024(w_100_024, w_040_000);
  not1 I100_025(w_100_025, w_070_043);
  nand2 I100_026(w_100_026, w_028_014, w_085_086);
  or2  I100_027(w_100_027, w_091_023, w_035_005);
  and2 I100_028(w_100_028, w_017_032, w_005_000);
  or2  I100_029(w_100_029, w_096_039, w_007_006);
  and2 I100_030(w_100_030, w_045_006, w_069_006);
  not1 I100_031(w_100_031, w_009_007);
  or2  I100_032(w_100_032, w_079_006, w_024_059);
  or2  I100_033(w_100_033, w_061_045, w_058_005);
  or2  I100_034(w_100_034, w_093_010, w_037_062);
  nand2 I100_035(w_100_035, w_094_033, w_088_010);
  and2 I100_036(w_100_036, w_095_000, w_048_040);
  or2  I100_037(w_100_037, w_069_068, w_048_035);
  nand2 I100_038(w_100_038, w_069_009, w_041_017);
  and2 I100_039(w_100_039, w_070_006, w_018_028);

  initial begin
    $get_module_info();
  end
endmodule

// ****** Combined Logic Module Defination ******

// ****** TestBench Module Defination ******

/*
module tb();
  wire  w_000_000, w_000_001, w_000_002, w_000_003, w_000_004, w_000_005, w_000_006, w_000_007, w_000_008, w_000_009, w_000_010, w_000_011, w_000_012, w_000_013, w_000_014, w_000_015, w_000_016, w_000_018, w_000_019, w_000_020, w_000_021, w_000_022, w_000_023, w_000_024, w_000_025, w_000_026, w_000_027, w_000_028, w_000_029, w_000_030, w_000_031, w_000_032, w_000_033, w_000_034, w_000_035, w_000_036, w_000_037, w_000_038, w_000_039, w_000_040, w_000_041, w_000_042, w_000_043, w_000_044, w_000_045, w_000_046, w_000_047, w_000_048, w_000_049, w_000_050, w_000_051, w_000_052, w_000_053, w_000_054, w_000_055, w_000_056, w_000_057, w_000_058, w_000_059, w_000_060, w_000_061, w_000_062, w_000_064, w_000_065, w_000_066, w_000_067, w_000_068, w_000_069, w_000_070, w_000_071, w_000_072, w_000_073, w_000_074, w_000_076, w_000_077, w_000_078, w_000_079, w_000_082, w_000_083, w_000_084, w_000_085, w_000_086, w_000_087, w_000_088, w_000_089, w_000_090, w_000_091, w_000_092, w_000_096, w_100_000, w_100_001, w_100_002, w_100_003, w_100_004, w_100_005, w_100_006, w_100_007, w_100_008, w_100_009, w_100_010, w_100_011, w_100_012, w_100_013, w_100_014, w_100_015, w_100_016, w_100_017, w_100_018, w_100_019, w_100_020, w_100_021, w_100_022, w_100_023, w_100_024, w_100_025, w_100_026, w_100_027, w_100_028, w_100_029, w_100_030, w_100_031, w_100_032, w_100_033, w_100_034, w_100_035, w_100_036, w_100_037, w_100_038, w_100_039 ;
  combLogic I0(  w_000_000, w_000_001, w_000_002, w_000_003, w_000_004, w_000_005, w_000_006, w_000_007, w_000_008, w_000_009, w_000_010, w_000_011, w_000_012, w_000_013, w_000_014, w_000_015, w_000_016, w_000_018, w_000_019, w_000_020, w_000_021, w_000_022, w_000_023, w_000_024, w_000_025, w_000_026, w_000_027, w_000_028, w_000_029, w_000_030, w_000_031, w_000_032, w_000_033, w_000_034, w_000_035, w_000_036, w_000_037, w_000_038, w_000_039, w_000_040, w_000_041, w_000_042, w_000_043, w_000_044, w_000_045, w_000_046, w_000_047, w_000_048, w_000_049, w_000_050, w_000_051, w_000_052, w_000_053, w_000_054, w_000_055, w_000_056, w_000_057, w_000_058, w_000_059, w_000_060, w_000_061, w_000_062, w_000_064, w_000_065, w_000_066, w_000_067, w_000_068, w_000_069, w_000_070, w_000_071, w_000_072, w_000_073, w_000_074, w_000_076, w_000_077, w_000_078, w_000_079, w_000_082, w_000_083, w_000_084, w_000_085, w_000_086, w_000_087, w_000_088, w_000_089, w_000_090, w_000_091, w_000_092, w_000_096, w_100_000, w_100_001, w_100_002, w_100_003, w_100_004, w_100_005, w_100_006, w_100_007, w_100_008, w_100_009, w_100_010, w_100_011, w_100_012, w_100_013, w_100_014, w_100_015, w_100_016, w_100_017, w_100_018, w_100_019, w_100_020, w_100_021, w_100_022, w_100_023, w_100_024, w_100_025, w_100_026, w_100_027, w_100_028, w_100_029, w_100_030, w_100_031, w_100_032, w_100_033, w_100_034, w_100_035, w_100_036, w_100_037, w_100_038, w_100_039  );

  reg r0, r1, r2, r3, r4, r5, r6, r7, r8, r9, r10, r11, r12, r13, r14, r15, r16, r17, r18, r19, r20, r21, r22, r23, r24, r25, r26, r27, r28, r29, r30, r31, r32, r33, r34, r35, r36, r37, r38, r39, r40, r41, r42, r43, r44, r45, r46, r47, r48, r49, r50, r51, r52, r53, r54, r55, r56, r57, r58, r59, r60, r61, r62, r63, r64, r65, r66, r67, r68, r69, r70, r71, r72, r73, r74, r75, r76, r77, r78, r79, r80, r81, r82, r83, r84, r85, r86, r87, r88, r89, r90, r91, r92, r93, r94, r95, r96, r97, r98, rEnd; 

  assign w_000_000 = r0;
  assign w_000_001 = r1;
  assign w_000_002 = r2;
  assign w_000_003 = r3;
  assign w_000_004 = r4;
  assign w_000_005 = r5;
  assign w_000_006 = r6;
  assign w_000_007 = r7;
  assign w_000_008 = r8;
  assign w_000_009 = r9;
  assign w_000_010 = r10;
  assign w_000_011 = r11;
  assign w_000_012 = r12;
  assign w_000_013 = r13;
  assign w_000_014 = r14;
  assign w_000_015 = r15;
  assign w_000_016 = r16;
  assign w_000_017 = r17;
  assign w_000_018 = r18;
  assign w_000_019 = r19;
  assign w_000_020 = r20;
  assign w_000_021 = r21;
  assign w_000_022 = r22;
  assign w_000_023 = r23;
  assign w_000_024 = r24;
  assign w_000_025 = r25;
  assign w_000_026 = r26;
  assign w_000_027 = r27;
  assign w_000_028 = r28;
  assign w_000_029 = r29;
  assign w_000_030 = r30;
  assign w_000_031 = r31;
  assign w_000_032 = r32;
  assign w_000_033 = r33;
  assign w_000_034 = r34;
  assign w_000_035 = r35;
  assign w_000_036 = r36;
  assign w_000_037 = r37;
  assign w_000_038 = r38;
  assign w_000_039 = r39;
  assign w_000_040 = r40;
  assign w_000_041 = r41;
  assign w_000_042 = r42;
  assign w_000_043 = r43;
  assign w_000_044 = r44;
  assign w_000_045 = r45;
  assign w_000_046 = r46;
  assign w_000_047 = r47;
  assign w_000_048 = r48;
  assign w_000_049 = r49;
  assign w_000_050 = r50;
  assign w_000_051 = r51;
  assign w_000_052 = r52;
  assign w_000_053 = r53;
  assign w_000_054 = r54;
  assign w_000_055 = r55;
  assign w_000_056 = r56;
  assign w_000_057 = r57;
  assign w_000_058 = r58;
  assign w_000_059 = r59;
  assign w_000_060 = r60;
  assign w_000_061 = r61;
  assign w_000_062 = r62;
  assign w_000_063 = r63;
  assign w_000_064 = r64;
  assign w_000_065 = r65;
  assign w_000_066 = r66;
  assign w_000_067 = r67;
  assign w_000_068 = r68;
  assign w_000_069 = r69;
  assign w_000_070 = r70;
  assign w_000_071 = r71;
  assign w_000_072 = r72;
  assign w_000_073 = r73;
  assign w_000_074 = r74;
  assign w_000_075 = r75;
  assign w_000_076 = r76;
  assign w_000_077 = r77;
  assign w_000_078 = r78;
  assign w_000_079 = r79;
  assign w_000_080 = r80;
  assign w_000_081 = r81;
  assign w_000_082 = r82;
  assign w_000_083 = r83;
  assign w_000_084 = r84;
  assign w_000_085 = r85;
  assign w_000_086 = r86;
  assign w_000_087 = r87;
  assign w_000_088 = r88;
  assign w_000_089 = r89;
  assign w_000_090 = r90;
  assign w_000_091 = r91;
  assign w_000_092 = r92;
  assign w_000_093 = r93;
  assign w_000_094 = r94;
  assign w_000_095 = r95;
  assign w_000_096 = r96;
  assign w_000_097 = r97;
  assign w_000_098 = r98;

  initial begin 
    r0 = 1'b0; 
    r1 = 1'b0; 
    r2 = 1'b0; 
    r3 = 1'b0; 
    r4 = 1'b0; 
    r5 = 1'b0; 
    r6 = 1'b0; 
    r7 = 1'b0; 
    r8 = 1'b0; 
    r9 = 1'b0; 
    r10 = 1'b0; 
    r11 = 1'b0; 
    r12 = 1'b0; 
    r13 = 1'b0; 
    r14 = 1'b0; 
    r15 = 1'b0; 
    r16 = 1'b0; 
    r17 = 1'b0; 
    r18 = 1'b0; 
    r19 = 1'b0; 
    r20 = 1'b0; 
    r21 = 1'b0; 
    r22 = 1'b0; 
    r23 = 1'b0; 
    r24 = 1'b0; 
    r25 = 1'b0; 
    r26 = 1'b0; 
    r27 = 1'b0; 
    r28 = 1'b0; 
    r29 = 1'b0; 
    r30 = 1'b0; 
    r31 = 1'b0; 
    r32 = 1'b0; 
    r33 = 1'b0; 
    r34 = 1'b0; 
    r35 = 1'b0; 
    r36 = 1'b0; 
    r37 = 1'b0; 
    r38 = 1'b0; 
    r39 = 1'b0; 
    r40 = 1'b0; 
    r41 = 1'b0; 
    r42 = 1'b0; 
    r43 = 1'b0; 
    r44 = 1'b0; 
    r45 = 1'b0; 
    r46 = 1'b0; 
    r47 = 1'b0; 
    r48 = 1'b0; 
    r49 = 1'b0; 
    r50 = 1'b0; 
    r51 = 1'b0; 
    r52 = 1'b0; 
    r53 = 1'b0; 
    r54 = 1'b0; 
    r55 = 1'b0; 
    r56 = 1'b0; 
    r57 = 1'b0; 
    r58 = 1'b0; 
    r59 = 1'b0; 
    r60 = 1'b0; 
    r61 = 1'b0; 
    r62 = 1'b0; 
    r63 = 1'b0; 
    r64 = 1'b0; 
    r65 = 1'b0; 
    r66 = 1'b0; 
    r67 = 1'b0; 
    r68 = 1'b0; 
    r69 = 1'b0; 
    r70 = 1'b0; 
    r71 = 1'b0; 
    r72 = 1'b0; 
    r73 = 1'b0; 
    r74 = 1'b0; 
    r75 = 1'b0; 
    r76 = 1'b0; 
    r77 = 1'b0; 
    r78 = 1'b0; 
    r79 = 1'b0; 
    r80 = 1'b0; 
    r81 = 1'b0; 
    r82 = 1'b0; 
    r83 = 1'b0; 
    r84 = 1'b0; 
    r85 = 1'b0; 
    r86 = 1'b0; 
    r87 = 1'b0; 
    r88 = 1'b0; 
    r89 = 1'b0; 
    r90 = 1'b0; 
    r91 = 1'b0; 
    r92 = 1'b0; 
    r93 = 1'b0; 
    r94 = 1'b0; 
    r95 = 1'b0; 
    r96 = 1'b0; 
    r97 = 1'b0; 
    r98 = 1'b0; 
    $monitor("%t %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b  ", $time, w_000_000, w_000_001, w_000_002, w_000_003, w_000_004, w_000_005, w_000_006, w_000_007, w_000_008, w_000_009, w_000_010, w_000_011, w_000_012, w_000_013, w_000_014, w_000_015, w_000_016, w_000_017, w_000_018, w_000_019, w_000_020, w_000_021, w_000_022, w_000_023, w_000_024, w_000_025, w_000_026, w_000_027, w_000_028, w_000_029, w_000_030, w_000_031, w_000_032, w_000_033, w_000_034, w_000_035, w_000_036, w_000_037, w_000_038, w_000_039, w_000_040, w_000_041, w_000_042, w_000_043, w_000_044, w_000_045, w_000_046, w_000_047, w_000_048, w_000_049, w_000_050, w_000_051, w_000_052, w_000_053, w_000_054, w_000_055, w_000_056, w_000_057, w_000_058, w_000_059, w_000_060, w_000_061, w_000_062, w_000_063, w_000_064, w_000_065, w_000_066, w_000_067, w_000_068, w_000_069, w_000_070, w_000_071, w_000_072, w_000_073, w_000_074, w_000_075, w_000_076, w_000_077, w_000_078, w_000_079, w_000_080, w_000_081, w_000_082, w_000_083, w_000_084, w_000_085, w_000_086, w_000_087, w_000_088, w_000_089, w_000_090, w_000_091, w_000_092, w_000_093, w_000_094, w_000_095, w_000_096, w_000_097, w_000_098, w_100_000, w_100_001, w_100_002, w_100_003, w_100_004, w_100_005, w_100_006, w_100_007, w_100_008, w_100_009, w_100_010, w_100_011, w_100_012, w_100_013, w_100_014, w_100_015, w_100_016, w_100_017, w_100_018, w_100_019, w_100_020, w_100_021, w_100_022, w_100_023, w_100_024, w_100_025, w_100_026, w_100_027, w_100_028, w_100_029, w_100_030, w_100_031, w_100_032, w_100_033, w_100_034, w_100_035, w_100_036, w_100_037, w_100_038, w_100_039);
    #100;
    $finish;
  end
  always #1 r0 = ~r0;
  always #2 r1 = ~r1;
  always #4 r2 = ~r2;
  always #8 r3 = ~r3;
  always #16 r4 = ~r4;
  always #32 r5 = ~r5;
  always #64 r6 = ~r6;
  always #128 r7 = ~r7;
  always #256 r8 = ~r8;
  always #512 r9 = ~r9;
  always #1024 r10 = ~r10;
  always #2048 r11 = ~r11;
  always #4096 r12 = ~r12;
  always #8192 r13 = ~r13;
  always #16384 r14 = ~r14;
  always #32768 r15 = ~r15;
  always #65536 r16 = ~r16;
  always #131072 r17 = ~r17;
  always #262144 r18 = ~r18;
  always #524288 r19 = ~r19;
  always #1048576 r20 = ~r20;
  always #2097152 r21 = ~r21;
  always #4194304 r22 = ~r22;
  always #8388608 r23 = ~r23;
  always #16777216 r24 = ~r24;
  always #33554432 r25 = ~r25;
  always #67108864 r26 = ~r26;
  always #134217728 r27 = ~r27;
  always #268435456 r28 = ~r28;
  always #536870912 r29 = ~r29;
  always #1073741824 r30 = ~r30;
  always #2147483648 r31 = ~r31;
  always #4294967296 r32 = ~r32;
  always #8589934592 r33 = ~r33;
  always #17179869184 r34 = ~r34;
  always #34359738368 r35 = ~r35;
  always #68719476736 r36 = ~r36;
  always #137438953472 r37 = ~r37;
  always #274877906944 r38 = ~r38;
  always #549755813888 r39 = ~r39;
  always #1099511627776 r40 = ~r40;
  always #2199023255552 r41 = ~r41;
  always #4398046511104 r42 = ~r42;
  always #8796093022208 r43 = ~r43;
  always #17592186044416 r44 = ~r44;
  always #35184372088832 r45 = ~r45;
  always #70368744177664 r46 = ~r46;
  always #140737488355328 r47 = ~r47;
  always #281474976710656 r48 = ~r48;
  always #562949953421312 r49 = ~r49;
  always #1125899906842624 r50 = ~r50;
  always #2251799813685248 r51 = ~r51;
  always #4503599627370496 r52 = ~r52;
  always #9007199254740992 r53 = ~r53;
  always #18014398509481984 r54 = ~r54;
  always #36028797018963968 r55 = ~r55;
  always #72057594037927936 r56 = ~r56;
  always #144115188075855872 r57 = ~r57;
  always #288230376151711744 r58 = ~r58;
  always #576460752303423488 r59 = ~r59;
  always #1152921504606846976 r60 = ~r60;
  always #2305843009213693952 r61 = ~r61;
  always #4611686018427387904 r62 = ~r62;
  always #9223372036854775808 r63 = ~r63;
  always #1 r64 = ~r64;
  always #2 r65 = ~r65;
  always #4 r66 = ~r66;
  always #8 r67 = ~r67;
  always #16 r68 = ~r68;
  always #32 r69 = ~r69;
  always #64 r70 = ~r70;
  always #128 r71 = ~r71;
  always #256 r72 = ~r72;
  always #512 r73 = ~r73;
  always #1024 r74 = ~r74;
  always #2048 r75 = ~r75;
  always #4096 r76 = ~r76;
  always #8192 r77 = ~r77;
  always #16384 r78 = ~r78;
  always #32768 r79 = ~r79;
  always #65536 r80 = ~r80;
  always #131072 r81 = ~r81;
  always #262144 r82 = ~r82;
  always #524288 r83 = ~r83;
  always #1048576 r84 = ~r84;
  always #2097152 r85 = ~r85;
  always #4194304 r86 = ~r86;
  always #8388608 r87 = ~r87;
  always #16777216 r88 = ~r88;
  always #33554432 r89 = ~r89;
  always #67108864 r90 = ~r90;
  always #134217728 r91 = ~r91;
  always #268435456 r92 = ~r92;
  always #536870912 r93 = ~r93;
  always #1073741824 r94 = ~r94;
  always #2147483648 r95 = ~r95;
  always #4294967296 r96 = ~r96;
  always #8589934592 r97 = ~r97;
  always #17179869184 r98 = ~r98;
endmodule
*/
// ****** TestBench Module Defination End ******

/*
// ******* The results for this case *********
******* result_1.txt *********
1)
  Loop Signals: w_012_052, w_012_053, w_012_054, w_012_055, 
  Loop Gates: I012_051.port1, I012_052.port1, I012_053.port1, I012_054.port1, 

2)
  Loop Signals: w_012_055, w_012_059, w_012_060, w_012_061, w_012_062, w_012_063, w_012_064, w_012_065, w_012_067, 
  Loop Gates: I012_053.port2, I012_055.port1, I012_056.port1, I012_057.port1, I012_058.port1, I012_059.port1, I012_060.port1, I012_061.port1, I012_062.port2, 

3)
  Loop Signals: w_005_002, w_005_003, w_005_004, w_005_005, 
  Loop Gates: I005_001.port2, I005_002.port1, I005_003.port1, I005_004.port2, 

4)
  Loop Signals: w_005_004, w_005_009, w_005_010, w_005_011, w_005_012, w_005_013, w_005_014, w_005_015, w_005_016, w_005_018, 
  Loop Gates: I005_002.port2, I005_005.port1, I005_006.port2, I005_007.port2, I005_008.port1, I005_009.port1, I005_010.port1, I005_011.port2, I005_012.port1, I005_013.port2, 

5)
  Loop Signals: w_062_004, w_062_005, w_062_006, w_062_007, w_062_008, w_062_009, w_062_010, w_062_011, w_062_012, 
  Loop Gates: I062_003.port1, I062_004.port1, I062_005.port2, I062_006.port2, I062_007.port1, I062_008.port2, I062_009.port1, I062_010.port2, I062_011.port1, 

6)
  Loop Signals: w_070_080, w_070_081, w_070_082, 
  Loop Gates: I070_079.port1, I070_080.port1, I070_081.port2, 

7)
  Loop Signals: w_020_011, w_020_012, w_020_013, w_020_014, w_020_015, w_020_016, w_020_017, w_020_018, w_020_019, w_020_020, 
  Loop Gates: I020_010.port2, I020_011.port1, I020_012.port1, I020_013.port2, I020_014.port2, I020_015.port1, I020_016.port2, I020_017.port2, I020_018.port2, I020_019.port2, 

8)
  Loop Signals: w_097_046, w_097_047, w_097_048, w_097_049, w_097_050, 
  Loop Gates: I097_045.port1, I097_046.port1, I097_047.port1, I097_048.port1, I097_049.port1, 

9)
  Loop Signals: w_032_004, w_032_005, w_032_006, w_032_007, w_032_008, w_032_009, 
  Loop Gates: I032_003.port2, I032_004.port1, I032_005.port1, I032_006.port2, I032_007.port1, I032_008.port1, 

10)
  Loop Signals: w_032_007, w_032_013, w_032_014, w_032_015, w_032_016, w_032_018, 
  Loop Gates: I032_005.port2, I032_009.port1, I032_010.port1, I032_011.port1, I032_012.port1, I032_013.port2, 

11)
  Loop Signals: w_052_043, w_052_044, w_052_045, w_052_046, w_052_047, w_052_048, 
  Loop Gates: I052_042.port1, I052_043.port2, I052_044.port1, I052_045.port2, I052_046.port1, I052_047.port1, 

12)
  Loop Signals: w_046_037, w_046_038, w_046_039, 
  Loop Gates: I046_036.port1, I046_037.port1, I046_038.port2, 

13)
  Loop Signals: w_046_037, w_046_043, w_046_044, w_046_045, w_046_046, w_046_047, w_046_048, w_046_050, 
  Loop Gates: I046_038.port1, I046_039.port1, I046_040.port2, I046_041.port1, I046_042.port1, I046_043.port1, I046_044.port1, I046_045.port2, 

14)
  Loop Signals: w_023_069, w_023_070, w_023_071, w_023_072, w_023_073, w_023_074, w_023_075, 
  Loop Gates: I023_068.port2, I023_069.port1, I023_070.port1, I023_071.port1, I023_072.port1, I023_073.port1, I023_074.port1, 

15)
  Loop Signals: w_023_072, w_023_079, w_023_080, w_023_081, w_023_082, w_023_083, w_023_084, w_023_085, w_023_086, w_023_087, w_023_088, w_023_089, w_023_090, w_023_092, 
  Loop Gates: I023_070.port2, I023_075.port1, I023_076.port2, I023_077.port2, I023_078.port1, I023_079.port2, I023_080.port2, I023_081.port2, I023_082.port1, I023_083.port2, I023_084.port1, I023_085.port1, I023_086.port1, I023_087.port2, 

16)
  Loop Signals: w_047_088, w_047_089, w_047_090, w_047_091, w_047_092, w_047_093, w_047_094, w_047_095, w_047_096, w_047_097, 
  Loop Gates: I047_088.port2, I047_089.port1, I047_090.port1, I047_091.port1, I047_092.port1, I047_093.port2, I047_094.port2, I047_095.port2, I047_096.port1, I047_097.port1, 

17)
  Loop Signals: w_047_095, w_047_101, w_047_102, w_047_103, w_047_105, 
  Loop Gates: I047_094.port1, I047_098.port1, I047_099.port2, I047_100.port1, I047_101.port2, 

18)
  Loop Signals: w_084_005, w_084_006, w_084_007, w_084_008, w_084_009, w_084_010, w_084_011, w_084_012, 
  Loop Gates: I084_004.port1, I084_005.port1, I084_006.port1, I084_007.port1, I084_008.port1, I084_009.port1, I084_010.port1, I084_011.port1, 

19)
  Loop Signals: w_084_007, w_084_016, w_084_017, w_084_018, w_084_019, w_084_020, w_084_021, w_084_022, w_084_023, w_084_024, w_084_025, w_084_026, w_084_027, w_084_029, 
  Loop Gates: I084_005.port2, I084_012.port1, I084_013.port1, I084_014.port2, I084_015.port2, I084_016.port2, I084_017.port1, I084_018.port1, I084_019.port1, I084_020.port2, I084_021.port2, I084_022.port1, I084_023.port1, I084_024.port2, 

20)
  Loop Signals: w_004_036, w_004_037, w_004_038, 
  Loop Gates: I004_035.port1, I004_036.port1, I004_037.port1, 

******* result_2.txt *********
1)
  Loop Signals: w_005_004, w_005_009, w_005_010, w_005_011, w_005_012, w_005_013, w_005_014, w_005_015, w_005_016, w_005_018, 
  Loop Gates: I005_002.port2, I005_005.port1, I005_006.port2, I005_007.port2, I005_008.port1, I005_009.port1, I005_010.port1, I005_011.port2, I005_012.port1, I005_013.port2, 

2)
  Loop Signals: w_070_080, w_070_081, w_070_082, 
  Loop Gates: I070_079.port1, I070_080.port1, I070_081.port2, 

3)
  Loop Signals: w_032_004, w_032_005, w_032_006, w_032_007, w_032_008, w_032_009, 
  Loop Gates: I032_003.port2, I032_004.port1, I032_005.port1, I032_006.port2, I032_007.port1, I032_008.port1, 

4)
  Loop Signals: w_032_007, w_032_013, w_032_014, w_032_015, w_032_016, w_032_018, 
  Loop Gates: I032_005.port2, I032_009.port1, I032_010.port1, I032_011.port1, I032_012.port1, I032_013.port2, 

5)
  Loop Signals: w_052_043, w_052_044, w_052_045, w_052_046, w_052_047, w_052_048, 
  Loop Gates: I052_042.port1, I052_043.port2, I052_044.port1, I052_045.port2, I052_046.port1, I052_047.port1, 

6)
  Loop Signals: w_046_037, w_046_043, w_046_044, w_046_045, w_046_046, w_046_047, w_046_048, w_046_050, 
  Loop Gates: I046_038.port1, I046_039.port1, I046_040.port2, I046_041.port1, I046_042.port1, I046_043.port1, I046_044.port1, I046_045.port2, 

7)
  Loop Signals: w_023_069, w_023_070, w_023_071, w_023_072, w_023_073, w_023_074, w_023_075, 
  Loop Gates: I023_068.port2, I023_069.port1, I023_070.port1, I023_071.port1, I023_072.port1, I023_073.port1, I023_074.port1, 

8)
  Loop Signals: w_047_088, w_047_089, w_047_090, w_047_091, w_047_092, w_047_093, w_047_094, w_047_095, w_047_096, w_047_097, 
  Loop Gates: I047_088.port2, I047_089.port1, I047_090.port1, I047_091.port1, I047_092.port1, I047_093.port2, I047_094.port2, I047_095.port2, I047_096.port1, I047_097.port1, 

9)
  Loop Signals: w_047_095, w_047_101, w_047_102, w_047_103, w_047_105, 
  Loop Gates: I047_094.port1, I047_098.port1, I047_099.port2, I047_100.port1, I047_101.port2, 

10)
  Loop Signals: w_004_036, w_004_037, w_004_038, 
  Loop Gates: I004_035.port1, I004_036.port1, I004_037.port1, 

******* result_3.txt *********
1)
  Loop Signals: w_012_052, w_012_053, w_012_054, w_012_055, 
  Loop Gates: I012_051.port1, I012_052.port1, I012_053.port1, I012_054.port1, 
  Loop Conditions: I012_053.port2=1, 
  (Signal Values: w_012_067=1, )

2)
  Loop Signals: w_012_055, w_012_059, w_012_060, w_012_061, w_012_062, w_012_063, w_012_064, w_012_065, w_012_067, 
  Loop Gates: I012_053.port2, I012_055.port1, I012_056.port1, I012_057.port1, I012_058.port1, I012_059.port1, I012_060.port1, I012_061.port1, I012_062.port2, 
  Loop Conditions: I012_053.port2=1, I012_057.port2=1, I012_058.port2=1, I012_060.port2=1, I012_062.port2=1, 
  (Signal Values: w_003_007=1, w_004_019=1, w_008_028=1, w_012_065=1, w_012_067=1, )

3)
  Loop Signals: w_005_002, w_005_003, w_005_004, w_005_005, 
  Loop Gates: I005_001.port2, I005_002.port1, I005_003.port1, I005_004.port2, 
  Loop Conditions: I005_001.port1=1, I005_002.port2=0, I005_004.port1=1, 
  (Signal Values: w_004_005=1, w_004_028=1, w_005_018=0, )

4)
  Loop Signals: w_062_004, w_062_005, w_062_006, w_062_007, w_062_008, w_062_009, w_062_010, w_062_011, w_062_012, 
  Loop Gates: I062_003.port1, I062_004.port1, I062_005.port2, I062_006.port2, I062_007.port1, I062_008.port2, I062_009.port1, I062_010.port2, I062_011.port1, 
  Loop Conditions: I062_003.port2=1, I062_005.port1=1, I062_006.port1=0, I062_007.port2=1, I062_008.port1=0, I062_009.port2=0, I062_010.port1=1, 
  (Signal Values: w_009_002=0, w_028_015=1, w_028_009=1, w_031_022=1, w_041_030=0, w_056_000=0, w_059_032=1, )

5)
  Loop Signals: w_020_011, w_020_012, w_020_013, w_020_014, w_020_015, w_020_016, w_020_017, w_020_018, w_020_019, w_020_020, 
  Loop Gates: I020_010.port2, I020_011.port1, I020_012.port1, I020_013.port2, I020_014.port2, I020_015.port1, I020_016.port2, I020_017.port2, I020_018.port2, I020_019.port2, 
  Loop Conditions: I020_010.port1=1, I020_011.port2=0, I020_013.port1=1, I020_014.port1=1, I020_016.port1=1, I020_017.port1=0, I020_018.port1=0, I020_019.port1=0, 
  (Signal Values: w_007_007=0, w_008_001=0, w_008_075=1, w_016_000=1, w_016_004=1, w_019_002=1, w_019_007=0, w_019_019=0, )

6)
  Loop Signals: w_097_046, w_097_047, w_097_048, w_097_049, w_097_050, 
  Loop Gates: I097_045.port1, I097_046.port1, I097_047.port1, I097_048.port1, I097_049.port1, 
  Loop Conditions: I097_045.port2=1, I097_046.port2=1, I097_047.port2=0, I097_048.port2=0, I097_049.port2=0, 
  (Signal Values: w_047_029=0, w_068_006=1, w_071_013=0, w_072_027=0, w_092_059=1, )

7)
  Loop Signals: w_046_037, w_046_038, w_046_039, 
  Loop Gates: I046_036.port1, I046_037.port1, I046_038.port2, 
  Loop Conditions: I046_037.port2=1, I046_038.port2=1, 
  (Signal Values: w_011_050=1, w_046_039=1, )

8)
  Loop Signals: w_023_072, w_023_079, w_023_080, w_023_081, w_023_082, w_023_083, w_023_084, w_023_085, w_023_086, w_023_087, w_023_088, w_023_089, w_023_090, w_023_092, 
  Loop Gates: I023_070.port2, I023_075.port1, I023_076.port2, I023_077.port2, I023_078.port1, I023_079.port2, I023_080.port2, I023_081.port2, I023_082.port1, I023_083.port2, I023_084.port1, I023_085.port1, I023_086.port1, I023_087.port2, 
  Loop Conditions: I023_070.port2=1, I023_076.port1=1, I023_077.port1=1, I023_078.port2=0, I023_079.port1=0, I023_080.port1=0, I023_081.port1=1, I023_082.port2=0, I023_083.port1=1, I023_084.port2=1, I023_087.port2=1, 
  (Signal Values: w_001_003=1, w_001_031=0, w_002_066=0, w_006_000=1, w_010_063=0, w_012_065=0, w_014_024=1, w_016_004=1, w_005_007=1, w_023_090=1, w_023_092=1, )

9)
  Loop Signals: w_084_005, w_084_006, w_084_007, w_084_008, w_084_009, w_084_010, w_084_011, w_084_012, 
  Loop Gates: I084_004.port1, I084_005.port1, I084_006.port1, I084_007.port1, I084_008.port1, I084_009.port1, I084_010.port1, I084_011.port1, 
  Loop Conditions: I084_005.port2=0, I084_008.port2=1, I084_009.port2=1, I084_010.port2=1, I084_011.port2=0, 
  (Signal Values: w_011_025=1, w_016_000=0, w_057_009=1, w_069_043=1, w_084_029=0, )

10)
  Loop Signals: w_084_007, w_084_016, w_084_017, w_084_018, w_084_019, w_084_020, w_084_021, w_084_022, w_084_023, w_084_024, w_084_025, w_084_026, w_084_027, w_084_029, 
  Loop Gates: I084_005.port2, I084_012.port1, I084_013.port1, I084_014.port2, I084_015.port2, I084_016.port2, I084_017.port1, I084_018.port1, I084_019.port1, I084_020.port2, I084_021.port2, I084_022.port1, I084_023.port1, I084_024.port2, 
  Loop Conditions: I084_005.port2=0, I084_012.port2=0, I084_013.port2=1, I084_014.port1=1, I084_015.port1=1, I084_016.port1=1, I084_017.port2=1, I084_018.port2=1, I084_019.port2=1, I084_020.port1=1, I084_021.port1=1, I084_022.port2=1, I084_024.port2=1, 
  (Signal Values: w_017_030=1, w_018_032=1, w_024_003=1, w_037_054=1, w_039_004=1, w_058_061=1, w_063_023=1, w_064_040=0, w_065_059=1, w_005_016=1, w_023_086=1, w_084_027=1, w_084_029=0, )

******* result_4.txt *********
1)
  Loop Breaker: I012_053.port0-w_012_055-Register-w_012_055'-I012_054.port1 

2)
  Loop Breaker: I012_053.port0-w_012_055-Register-w_012_055'-I012_061.port1 

3)
  Loop Breaker: I005_002.port0-w_005_004-Register-w_005_004'-I005_003.port1 

4)
  Loop Breaker: I062_003.port0-w_062_005-Register-w_062_005'-I062_004.port1 

5)
  Loop Breaker: I020_010.port0-w_020_012-Register-w_020_012'-I020_011.port1 

6)
  Loop Breaker: I097_045.port0-w_097_047-Register-w_097_047'-I097_046.port1 

7)
  Loop Breaker: I046_038.port0-w_046_037-Register-w_046_037'-I046_036.port1 

8)
  Loop Breaker: I023_070.port0-w_023_072-Register-w_023_072'-I023_086.port1 

9)
  Loop Breaker: I084_005.port0-w_084_007-Register-w_084_007'-I084_006.port1 

10)
  Loop Breaker: I084_005.port0-w_084_007-Register-w_084_007'-I084_023.port1 

// ******* The results for this case End *********
*/

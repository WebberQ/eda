// ****** Basic Gate Module Defination ******
module or2(out, in1, in2);
  output out;
  input in1, in2;
  wire in1, in2, out;
  assign out = in1 || in2;
endmodule

module and2(out, in1, in2);
  output out;
  input in1, in2;
  wire in1, in2, out;
  assign out = in1 && in2;
endmodule

module not1(out, in);
  output out;
  input in;
  wire in,out;
  assign out = ~in;
endmodule

module nand2(out, in1, in2);
  output out;
  input in1, in2;
  wire in1, in2, out;
  assign out = ~(in1 && in2);
endmodule
// ****** Basic Gate Module Defination End ******

// ****** Combined Logic Module Defination ******
module combLogic( w_000_000, w_000_001, w_000_002, w_000_003, w_000_004, w_000_005, w_000_006, w_000_007, w_000_008, w_000_009, w_000_010, w_000_011, w_000_012, w_000_013, w_000_014, w_000_015, w_000_016, w_000_017, w_000_018, w_000_019, w_000_020, w_000_021, w_000_022, w_000_023, w_000_024, w_000_025, w_000_026, w_000_027, w_000_028, w_000_029, w_000_030, w_000_031, w_000_032, w_000_033, w_000_034, w_000_035, w_000_036, w_000_037, w_000_038, w_000_039, w_000_040, w_000_041, w_000_042, w_000_043, w_000_044, w_000_045, w_000_046, w_000_047, w_000_048, w_000_049, w_000_050, w_000_051, w_000_052, w_000_053, w_000_054, w_000_055, w_000_056, w_000_057, w_000_058, w_000_059, w_000_060, w_000_061, w_000_062, w_000_063, w_000_064, w_000_065, w_000_066, w_000_067, w_000_068, w_000_069, w_000_070, w_000_071, w_000_072, w_000_073, w_000_074, w_000_075, w_000_076, w_000_077, w_000_078, w_000_079, w_000_080, w_000_081, w_000_082, w_000_083, w_000_084, w_000_085, w_000_086, w_000_087, w_000_088, w_000_089, w_000_090, w_000_091, w_000_092, w_000_093, w_000_094, w_000_095, w_000_096, w_000_097, w_000_098, w_000_099, w_000_100, w_000_101, w_000_102, w_000_103, w_000_104, w_000_105, w_000_106, w_000_107, w_000_108, w_000_109, w_000_110, w_000_111, w_000_112, w_000_113, w_000_114, w_000_115, w_000_116, w_000_117, w_000_118, w_000_119, w_000_120, w_000_121, w_000_122, w_000_123, w_000_124, w_000_125, w_000_126, w_000_127, w_000_128, w_000_129, w_000_130, w_000_131, w_000_132, w_000_133, w_000_134, w_000_135, w_000_136, w_000_137, w_000_138, w_000_139, w_000_140, w_000_141, w_000_142, w_000_143, w_000_144, w_000_145, w_000_146, w_000_147, w_000_148, w_000_149, w_000_150, w_000_151, w_000_152, w_000_153, w_000_154, w_000_155, w_000_156, w_000_157, w_000_158, w_000_159, w_000_160, w_000_161, w_000_162, w_000_163, w_000_164, w_000_165, w_000_166, w_000_167, w_000_169, w_000_170, w_000_171, w_000_172, w_000_173, w_000_174, w_000_175, w_000_176, w_000_177, w_000_178, w_000_179, w_000_180, w_000_181, w_000_182, w_000_183, w_000_184, w_000_185, w_000_186, w_000_187, w_000_188, w_000_189, w_000_190, w_000_191, w_000_192, w_000_193, w_000_194, w_000_195, w_000_196, w_000_197, w_000_198, w_000_199, w_000_200, w_000_202, w_000_203, w_000_204, w_000_205, w_000_206, w_000_207, w_000_208, w_000_209, w_000_210, w_000_211, w_000_212, w_000_213, w_000_214, w_000_215, w_000_216, w_000_217, w_000_218, w_000_219, w_000_220, w_000_221, w_000_222, w_000_223, w_000_224, w_000_225, w_000_226, w_000_227, w_000_228, w_000_229, w_000_230, w_000_231, w_000_232, w_000_233, w_000_234, w_000_235, w_000_236, w_000_237, w_000_238, w_000_239, w_000_240, w_000_241, w_000_242, w_000_243, w_000_244, w_000_245, w_000_246, w_000_247, w_000_248, w_000_249, w_000_250, w_000_251, w_000_252, w_000_253, w_000_254, w_000_255, w_000_256, w_000_257, w_000_258, w_000_259, w_000_260, w_000_261, w_000_262, w_000_263, w_000_264, w_000_265, w_000_266, w_000_267, w_000_268, w_000_269, w_000_270, w_000_271, w_000_272, w_000_273, w_000_274, w_000_275, w_000_276, w_000_277, w_000_278, w_000_279, w_000_280, w_000_281, w_000_282, w_000_283, w_000_284, w_000_285, w_000_286, w_000_287, w_000_288, w_000_289, w_000_290, w_000_291, w_000_292, w_000_293, w_000_294, w_000_295, w_000_296, w_000_297, w_000_298, w_000_299, w_000_300, w_000_301, w_000_302, w_000_303, w_000_304, w_000_305, w_000_306, w_000_307, w_000_308, w_000_309, w_000_310, w_000_311, w_000_312, w_000_313, w_000_314, w_000_315, w_000_316, w_000_317, w_000_318, w_000_319, w_000_320, w_000_321, w_000_322, w_000_323, w_000_324, w_000_325, w_000_326, w_000_327, w_000_328, w_000_329, w_000_330, w_000_331, w_000_332, w_000_333, w_000_334, w_000_335, w_000_336, w_000_337, w_000_338, w_000_339, w_000_340, w_000_341, w_000_342, w_000_343, w_000_344, w_000_345, w_000_346, w_000_347, w_000_348, w_000_349, w_000_350, w_000_351, w_000_352, w_000_353, w_000_354, w_000_355, w_000_356, w_000_357, w_000_358, w_000_359, w_000_360, w_000_361, w_000_362, w_000_363, w_000_364, w_000_365, w_000_366, w_000_367, w_000_368, w_000_370, w_000_371, w_000_372, w_000_373, w_000_374, w_000_375, w_000_376, w_000_377, w_000_378, w_000_379, w_000_380, w_000_381, w_000_382, w_000_383, w_000_384, w_000_385, w_000_386, w_000_387, w_000_388, w_000_389, w_000_390, w_000_391, w_000_392, w_000_393, w_000_394, w_000_395, w_000_396, w_000_397, w_000_398, w_000_399, w_000_400, w_000_401, w_000_402, w_000_403, w_000_404, w_000_405, w_000_406, w_000_408, w_000_409, w_000_410, w_000_411, w_000_412, w_000_413, w_000_414, w_000_415, w_000_416, w_000_417, w_000_418, w_000_419, w_000_420, w_000_421, w_000_422, w_000_423, w_000_424, w_000_425, w_000_426, w_000_427, w_000_428, w_000_429, w_000_430, w_000_431, w_000_432, w_000_433, w_000_434, w_000_435, w_000_436, w_000_437, w_000_438, w_000_439, w_000_440, w_000_441, w_000_442, w_000_443, w_000_444, w_000_445, w_000_446, w_000_447, w_000_448, w_000_449, w_000_450, w_000_451, w_000_452, w_000_453, w_000_454, w_000_455, w_000_456, w_000_457, w_000_458, w_000_459, w_000_460, w_000_461, w_000_462, w_000_463, w_000_464, w_000_465, w_000_466, w_000_467, w_000_468, w_000_469, w_000_470, w_000_471, w_000_472, w_000_473, w_000_474, w_000_475, w_000_476, w_000_477, w_000_478, w_000_479, w_000_480, w_000_481, w_000_482, w_000_483, w_000_484, w_000_485, w_000_486, w_000_487, w_000_488, w_000_489, w_000_490, w_000_491, w_000_492, w_000_493, w_000_494, w_000_495, w_000_496, w_000_497, w_000_498, w_000_499, w_000_500, w_000_501, w_000_502, w_000_503, w_000_504, w_000_505, w_000_506, w_000_507, w_000_508, w_000_510, w_000_511, w_000_512, w_000_513, w_000_514, w_000_515, w_000_516, w_000_517, w_000_518, w_000_519, w_000_520, w_000_521, w_000_522, w_000_523, w_000_524, w_000_525, w_000_526, w_000_527, w_000_528, w_000_529, w_000_530, w_000_531, w_000_532, w_000_533, w_000_534, w_000_535, w_000_536, w_000_537, w_000_538, w_000_540, w_000_541, w_000_542, w_000_543, w_000_544, w_000_545, w_000_546, w_000_547, w_000_548, w_000_549, w_000_550, w_000_551, w_000_552, w_000_553, w_000_554, w_000_555, w_000_556, w_000_557, w_000_558, w_000_559, w_000_560, w_000_561, w_000_563, w_000_564, w_000_565, w_000_566, w_000_567, w_000_568, w_000_569, w_000_570, w_000_571, w_000_572, w_000_573, w_000_574, w_000_575, w_000_576, w_000_577, w_000_578, w_000_579, w_000_580, w_000_581, w_000_582, w_000_583, w_000_584, w_000_585, w_000_586, w_000_587, w_000_588, w_000_589, w_000_590, w_000_591, w_000_592, w_000_593, w_000_594, w_000_595, w_000_596, w_000_597, w_000_598, w_000_599, w_000_600, w_000_601, w_000_602, w_000_603, w_000_604, w_000_605, w_000_606, w_000_607, w_000_608, w_000_609, w_000_610, w_000_611, w_000_612, w_000_613, w_000_614, w_000_615, w_000_616, w_000_617, w_000_618, w_000_619, w_000_620, w_000_621, w_000_622, w_000_623, w_000_624, w_000_625, w_000_626, w_000_627, w_000_628, w_000_629, w_000_630, w_000_632, w_000_634, w_000_635, w_000_636, w_000_637, w_000_638, w_000_639, w_000_640, w_000_641, w_000_642, w_000_643, w_000_644, w_000_645, w_000_646, w_000_647, w_000_648, w_000_649, w_000_650, w_000_651, w_000_652, w_000_653, w_000_654, w_000_655, w_000_656, w_000_657, w_000_658, w_000_659, w_000_660, w_000_661, w_000_662, w_000_663, w_000_664, w_000_665, w_000_666, w_000_667, w_000_668, w_000_671, w_000_674, w_000_675, w_000_676, w_000_679, w_000_680, w_000_681, w_000_682, w_000_683, w_000_684, w_000_685, w_000_687, w_000_688, w_000_689, w_000_690, w_000_691, w_000_692, w_000_693, w_000_694, w_000_695, w_000_696, w_000_697, w_000_698, w_000_699, w_000_701, w_000_702, w_000_703, w_000_704, w_000_705, w_000_706, w_000_707, w_000_708, w_000_709, w_000_710, w_000_711, w_000_712, w_000_713, w_000_714, w_000_715, w_000_716, w_000_717, w_000_718, w_000_720, w_000_722, w_000_724, w_000_725, w_000_726, w_000_727, w_000_728, w_000_731, w_000_732, w_000_733, w_000_734, w_000_735, w_000_736, w_000_738, w_000_739, w_000_740, w_000_741, w_000_743, w_000_744, w_000_745, w_000_747, w_000_748, w_000_749, w_000_751, w_000_754, w_000_756, w_000_757, w_000_758, w_000_759, w_000_762, w_000_763, w_000_768, w_000_770, w_000_772, w_000_776, w_000_777, w_000_780, w_000_783, w_800_000, w_800_001, w_800_002, w_800_003, w_800_004, w_800_005, w_800_006, w_800_007, w_800_008, w_800_009, w_800_010, w_800_011, w_800_012, w_800_013, w_800_014, w_800_015, w_800_016, w_800_017, w_800_018, w_800_019, w_800_020, w_800_021, w_800_022, w_800_023, w_800_024, w_800_025, w_800_026, w_800_027, w_800_028, w_800_029, w_800_030, w_800_031, w_800_032, w_800_033, w_800_034, w_800_035, w_800_036, w_800_037, w_800_038, w_800_039, w_800_040, w_800_041, w_800_042, w_800_043, w_800_044, w_800_045, w_800_046, w_800_047, w_800_048, w_800_049, w_800_050, w_800_051, w_800_052, w_800_053, w_800_054, w_800_055, w_800_056, w_800_057, w_800_058, w_800_059, w_800_060, w_800_061, w_800_062, w_800_063, w_800_064, w_800_065, w_800_066, w_800_067, w_800_068, w_800_069, w_800_070, w_800_071, w_800_072, w_800_073, w_800_074, w_800_075, w_800_076, w_800_077, w_800_078, w_800_079, w_800_080, w_800_081, w_800_082, w_800_083, w_800_084, w_800_085, w_800_086, w_800_087, w_800_088, w_800_089, w_800_090, w_800_091, w_800_092, w_800_093, w_800_094, w_800_095, w_800_096, w_800_097, w_800_098, w_800_099, w_800_100, w_800_101, w_800_102, w_800_103, w_800_104, w_800_105, w_800_106, w_800_107, w_800_108, w_800_109, w_800_110, w_800_111, w_800_112, w_800_113, w_800_114, w_800_115, w_800_116, w_800_117, w_800_118, w_800_119, w_800_120, w_800_121, w_800_122, w_800_123, w_800_124, w_800_125, w_800_126, w_800_127, w_800_128, w_800_129, w_800_130, w_800_131, w_800_132, w_800_133, w_800_134, w_800_135, w_800_136, w_800_137, w_800_138, w_800_139, w_800_140, w_800_141, w_800_142, w_800_143, w_800_144, w_800_145, w_800_146, w_800_147, w_800_148, w_800_149, w_800_150, w_800_151, w_800_152, w_800_153, w_800_154, w_800_155, w_800_156, w_800_157, w_800_158, w_800_159, w_800_160, w_800_161, w_800_162, w_800_163, w_800_164, w_800_165, w_800_166, w_800_167, w_800_168, w_800_169, w_800_170, w_800_171, w_800_172, w_800_173, w_800_174, w_800_175, w_800_176, w_800_177, w_800_178, w_800_179, w_800_180, w_800_181, w_800_182, w_800_183, w_800_184, w_800_185, w_800_186, w_800_187, w_800_188, w_800_189, w_800_190, w_800_191, w_800_192, w_800_193, w_800_194, w_800_195, w_800_196, w_800_197, w_800_198, w_800_199, w_800_200, w_800_201, w_800_202, w_800_203, w_800_204, w_800_205, w_800_206, w_800_207, w_800_208, w_800_209, w_800_210, w_800_211, w_800_212, w_800_213, w_800_214, w_800_215, w_800_216, w_800_217, w_800_218, w_800_219, w_800_220, w_800_221, w_800_222, w_800_223, w_800_224, w_800_225, w_800_226, w_800_227, w_800_228, w_800_229, w_800_230, w_800_231, w_800_232, w_800_233, w_800_234, w_800_235, w_800_236, w_800_237, w_800_238, w_800_239, w_800_240, w_800_241, w_800_242, w_800_243, w_800_244, w_800_245, w_800_246, w_800_247, w_800_248, w_800_249, w_800_250, w_800_251, w_800_252, w_800_253, w_800_254, w_800_255, w_800_256, w_800_257, w_800_258, w_800_259, w_800_260, w_800_261, w_800_262, w_800_263, w_800_264, w_800_265, w_800_266, w_800_267, w_800_268, w_800_269, w_800_270, w_800_271, w_800_272, w_800_273, w_800_274, w_800_275, w_800_276, w_800_277, w_800_278, w_800_279, w_800_280, w_800_281, w_800_282, w_800_283, w_800_284, w_800_285, w_800_286, w_800_287, w_800_288, w_800_289, w_800_290, w_800_291, w_800_292, w_800_293, w_800_294, w_800_295, w_800_296, w_800_297, w_800_298, w_800_299, w_800_300, w_800_301, w_800_302, w_800_303, w_800_304, w_800_305, w_800_306, w_800_307, w_800_308, w_800_309, w_800_310, w_800_311, w_800_312, w_800_313, w_800_314, w_800_315, w_800_316, w_800_317, w_800_318, w_800_319, w_800_320, w_800_321, w_800_322, w_800_323, w_800_324, w_800_325, w_800_326, w_800_327, w_800_328, w_800_329, w_800_330, w_800_331, w_800_332, w_800_333, w_800_334, w_800_335, w_800_336, w_800_337, w_800_338, w_800_339, w_800_340, w_800_341, w_800_342, w_800_343, w_800_344, w_800_345, w_800_346, w_800_347, w_800_348, w_800_349, w_800_350, w_800_351, w_800_352, w_800_353, w_800_354, w_800_355, w_800_356, w_800_357, w_800_358, w_800_359, w_800_360, w_800_361, w_800_362, w_800_363, w_800_364, w_800_365, w_800_366, w_800_367, w_800_368, w_800_369, w_800_370, w_800_371, w_800_372, w_800_373, w_800_374, w_800_375, w_800_376, w_800_377, w_800_378, w_800_379, w_800_380, w_800_381, w_800_382, w_800_383, w_800_384, w_800_385, w_800_386, w_800_387, w_800_388, w_800_389, w_800_390, w_800_391, w_800_392, w_800_393, w_800_394, w_800_395, w_800_396, w_800_397, w_800_398, w_800_399, w_800_400, w_800_401, w_800_402, w_800_403, w_800_404, w_800_405, w_800_406, w_800_407, w_800_408, w_800_409, w_800_410, w_800_411, w_800_412, w_800_413, w_800_414, w_800_415, w_800_416, w_800_417, w_800_418, w_800_419, w_800_420, w_800_421, w_800_422, w_800_423, w_800_424, w_800_425, w_800_426, w_800_427, w_800_428, w_800_429, w_800_430, w_800_431, w_800_432, w_800_433, w_800_434, w_800_435, w_800_436, w_800_437, w_800_438, w_800_439, w_800_440, w_800_441, w_800_442, w_800_443, w_800_444, w_800_445, w_800_446, w_800_447, w_800_448, w_800_449, w_800_450, w_800_451, w_800_452, w_800_453, w_800_454, w_800_455, w_800_456, w_800_457, w_800_458, w_800_459, w_800_460, w_800_461, w_800_462, w_800_463, w_800_464, w_800_465, w_800_466, w_800_467, w_800_468, w_800_469, w_800_470, w_800_471, w_800_472, w_800_473, w_800_474, w_800_475, w_800_476, w_800_477, w_800_478, w_800_479, w_800_480, w_800_481, w_800_482, w_800_483, w_800_484, w_800_485, w_800_486, w_800_487, w_800_488, w_800_489, w_800_490, w_800_491, w_800_492, w_800_493, w_800_494, w_800_495, w_800_496, w_800_497, w_800_498, w_800_499, w_800_500, w_800_501, w_800_502, w_800_503, w_800_504, w_800_505, w_800_506, w_800_507, w_800_508, w_800_509, w_800_510, w_800_511, w_800_512, w_800_513, w_800_514, w_800_515, w_800_516, w_800_517, w_800_518, w_800_519, w_800_520, w_800_521, w_800_522, w_800_523, w_800_524, w_800_525, w_800_526, w_800_527, w_800_528, w_800_529, w_800_530, w_800_531, w_800_532, w_800_533, w_800_534, w_800_535, w_800_536, w_800_537, w_800_538, w_800_539, w_800_540, w_800_541, w_800_542, w_800_543, w_800_544, w_800_545, w_800_546, w_800_547, w_800_548, w_800_549, w_800_550, w_800_551, w_800_552, w_800_553, w_800_554, w_800_555, w_800_556, w_800_557, w_800_558, w_800_559, w_800_560, w_800_561, w_800_562, w_800_563, w_800_564, w_800_565, w_800_566, w_800_567, w_800_568, w_800_569, w_800_570, w_800_571, w_800_572, w_800_573, w_800_574, w_800_575, w_800_576, w_800_577, w_800_578, w_800_579, w_800_580, w_800_581, w_800_582, w_800_583, w_800_584, w_800_585, w_800_586, w_800_587, w_800_588, w_800_589, w_800_590, w_800_591, w_800_592, w_800_593, w_800_594, w_800_595, w_800_596, w_800_597, w_800_598, w_800_599, w_800_600, w_800_601, w_800_602, w_800_603, w_800_604, w_800_605, w_800_606, w_800_607, w_800_608, w_800_609, w_800_610, w_800_611, w_800_612, w_800_613, w_800_614, w_800_615, w_800_616, w_800_617, w_800_618, w_800_619, w_800_620, w_800_621, w_800_622, w_800_623, w_800_624, w_800_625, w_800_626, w_800_627, w_800_628, w_800_629, w_800_630, w_800_631, w_800_632, w_800_633, w_800_634, w_800_635, w_800_636, w_800_637, w_800_638, w_800_639, w_800_640, w_800_641, w_800_642, w_800_643, w_800_644, w_800_645, w_800_646, w_800_647, w_800_648, w_800_649, w_800_650, w_800_651, w_800_652, w_800_653, w_800_654, w_800_655, w_800_656, w_800_657, w_800_658, w_800_659, w_800_660, w_800_661, w_800_662, w_800_663, w_800_664, w_800_665, w_800_666, w_800_667, w_800_668, w_800_669, w_800_670, w_800_671, w_800_672, w_800_673, w_800_674, w_800_675, w_800_676, w_800_677, w_800_678, w_800_679, w_800_680, w_800_681, w_800_682, w_800_683, w_800_684, w_800_685, w_800_686, w_800_687, w_800_688, w_800_689, w_800_690, w_800_691, w_800_692, w_800_693, w_800_694, w_800_695, w_800_696, w_800_697, w_800_698, w_800_699, w_800_700, w_800_701, w_800_702, w_800_703, w_800_704, w_800_705, w_800_706, w_800_707, w_800_708, w_800_709, w_800_710, w_800_711, w_800_712, w_800_713, w_800_714, w_800_715, w_800_716, w_800_717 );
  inout w_000_000, w_000_001, w_000_002, w_000_003, w_000_004, w_000_005, w_000_006, w_000_007, w_000_008, w_000_009, w_000_010, w_000_011, w_000_012, w_000_013, w_000_014, w_000_015, w_000_016, w_000_017, w_000_018, w_000_019, w_000_020, w_000_021, w_000_022, w_000_023, w_000_024, w_000_025, w_000_026, w_000_027, w_000_028, w_000_029, w_000_030, w_000_031, w_000_032, w_000_033, w_000_034, w_000_035, w_000_036, w_000_037, w_000_038, w_000_039, w_000_040, w_000_041, w_000_042, w_000_043, w_000_044, w_000_045, w_000_046, w_000_047, w_000_048, w_000_049, w_000_050, w_000_051, w_000_052, w_000_053, w_000_054, w_000_055, w_000_056, w_000_057, w_000_058, w_000_059, w_000_060, w_000_061, w_000_062, w_000_063, w_000_064, w_000_065, w_000_066, w_000_067, w_000_068, w_000_069, w_000_070, w_000_071, w_000_072, w_000_073, w_000_074, w_000_075, w_000_076, w_000_077, w_000_078, w_000_079, w_000_080, w_000_081, w_000_082, w_000_083, w_000_084, w_000_085, w_000_086, w_000_087, w_000_088, w_000_089, w_000_090, w_000_091, w_000_092, w_000_093, w_000_094, w_000_095, w_000_096, w_000_097, w_000_098, w_000_099, w_000_100, w_000_101, w_000_102, w_000_103, w_000_104, w_000_105, w_000_106, w_000_107, w_000_108, w_000_109, w_000_110, w_000_111, w_000_112, w_000_113, w_000_114, w_000_115, w_000_116, w_000_117, w_000_118, w_000_119, w_000_120, w_000_121, w_000_122, w_000_123, w_000_124, w_000_125, w_000_126, w_000_127, w_000_128, w_000_129, w_000_130, w_000_131, w_000_132, w_000_133, w_000_134, w_000_135, w_000_136, w_000_137, w_000_138, w_000_139, w_000_140, w_000_141, w_000_142, w_000_143, w_000_144, w_000_145, w_000_146, w_000_147, w_000_148, w_000_149, w_000_150, w_000_151, w_000_152, w_000_153, w_000_154, w_000_155, w_000_156, w_000_157, w_000_158, w_000_159, w_000_160, w_000_161, w_000_162, w_000_163, w_000_164, w_000_165, w_000_166, w_000_167, w_000_169, w_000_170, w_000_171, w_000_172, w_000_173, w_000_174, w_000_175, w_000_176, w_000_177, w_000_178, w_000_179, w_000_180, w_000_181, w_000_182, w_000_183, w_000_184, w_000_185, w_000_186, w_000_187, w_000_188, w_000_189, w_000_190, w_000_191, w_000_192, w_000_193, w_000_194, w_000_195, w_000_196, w_000_197, w_000_198, w_000_199, w_000_200, w_000_202, w_000_203, w_000_204, w_000_205, w_000_206, w_000_207, w_000_208, w_000_209, w_000_210, w_000_211, w_000_212, w_000_213, w_000_214, w_000_215, w_000_216, w_000_217, w_000_218, w_000_219, w_000_220, w_000_221, w_000_222, w_000_223, w_000_224, w_000_225, w_000_226, w_000_227, w_000_228, w_000_229, w_000_230, w_000_231, w_000_232, w_000_233, w_000_234, w_000_235, w_000_236, w_000_237, w_000_238, w_000_239, w_000_240, w_000_241, w_000_242, w_000_243, w_000_244, w_000_245, w_000_246, w_000_247, w_000_248, w_000_249, w_000_250, w_000_251, w_000_252, w_000_253, w_000_254, w_000_255, w_000_256, w_000_257, w_000_258, w_000_259, w_000_260, w_000_261, w_000_262, w_000_263, w_000_264, w_000_265, w_000_266, w_000_267, w_000_268, w_000_269, w_000_270, w_000_271, w_000_272, w_000_273, w_000_274, w_000_275, w_000_276, w_000_277, w_000_278, w_000_279, w_000_280, w_000_281, w_000_282, w_000_283, w_000_284, w_000_285, w_000_286, w_000_287, w_000_288, w_000_289, w_000_290, w_000_291, w_000_292, w_000_293, w_000_294, w_000_295, w_000_296, w_000_297, w_000_298, w_000_299, w_000_300, w_000_301, w_000_302, w_000_303, w_000_304, w_000_305, w_000_306, w_000_307, w_000_308, w_000_309, w_000_310, w_000_311, w_000_312, w_000_313, w_000_314, w_000_315, w_000_316, w_000_317, w_000_318, w_000_319, w_000_320, w_000_321, w_000_322, w_000_323, w_000_324, w_000_325, w_000_326, w_000_327, w_000_328, w_000_329, w_000_330, w_000_331, w_000_332, w_000_333, w_000_334, w_000_335, w_000_336, w_000_337, w_000_338, w_000_339, w_000_340, w_000_341, w_000_342, w_000_343, w_000_344, w_000_345, w_000_346, w_000_347, w_000_348, w_000_349, w_000_350, w_000_351, w_000_352, w_000_353, w_000_354, w_000_355, w_000_356, w_000_357, w_000_358, w_000_359, w_000_360, w_000_361, w_000_362, w_000_363, w_000_364, w_000_365, w_000_366, w_000_367, w_000_368, w_000_370, w_000_371, w_000_372, w_000_373, w_000_374, w_000_375, w_000_376, w_000_377, w_000_378, w_000_379, w_000_380, w_000_381, w_000_382, w_000_383, w_000_384, w_000_385, w_000_386, w_000_387, w_000_388, w_000_389, w_000_390, w_000_391, w_000_392, w_000_393, w_000_394, w_000_395, w_000_396, w_000_397, w_000_398, w_000_399, w_000_400, w_000_401, w_000_402, w_000_403, w_000_404, w_000_405, w_000_406, w_000_408, w_000_409, w_000_410, w_000_411, w_000_412, w_000_413, w_000_414, w_000_415, w_000_416, w_000_417, w_000_418, w_000_419, w_000_420, w_000_421, w_000_422, w_000_423, w_000_424, w_000_425, w_000_426, w_000_427, w_000_428, w_000_429, w_000_430, w_000_431, w_000_432, w_000_433, w_000_434, w_000_435, w_000_436, w_000_437, w_000_438, w_000_439, w_000_440, w_000_441, w_000_442, w_000_443, w_000_444, w_000_445, w_000_446, w_000_447, w_000_448, w_000_449, w_000_450, w_000_451, w_000_452, w_000_453, w_000_454, w_000_455, w_000_456, w_000_457, w_000_458, w_000_459, w_000_460, w_000_461, w_000_462, w_000_463, w_000_464, w_000_465, w_000_466, w_000_467, w_000_468, w_000_469, w_000_470, w_000_471, w_000_472, w_000_473, w_000_474, w_000_475, w_000_476, w_000_477, w_000_478, w_000_479, w_000_480, w_000_481, w_000_482, w_000_483, w_000_484, w_000_485, w_000_486, w_000_487, w_000_488, w_000_489, w_000_490, w_000_491, w_000_492, w_000_493, w_000_494, w_000_495, w_000_496, w_000_497, w_000_498, w_000_499, w_000_500, w_000_501, w_000_502, w_000_503, w_000_504, w_000_505, w_000_506, w_000_507, w_000_508, w_000_510, w_000_511, w_000_512, w_000_513, w_000_514, w_000_515, w_000_516, w_000_517, w_000_518, w_000_519, w_000_520, w_000_521, w_000_522, w_000_523, w_000_524, w_000_525, w_000_526, w_000_527, w_000_528, w_000_529, w_000_530, w_000_531, w_000_532, w_000_533, w_000_534, w_000_535, w_000_536, w_000_537, w_000_538, w_000_540, w_000_541, w_000_542, w_000_543, w_000_544, w_000_545, w_000_546, w_000_547, w_000_548, w_000_549, w_000_550, w_000_551, w_000_552, w_000_553, w_000_554, w_000_555, w_000_556, w_000_557, w_000_558, w_000_559, w_000_560, w_000_561, w_000_563, w_000_564, w_000_565, w_000_566, w_000_567, w_000_568, w_000_569, w_000_570, w_000_571, w_000_572, w_000_573, w_000_574, w_000_575, w_000_576, w_000_577, w_000_578, w_000_579, w_000_580, w_000_581, w_000_582, w_000_583, w_000_584, w_000_585, w_000_586, w_000_587, w_000_588, w_000_589, w_000_590, w_000_591, w_000_592, w_000_593, w_000_594, w_000_595, w_000_596, w_000_597, w_000_598, w_000_599, w_000_600, w_000_601, w_000_602, w_000_603, w_000_604, w_000_605, w_000_606, w_000_607, w_000_608, w_000_609, w_000_610, w_000_611, w_000_612, w_000_613, w_000_614, w_000_615, w_000_616, w_000_617, w_000_618, w_000_619, w_000_620, w_000_621, w_000_622, w_000_623, w_000_624, w_000_625, w_000_626, w_000_627, w_000_628, w_000_629, w_000_630, w_000_632, w_000_634, w_000_635, w_000_636, w_000_637, w_000_638, w_000_639, w_000_640, w_000_641, w_000_642, w_000_643, w_000_644, w_000_645, w_000_646, w_000_647, w_000_648, w_000_649, w_000_650, w_000_651, w_000_652, w_000_653, w_000_654, w_000_655, w_000_656, w_000_657, w_000_658, w_000_659, w_000_660, w_000_661, w_000_662, w_000_663, w_000_664, w_000_665, w_000_666, w_000_667, w_000_668, w_000_671, w_000_674, w_000_675, w_000_676, w_000_679, w_000_680, w_000_681, w_000_682, w_000_683, w_000_684, w_000_685, w_000_687, w_000_688, w_000_689, w_000_690, w_000_691, w_000_692, w_000_693, w_000_694, w_000_695, w_000_696, w_000_697, w_000_698, w_000_699, w_000_701, w_000_702, w_000_703, w_000_704, w_000_705, w_000_706, w_000_707, w_000_708, w_000_709, w_000_710, w_000_711, w_000_712, w_000_713, w_000_714, w_000_715, w_000_716, w_000_717, w_000_718, w_000_720, w_000_722, w_000_724, w_000_725, w_000_726, w_000_727, w_000_728, w_000_731, w_000_732, w_000_733, w_000_734, w_000_735, w_000_736, w_000_738, w_000_739, w_000_740, w_000_741, w_000_743, w_000_744, w_000_745, w_000_747, w_000_748, w_000_749, w_000_751, w_000_754, w_000_756, w_000_757, w_000_758, w_000_759, w_000_762, w_000_763, w_000_768, w_000_770, w_000_772, w_000_776, w_000_777, w_000_780, w_000_783;
  output w_800_000, w_800_001, w_800_002, w_800_003, w_800_004, w_800_005, w_800_006, w_800_007, w_800_008, w_800_009, w_800_010, w_800_011, w_800_012, w_800_013, w_800_014, w_800_015, w_800_016, w_800_017, w_800_018, w_800_019, w_800_020, w_800_021, w_800_022, w_800_023, w_800_024, w_800_025, w_800_026, w_800_027, w_800_028, w_800_029, w_800_030, w_800_031, w_800_032, w_800_033, w_800_034, w_800_035, w_800_036, w_800_037, w_800_038, w_800_039, w_800_040, w_800_041, w_800_042, w_800_043, w_800_044, w_800_045, w_800_046, w_800_047, w_800_048, w_800_049, w_800_050, w_800_051, w_800_052, w_800_053, w_800_054, w_800_055, w_800_056, w_800_057, w_800_058, w_800_059, w_800_060, w_800_061, w_800_062, w_800_063, w_800_064, w_800_065, w_800_066, w_800_067, w_800_068, w_800_069, w_800_070, w_800_071, w_800_072, w_800_073, w_800_074, w_800_075, w_800_076, w_800_077, w_800_078, w_800_079, w_800_080, w_800_081, w_800_082, w_800_083, w_800_084, w_800_085, w_800_086, w_800_087, w_800_088, w_800_089, w_800_090, w_800_091, w_800_092, w_800_093, w_800_094, w_800_095, w_800_096, w_800_097, w_800_098, w_800_099, w_800_100, w_800_101, w_800_102, w_800_103, w_800_104, w_800_105, w_800_106, w_800_107, w_800_108, w_800_109, w_800_110, w_800_111, w_800_112, w_800_113, w_800_114, w_800_115, w_800_116, w_800_117, w_800_118, w_800_119, w_800_120, w_800_121, w_800_122, w_800_123, w_800_124, w_800_125, w_800_126, w_800_127, w_800_128, w_800_129, w_800_130, w_800_131, w_800_132, w_800_133, w_800_134, w_800_135, w_800_136, w_800_137, w_800_138, w_800_139, w_800_140, w_800_141, w_800_142, w_800_143, w_800_144, w_800_145, w_800_146, w_800_147, w_800_148, w_800_149, w_800_150, w_800_151, w_800_152, w_800_153, w_800_154, w_800_155, w_800_156, w_800_157, w_800_158, w_800_159, w_800_160, w_800_161, w_800_162, w_800_163, w_800_164, w_800_165, w_800_166, w_800_167, w_800_168, w_800_169, w_800_170, w_800_171, w_800_172, w_800_173, w_800_174, w_800_175, w_800_176, w_800_177, w_800_178, w_800_179, w_800_180, w_800_181, w_800_182, w_800_183, w_800_184, w_800_185, w_800_186, w_800_187, w_800_188, w_800_189, w_800_190, w_800_191, w_800_192, w_800_193, w_800_194, w_800_195, w_800_196, w_800_197, w_800_198, w_800_199, w_800_200, w_800_201, w_800_202, w_800_203, w_800_204, w_800_205, w_800_206, w_800_207, w_800_208, w_800_209, w_800_210, w_800_211, w_800_212, w_800_213, w_800_214, w_800_215, w_800_216, w_800_217, w_800_218, w_800_219, w_800_220, w_800_221, w_800_222, w_800_223, w_800_224, w_800_225, w_800_226, w_800_227, w_800_228, w_800_229, w_800_230, w_800_231, w_800_232, w_800_233, w_800_234, w_800_235, w_800_236, w_800_237, w_800_238, w_800_239, w_800_240, w_800_241, w_800_242, w_800_243, w_800_244, w_800_245, w_800_246, w_800_247, w_800_248, w_800_249, w_800_250, w_800_251, w_800_252, w_800_253, w_800_254, w_800_255, w_800_256, w_800_257, w_800_258, w_800_259, w_800_260, w_800_261, w_800_262, w_800_263, w_800_264, w_800_265, w_800_266, w_800_267, w_800_268, w_800_269, w_800_270, w_800_271, w_800_272, w_800_273, w_800_274, w_800_275, w_800_276, w_800_277, w_800_278, w_800_279, w_800_280, w_800_281, w_800_282, w_800_283, w_800_284, w_800_285, w_800_286, w_800_287, w_800_288, w_800_289, w_800_290, w_800_291, w_800_292, w_800_293, w_800_294, w_800_295, w_800_296, w_800_297, w_800_298, w_800_299, w_800_300, w_800_301, w_800_302, w_800_303, w_800_304, w_800_305, w_800_306, w_800_307, w_800_308, w_800_309, w_800_310, w_800_311, w_800_312, w_800_313, w_800_314, w_800_315, w_800_316, w_800_317, w_800_318, w_800_319, w_800_320, w_800_321, w_800_322, w_800_323, w_800_324, w_800_325, w_800_326, w_800_327, w_800_328, w_800_329, w_800_330, w_800_331, w_800_332, w_800_333, w_800_334, w_800_335, w_800_336, w_800_337, w_800_338, w_800_339, w_800_340, w_800_341, w_800_342, w_800_343, w_800_344, w_800_345, w_800_346, w_800_347, w_800_348, w_800_349, w_800_350, w_800_351, w_800_352, w_800_353, w_800_354, w_800_355, w_800_356, w_800_357, w_800_358, w_800_359, w_800_360, w_800_361, w_800_362, w_800_363, w_800_364, w_800_365, w_800_366, w_800_367, w_800_368, w_800_369, w_800_370, w_800_371, w_800_372, w_800_373, w_800_374, w_800_375, w_800_376, w_800_377, w_800_378, w_800_379, w_800_380, w_800_381, w_800_382, w_800_383, w_800_384, w_800_385, w_800_386, w_800_387, w_800_388, w_800_389, w_800_390, w_800_391, w_800_392, w_800_393, w_800_394, w_800_395, w_800_396, w_800_397, w_800_398, w_800_399, w_800_400, w_800_401, w_800_402, w_800_403, w_800_404, w_800_405, w_800_406, w_800_407, w_800_408, w_800_409, w_800_410, w_800_411, w_800_412, w_800_413, w_800_414, w_800_415, w_800_416, w_800_417, w_800_418, w_800_419, w_800_420, w_800_421, w_800_422, w_800_423, w_800_424, w_800_425, w_800_426, w_800_427, w_800_428, w_800_429, w_800_430, w_800_431, w_800_432, w_800_433, w_800_434, w_800_435, w_800_436, w_800_437, w_800_438, w_800_439, w_800_440, w_800_441, w_800_442, w_800_443, w_800_444, w_800_445, w_800_446, w_800_447, w_800_448, w_800_449, w_800_450, w_800_451, w_800_452, w_800_453, w_800_454, w_800_455, w_800_456, w_800_457, w_800_458, w_800_459, w_800_460, w_800_461, w_800_462, w_800_463, w_800_464, w_800_465, w_800_466, w_800_467, w_800_468, w_800_469, w_800_470, w_800_471, w_800_472, w_800_473, w_800_474, w_800_475, w_800_476, w_800_477, w_800_478, w_800_479, w_800_480, w_800_481, w_800_482, w_800_483, w_800_484, w_800_485, w_800_486, w_800_487, w_800_488, w_800_489, w_800_490, w_800_491, w_800_492, w_800_493, w_800_494, w_800_495, w_800_496, w_800_497, w_800_498, w_800_499, w_800_500, w_800_501, w_800_502, w_800_503, w_800_504, w_800_505, w_800_506, w_800_507, w_800_508, w_800_509, w_800_510, w_800_511, w_800_512, w_800_513, w_800_514, w_800_515, w_800_516, w_800_517, w_800_518, w_800_519, w_800_520, w_800_521, w_800_522, w_800_523, w_800_524, w_800_525, w_800_526, w_800_527, w_800_528, w_800_529, w_800_530, w_800_531, w_800_532, w_800_533, w_800_534, w_800_535, w_800_536, w_800_537, w_800_538, w_800_539, w_800_540, w_800_541, w_800_542, w_800_543, w_800_544, w_800_545, w_800_546, w_800_547, w_800_548, w_800_549, w_800_550, w_800_551, w_800_552, w_800_553, w_800_554, w_800_555, w_800_556, w_800_557, w_800_558, w_800_559, w_800_560, w_800_561, w_800_562, w_800_563, w_800_564, w_800_565, w_800_566, w_800_567, w_800_568, w_800_569, w_800_570, w_800_571, w_800_572, w_800_573, w_800_574, w_800_575, w_800_576, w_800_577, w_800_578, w_800_579, w_800_580, w_800_581, w_800_582, w_800_583, w_800_584, w_800_585, w_800_586, w_800_587, w_800_588, w_800_589, w_800_590, w_800_591, w_800_592, w_800_593, w_800_594, w_800_595, w_800_596, w_800_597, w_800_598, w_800_599, w_800_600, w_800_601, w_800_602, w_800_603, w_800_604, w_800_605, w_800_606, w_800_607, w_800_608, w_800_609, w_800_610, w_800_611, w_800_612, w_800_613, w_800_614, w_800_615, w_800_616, w_800_617, w_800_618, w_800_619, w_800_620, w_800_621, w_800_622, w_800_623, w_800_624, w_800_625, w_800_626, w_800_627, w_800_628, w_800_629, w_800_630, w_800_631, w_800_632, w_800_633, w_800_634, w_800_635, w_800_636, w_800_637, w_800_638, w_800_639, w_800_640, w_800_641, w_800_642, w_800_643, w_800_644, w_800_645, w_800_646, w_800_647, w_800_648, w_800_649, w_800_650, w_800_651, w_800_652, w_800_653, w_800_654, w_800_655, w_800_656, w_800_657, w_800_658, w_800_659, w_800_660, w_800_661, w_800_662, w_800_663, w_800_664, w_800_665, w_800_666, w_800_667, w_800_668, w_800_669, w_800_670, w_800_671, w_800_672, w_800_673, w_800_674, w_800_675, w_800_676, w_800_677, w_800_678, w_800_679, w_800_680, w_800_681, w_800_682, w_800_683, w_800_684, w_800_685, w_800_686, w_800_687, w_800_688, w_800_689, w_800_690, w_800_691, w_800_692, w_800_693, w_800_694, w_800_695, w_800_696, w_800_697, w_800_698, w_800_699, w_800_700, w_800_701, w_800_702, w_800_703, w_800_704, w_800_705, w_800_706, w_800_707, w_800_708, w_800_709, w_800_710, w_800_711, w_800_712, w_800_713, w_800_714, w_800_715, w_800_716, w_800_717;
  wire w_000_000, w_000_001, w_000_002, w_000_003, w_000_004, w_000_005, w_000_006, w_000_007, w_000_008, w_000_009, w_000_010, w_000_011, w_000_012, w_000_013, w_000_014, w_000_015, w_000_016, w_000_017, w_000_018, w_000_019, w_000_020, w_000_021, w_000_022, w_000_023, w_000_024, w_000_025, w_000_026, w_000_027, w_000_028, w_000_029, w_000_030, w_000_031, w_000_032, w_000_033, w_000_034, w_000_035, w_000_036, w_000_037, w_000_038, w_000_039, w_000_040, w_000_041, w_000_042, w_000_043, w_000_044, w_000_045, w_000_046, w_000_047, w_000_048, w_000_049, w_000_050, w_000_051, w_000_052, w_000_053, w_000_054, w_000_055, w_000_056, w_000_057, w_000_058, w_000_059, w_000_060, w_000_061, w_000_062, w_000_063, w_000_064, w_000_065, w_000_066, w_000_067, w_000_068, w_000_069, w_000_070, w_000_071, w_000_072, w_000_073, w_000_074, w_000_075, w_000_076, w_000_077, w_000_078, w_000_079, w_000_080, w_000_081, w_000_082, w_000_083, w_000_084, w_000_085, w_000_086, w_000_087, w_000_088, w_000_089, w_000_090, w_000_091, w_000_092, w_000_093, w_000_094, w_000_095, w_000_096, w_000_097, w_000_098, w_000_099, w_000_100, w_000_101, w_000_102, w_000_103, w_000_104, w_000_105, w_000_106, w_000_107, w_000_108, w_000_109, w_000_110, w_000_111, w_000_112, w_000_113, w_000_114, w_000_115, w_000_116, w_000_117, w_000_118, w_000_119, w_000_120, w_000_121, w_000_122, w_000_123, w_000_124, w_000_125, w_000_126, w_000_127, w_000_128, w_000_129, w_000_130, w_000_131, w_000_132, w_000_133, w_000_134, w_000_135, w_000_136, w_000_137, w_000_138, w_000_139, w_000_140, w_000_141, w_000_142, w_000_143, w_000_144, w_000_145, w_000_146, w_000_147, w_000_148, w_000_149, w_000_150, w_000_151, w_000_152, w_000_153, w_000_154, w_000_155, w_000_156, w_000_157, w_000_158, w_000_159, w_000_160, w_000_161, w_000_162, w_000_163, w_000_164, w_000_165, w_000_166, w_000_167, w_000_169, w_000_170, w_000_171, w_000_172, w_000_173, w_000_174, w_000_175, w_000_176, w_000_177, w_000_178, w_000_179, w_000_180, w_000_181, w_000_182, w_000_183, w_000_184, w_000_185, w_000_186, w_000_187, w_000_188, w_000_189, w_000_190, w_000_191, w_000_192, w_000_193, w_000_194, w_000_195, w_000_196, w_000_197, w_000_198, w_000_199, w_000_200, w_000_202, w_000_203, w_000_204, w_000_205, w_000_206, w_000_207, w_000_208, w_000_209, w_000_210, w_000_211, w_000_212, w_000_213, w_000_214, w_000_215, w_000_216, w_000_217, w_000_218, w_000_219, w_000_220, w_000_221, w_000_222, w_000_223, w_000_224, w_000_225, w_000_226, w_000_227, w_000_228, w_000_229, w_000_230, w_000_231, w_000_232, w_000_233, w_000_234, w_000_235, w_000_236, w_000_237, w_000_238, w_000_239, w_000_240, w_000_241, w_000_242, w_000_243, w_000_244, w_000_245, w_000_246, w_000_247, w_000_248, w_000_249, w_000_250, w_000_251, w_000_252, w_000_253, w_000_254, w_000_255, w_000_256, w_000_257, w_000_258, w_000_259, w_000_260, w_000_261, w_000_262, w_000_263, w_000_264, w_000_265, w_000_266, w_000_267, w_000_268, w_000_269, w_000_270, w_000_271, w_000_272, w_000_273, w_000_274, w_000_275, w_000_276, w_000_277, w_000_278, w_000_279, w_000_280, w_000_281, w_000_282, w_000_283, w_000_284, w_000_285, w_000_286, w_000_287, w_000_288, w_000_289, w_000_290, w_000_291, w_000_292, w_000_293, w_000_294, w_000_295, w_000_296, w_000_297, w_000_298, w_000_299, w_000_300, w_000_301, w_000_302, w_000_303, w_000_304, w_000_305, w_000_306, w_000_307, w_000_308, w_000_309, w_000_310, w_000_311, w_000_312, w_000_313, w_000_314, w_000_315, w_000_316, w_000_317, w_000_318, w_000_319, w_000_320, w_000_321, w_000_322, w_000_323, w_000_324, w_000_325, w_000_326, w_000_327, w_000_328, w_000_329, w_000_330, w_000_331, w_000_332, w_000_333, w_000_334, w_000_335, w_000_336, w_000_337, w_000_338, w_000_339, w_000_340, w_000_341, w_000_342, w_000_343, w_000_344, w_000_345, w_000_346, w_000_347, w_000_348, w_000_349, w_000_350, w_000_351, w_000_352, w_000_353, w_000_354, w_000_355, w_000_356, w_000_357, w_000_358, w_000_359, w_000_360, w_000_361, w_000_362, w_000_363, w_000_364, w_000_365, w_000_366, w_000_367, w_000_368, w_000_370, w_000_371, w_000_372, w_000_373, w_000_374, w_000_375, w_000_376, w_000_377, w_000_378, w_000_379, w_000_380, w_000_381, w_000_382, w_000_383, w_000_384, w_000_385, w_000_386, w_000_387, w_000_388, w_000_389, w_000_390, w_000_391, w_000_392, w_000_393, w_000_394, w_000_395, w_000_396, w_000_397, w_000_398, w_000_399, w_000_400, w_000_401, w_000_402, w_000_403, w_000_404, w_000_405, w_000_406, w_000_408, w_000_409, w_000_410, w_000_411, w_000_412, w_000_413, w_000_414, w_000_415, w_000_416, w_000_417, w_000_418, w_000_419, w_000_420, w_000_421, w_000_422, w_000_423, w_000_424, w_000_425, w_000_426, w_000_427, w_000_428, w_000_429, w_000_430, w_000_431, w_000_432, w_000_433, w_000_434, w_000_435, w_000_436, w_000_437, w_000_438, w_000_439, w_000_440, w_000_441, w_000_442, w_000_443, w_000_444, w_000_445, w_000_446, w_000_447, w_000_448, w_000_449, w_000_450, w_000_451, w_000_452, w_000_453, w_000_454, w_000_455, w_000_456, w_000_457, w_000_458, w_000_459, w_000_460, w_000_461, w_000_462, w_000_463, w_000_464, w_000_465, w_000_466, w_000_467, w_000_468, w_000_469, w_000_470, w_000_471, w_000_472, w_000_473, w_000_474, w_000_475, w_000_476, w_000_477, w_000_478, w_000_479, w_000_480, w_000_481, w_000_482, w_000_483, w_000_484, w_000_485, w_000_486, w_000_487, w_000_488, w_000_489, w_000_490, w_000_491, w_000_492, w_000_493, w_000_494, w_000_495, w_000_496, w_000_497, w_000_498, w_000_499, w_000_500, w_000_501, w_000_502, w_000_503, w_000_504, w_000_505, w_000_506, w_000_507, w_000_508, w_000_510, w_000_511, w_000_512, w_000_513, w_000_514, w_000_515, w_000_516, w_000_517, w_000_518, w_000_519, w_000_520, w_000_521, w_000_522, w_000_523, w_000_524, w_000_525, w_000_526, w_000_527, w_000_528, w_000_529, w_000_530, w_000_531, w_000_532, w_000_533, w_000_534, w_000_535, w_000_536, w_000_537, w_000_538, w_000_540, w_000_541, w_000_542, w_000_543, w_000_544, w_000_545, w_000_546, w_000_547, w_000_548, w_000_549, w_000_550, w_000_551, w_000_552, w_000_553, w_000_554, w_000_555, w_000_556, w_000_557, w_000_558, w_000_559, w_000_560, w_000_561, w_000_563, w_000_564, w_000_565, w_000_566, w_000_567, w_000_568, w_000_569, w_000_570, w_000_571, w_000_572, w_000_573, w_000_574, w_000_575, w_000_576, w_000_577, w_000_578, w_000_579, w_000_580, w_000_581, w_000_582, w_000_583, w_000_584, w_000_585, w_000_586, w_000_587, w_000_588, w_000_589, w_000_590, w_000_591, w_000_592, w_000_593, w_000_594, w_000_595, w_000_596, w_000_597, w_000_598, w_000_599, w_000_600, w_000_601, w_000_602, w_000_603, w_000_604, w_000_605, w_000_606, w_000_607, w_000_608, w_000_609, w_000_610, w_000_611, w_000_612, w_000_613, w_000_614, w_000_615, w_000_616, w_000_617, w_000_618, w_000_619, w_000_620, w_000_621, w_000_622, w_000_623, w_000_624, w_000_625, w_000_626, w_000_627, w_000_628, w_000_629, w_000_630, w_000_632, w_000_634, w_000_635, w_000_636, w_000_637, w_000_638, w_000_639, w_000_640, w_000_641, w_000_642, w_000_643, w_000_644, w_000_645, w_000_646, w_000_647, w_000_648, w_000_649, w_000_650, w_000_651, w_000_652, w_000_653, w_000_654, w_000_655, w_000_656, w_000_657, w_000_658, w_000_659, w_000_660, w_000_661, w_000_662, w_000_663, w_000_664, w_000_665, w_000_666, w_000_667, w_000_668, w_000_671, w_000_674, w_000_675, w_000_676, w_000_679, w_000_680, w_000_681, w_000_682, w_000_683, w_000_684, w_000_685, w_000_687, w_000_688, w_000_689, w_000_690, w_000_691, w_000_692, w_000_693, w_000_694, w_000_695, w_000_696, w_000_697, w_000_698, w_000_699, w_000_701, w_000_702, w_000_703, w_000_704, w_000_705, w_000_706, w_000_707, w_000_708, w_000_709, w_000_710, w_000_711, w_000_712, w_000_713, w_000_714, w_000_715, w_000_716, w_000_717, w_000_718, w_000_720, w_000_722, w_000_724, w_000_725, w_000_726, w_000_727, w_000_728, w_000_731, w_000_732, w_000_733, w_000_734, w_000_735, w_000_736, w_000_738, w_000_739, w_000_740, w_000_741, w_000_743, w_000_744, w_000_745, w_000_747, w_000_748, w_000_749, w_000_751, w_000_754, w_000_756, w_000_757, w_000_758, w_000_759, w_000_762, w_000_763, w_000_768, w_000_770, w_000_772, w_000_776, w_000_777, w_000_780, w_000_783;
  wire w_001_000, w_001_001, w_001_002, w_001_003, w_001_004, w_001_005, w_001_006, w_001_007, w_001_008, w_001_009, w_001_010, w_001_011, w_001_012, w_001_013, w_001_014, w_001_015, w_001_016, w_001_017, w_001_018, w_001_019, w_001_020, w_001_021, w_001_022, w_001_023, w_001_024, w_001_025, w_001_026, w_001_027, w_001_028, w_001_029, w_001_030, w_001_031, w_001_032, w_001_033, w_001_034, w_001_035, w_001_036;
  wire w_002_000, w_002_001, w_002_002, w_002_003, w_002_004, w_002_005, w_002_006, w_002_007, w_002_008, w_002_009, w_002_010, w_002_011, w_002_012, w_002_013, w_002_014, w_002_015, w_002_016, w_002_017, w_002_018, w_002_019, w_002_020, w_002_021, w_002_022, w_002_023, w_002_024, w_002_025, w_002_026, w_002_027, w_002_028, w_002_029, w_002_030, w_002_031, w_002_032, w_002_033, w_002_034, w_002_035, w_002_036, w_002_037, w_002_038, w_002_039, w_002_040, w_002_041, w_002_042, w_002_043, w_002_044, w_002_045, w_002_046, w_002_047, w_002_048, w_002_049, w_002_050, w_002_051, w_002_052, w_002_053, w_002_054, w_002_055, w_002_056, w_002_057, w_002_058, w_002_059, w_002_060, w_002_061, w_002_062, w_002_063, w_002_064, w_002_065, w_002_066, w_002_067, w_002_068, w_002_069, w_002_070, w_002_071, w_002_072, w_002_073, w_002_074, w_002_075, w_002_076, w_002_077, w_002_078, w_002_079, w_002_080, w_002_081, w_002_082, w_002_083, w_002_084, w_002_085, w_002_086, w_002_087, w_002_088, w_002_090, w_002_091, w_002_092, w_002_093, w_002_094, w_002_096, w_002_097, w_002_098, w_002_099, w_002_100, w_002_101, w_002_102, w_002_103, w_002_104, w_002_105, w_002_106, w_002_107, w_002_108, w_002_109, w_002_110, w_002_112, w_002_113, w_002_114, w_002_115, w_002_116, w_002_118, w_002_119, w_002_120, w_002_121, w_002_123, w_002_124, w_002_125, w_002_127, w_002_128, w_002_129, w_002_130, w_002_133, w_002_134, w_002_135, w_002_137, w_002_139, w_002_141, w_002_142, w_002_144, w_002_145, w_002_146, w_002_147, w_002_148, w_002_149, w_002_150, w_002_151, w_002_152, w_002_154, w_002_155, w_002_157, w_002_158, w_002_159, w_002_161, w_002_162, w_002_163, w_002_165, w_002_166, w_002_167, w_002_168, w_002_170, w_002_171, w_002_172, w_002_173, w_002_174, w_002_175, w_002_176, w_002_178, w_002_179, w_002_180, w_002_181, w_002_182, w_002_183, w_002_184, w_002_186, w_002_188, w_002_189, w_002_190, w_002_191, w_002_192, w_002_193, w_002_194, w_002_195, w_002_196, w_002_198, w_002_200, w_002_201, w_002_202, w_002_204, w_002_205, w_002_206, w_002_207, w_002_209, w_002_210, w_002_211, w_002_212, w_002_213, w_002_214, w_002_215, w_002_216, w_002_217, w_002_218, w_002_219, w_002_220, w_002_221, w_002_222, w_002_223, w_002_224, w_002_225, w_002_226, w_002_227, w_002_228, w_002_229, w_002_230, w_002_231, w_002_233, w_002_234, w_002_236, w_002_237, w_002_238, w_002_239, w_002_240, w_002_243, w_002_244, w_002_246, w_002_247, w_002_249, w_002_250, w_002_251, w_002_252, w_002_253, w_002_256, w_002_257, w_002_258, w_002_259, w_002_260, w_002_261, w_002_262, w_002_263, w_002_264, w_002_265, w_002_266, w_002_267, w_002_268, w_002_269, w_002_270, w_002_271, w_002_272, w_002_273, w_002_274, w_002_275, w_002_276, w_002_277, w_002_278, w_002_279, w_002_280, w_002_282, w_002_283, w_002_285, w_002_286, w_002_287, w_002_288, w_002_289, w_002_290, w_002_291, w_002_292, w_002_293, w_002_295, w_002_296, w_002_297, w_002_298, w_002_299, w_002_300, w_002_301, w_002_302, w_002_303, w_002_304, w_002_305, w_002_306, w_002_307, w_002_308, w_002_309, w_002_310, w_002_311, w_002_312, w_002_313, w_002_315, w_002_316, w_002_317, w_002_318, w_002_319, w_002_320, w_002_321, w_002_322, w_002_323, w_002_324, w_002_326, w_002_327, w_002_328, w_002_329, w_002_330, w_002_331, w_002_334, w_002_335, w_002_337, w_002_338, w_002_340, w_002_341, w_002_342, w_002_343, w_002_344, w_002_345, w_002_346, w_002_347, w_002_349, w_002_350, w_002_351, w_002_352, w_002_353, w_002_354, w_002_357, w_002_358, w_002_359, w_002_360, w_002_361, w_002_362, w_002_363, w_002_365, w_002_366, w_002_367, w_002_368, w_002_369, w_002_370, w_002_372, w_002_373, w_002_374, w_002_375, w_002_376, w_002_377, w_002_378, w_002_379, w_002_380, w_002_383, w_002_384, w_002_385, w_002_386, w_002_389, w_002_390, w_002_391, w_002_392, w_002_393, w_002_396, w_002_397, w_002_398, w_002_400, w_002_401, w_002_402, w_002_403, w_002_405, w_002_406, w_002_407, w_002_408, w_002_409, w_002_411, w_002_412, w_002_413, w_002_414, w_002_415, w_002_416, w_002_417, w_002_418, w_002_419, w_002_420, w_002_421, w_002_423, w_002_424, w_002_425, w_002_426, w_002_427, w_002_428, w_002_429, w_002_433, w_002_434, w_002_435, w_002_436, w_002_438, w_002_439, w_002_440, w_002_441, w_002_442, w_002_443, w_002_444, w_002_445, w_002_446, w_002_447, w_002_448, w_002_449, w_002_450, w_002_451, w_002_452, w_002_453, w_002_455, w_002_457, w_002_458, w_002_459, w_002_460, w_002_461, w_002_462, w_002_464, w_002_465, w_002_466, w_002_467, w_002_468, w_002_469, w_002_470, w_002_471, w_002_472, w_002_473, w_002_474, w_002_475, w_002_477, w_002_478, w_002_479, w_002_480, w_002_481, w_002_482, w_002_485, w_002_486, w_002_487, w_002_488, w_002_489, w_002_490, w_002_491, w_002_493, w_002_494, w_002_495, w_002_496, w_002_497, w_002_498, w_002_499, w_002_500, w_002_501, w_002_502, w_002_503, w_002_504, w_002_505, w_002_507, w_002_509, w_002_510, w_002_511, w_002_512, w_002_513, w_002_514, w_002_515, w_002_516, w_002_517, w_002_518, w_002_519, w_002_520, w_002_522, w_002_523, w_002_524, w_002_526, w_002_528, w_002_529, w_002_530, w_002_531, w_002_532, w_002_533, w_002_534, w_002_535, w_002_536, w_002_537, w_002_538, w_002_540, w_002_541, w_002_542, w_002_543, w_002_545, w_002_547, w_002_548, w_002_549, w_002_550, w_002_551, w_002_552, w_002_553, w_002_554, w_002_557, w_002_558, w_002_560, w_002_561, w_002_562, w_002_563, w_002_564, w_002_565, w_002_566, w_002_567, w_002_568, w_002_569, w_002_570, w_002_571, w_002_572, w_002_574, w_002_575, w_002_576, w_002_577, w_002_578, w_002_579, w_002_580, w_002_581, w_002_582, w_002_583, w_002_584, w_002_585, w_002_586, w_002_587, w_002_588, w_002_589, w_002_590, w_002_591, w_002_592, w_002_593, w_002_594, w_002_595, w_002_596, w_002_597, w_002_598, w_002_599, w_002_600, w_002_601, w_002_602, w_002_603, w_002_604, w_002_605, w_002_606, w_002_607, w_002_608, w_002_609, w_002_610, w_002_612, w_002_613, w_002_614, w_002_615, w_002_616, w_002_617, w_002_618, w_002_619, w_002_620, w_002_621, w_002_622, w_002_623, w_002_624, w_002_625, w_002_626, w_002_627, w_002_628, w_002_629, w_002_631, w_002_632, w_002_633, w_002_634, w_002_635, w_002_636, w_002_638, w_002_639, w_002_640, w_002_642, w_002_643, w_002_644, w_002_645, w_002_646, w_002_647, w_002_648, w_002_650, w_002_651, w_002_652, w_002_653, w_002_654, w_002_655, w_002_656, w_002_657, w_002_658, w_002_659, w_002_660, w_002_661, w_002_662, w_002_664, w_002_665, w_002_666, w_002_667, w_002_668, w_002_669, w_002_671, w_002_672, w_002_673, w_002_674, w_002_676, w_002_677, w_002_678, w_002_679, w_002_681, w_002_682, w_002_683, w_002_684, w_002_685, w_002_686, w_002_688, w_002_690, w_002_691, w_002_692, w_002_693, w_002_694, w_002_695, w_002_696, w_002_697, w_002_698, w_002_699, w_002_701, w_002_702, w_002_703, w_002_705, w_002_706, w_002_707, w_002_708, w_002_709, w_002_710, w_002_711;
  wire w_003_000, w_003_001, w_003_002, w_003_003, w_003_004, w_003_005, w_003_006, w_003_007, w_003_008, w_003_009, w_003_010, w_003_011, w_003_012, w_003_013, w_003_014, w_003_015, w_003_016, w_003_017, w_003_018, w_003_019, w_003_020, w_003_021, w_003_022, w_003_023, w_003_024, w_003_025, w_003_026, w_003_027, w_003_028, w_003_029, w_003_030, w_003_031, w_003_032, w_003_033, w_003_034, w_003_035, w_003_036, w_003_037, w_003_038, w_003_039, w_003_040, w_003_041, w_003_042, w_003_043, w_003_044, w_003_045, w_003_046, w_003_047, w_003_048, w_003_049, w_003_050, w_003_051, w_003_052, w_003_053, w_003_054, w_003_055, w_003_056, w_003_057, w_003_058, w_003_059, w_003_060, w_003_061, w_003_062, w_003_063, w_003_064, w_003_065, w_003_066, w_003_067, w_003_068, w_003_069, w_003_070, w_003_071, w_003_072, w_003_073, w_003_074, w_003_075, w_003_076, w_003_077, w_003_078, w_003_079, w_003_080, w_003_081, w_003_082, w_003_083, w_003_084;
  wire w_004_000, w_004_001, w_004_002, w_004_003, w_004_004, w_004_005, w_004_006, w_004_007, w_004_008, w_004_009, w_004_010, w_004_011, w_004_012, w_004_013, w_004_014, w_004_015, w_004_016, w_004_017, w_004_019, w_004_020, w_004_021, w_004_022, w_004_023, w_004_024, w_004_025, w_004_026, w_004_027, w_004_028, w_004_029, w_004_030, w_004_031, w_004_032, w_004_033, w_004_034, w_004_035, w_004_036, w_004_037, w_004_038, w_004_039, w_004_040, w_004_041, w_004_042, w_004_043, w_004_044, w_004_045, w_004_046, w_004_047, w_004_048, w_004_049, w_004_050, w_004_051, w_004_052, w_004_053, w_004_054, w_004_055, w_004_056, w_004_057, w_004_058, w_004_059, w_004_060, w_004_061, w_004_062, w_004_063, w_004_064, w_004_065, w_004_066, w_004_067, w_004_068, w_004_069, w_004_070, w_004_071, w_004_072, w_004_074, w_004_075, w_004_076, w_004_077, w_004_078, w_004_079, w_004_081, w_004_082, w_004_083, w_004_084, w_004_085, w_004_086, w_004_087, w_004_088, w_004_089, w_004_090, w_004_091, w_004_092, w_004_093, w_004_094, w_004_095, w_004_096, w_004_097, w_004_098, w_004_099, w_004_100, w_004_101, w_004_102, w_004_103, w_004_104, w_004_105, w_004_106, w_004_107, w_004_108, w_004_109, w_004_110, w_004_111, w_004_113, w_004_114, w_004_115, w_004_116, w_004_117, w_004_118, w_004_119, w_004_120, w_004_121, w_004_122, w_004_123, w_004_124, w_004_125, w_004_126, w_004_128, w_004_129, w_004_130, w_004_131, w_004_132, w_004_133, w_004_134, w_004_135, w_004_136, w_004_137, w_004_138, w_004_139, w_004_140, w_004_141, w_004_142, w_004_143, w_004_144, w_004_145, w_004_146, w_004_147, w_004_148, w_004_149, w_004_150, w_004_151, w_004_152, w_004_153, w_004_154, w_004_155, w_004_156, w_004_157, w_004_158, w_004_159, w_004_160, w_004_161, w_004_162, w_004_163, w_004_164, w_004_165, w_004_166, w_004_167, w_004_168, w_004_169, w_004_170, w_004_171, w_004_172, w_004_173, w_004_174, w_004_175, w_004_176, w_004_177, w_004_178, w_004_179, w_004_180, w_004_181, w_004_182, w_004_183, w_004_184, w_004_185, w_004_186, w_004_187, w_004_188, w_004_190, w_004_191, w_004_192, w_004_193, w_004_194, w_004_195, w_004_196, w_004_197, w_004_198, w_004_199, w_004_200, w_004_201, w_004_202, w_004_203, w_004_204, w_004_205, w_004_206, w_004_207, w_004_208, w_004_209, w_004_210, w_004_211, w_004_212, w_004_213, w_004_214, w_004_215, w_004_216, w_004_217, w_004_218, w_004_219, w_004_220, w_004_221, w_004_222, w_004_223, w_004_224, w_004_225, w_004_226, w_004_227, w_004_228, w_004_229, w_004_230, w_004_231, w_004_232, w_004_235, w_004_236, w_004_237, w_004_238, w_004_239, w_004_240, w_004_241, w_004_242, w_004_243, w_004_244, w_004_245, w_004_246, w_004_247, w_004_248, w_004_249, w_004_250, w_004_252, w_004_253, w_004_254, w_004_255, w_004_256, w_004_257, w_004_259, w_004_260, w_004_261, w_004_262, w_004_263, w_004_264, w_004_265, w_004_266, w_004_267, w_004_268, w_004_269, w_004_270, w_004_271, w_004_272, w_004_273, w_004_274, w_004_275, w_004_276, w_004_277, w_004_278, w_004_279, w_004_280, w_004_281, w_004_282, w_004_283, w_004_284, w_004_285, w_004_286, w_004_287, w_004_288, w_004_289, w_004_290, w_004_291, w_004_292, w_004_293, w_004_294, w_004_295, w_004_296, w_004_297, w_004_299, w_004_301, w_004_302, w_004_304, w_004_305, w_004_307, w_004_308, w_004_309, w_004_310, w_004_311, w_004_314, w_004_315, w_004_316, w_004_317, w_004_319, w_004_320, w_004_321, w_004_322, w_004_325, w_004_326, w_004_328, w_004_329, w_004_330, w_004_331, w_004_332, w_004_333, w_004_335, w_004_336, w_004_337, w_004_338, w_004_340, w_004_341, w_004_343, w_004_344, w_004_345, w_004_346, w_004_347, w_004_348, w_004_349, w_004_350, w_004_351, w_004_352, w_004_353, w_004_354, w_004_355, w_004_357, w_004_359, w_004_360, w_004_361, w_004_362, w_004_363, w_004_364, w_004_365, w_004_366, w_004_367, w_004_368, w_004_369, w_004_370, w_004_371, w_004_372, w_004_373, w_004_374, w_004_375, w_004_376, w_004_377, w_004_378, w_004_379, w_004_380, w_004_382, w_004_383, w_004_384, w_004_386, w_004_387, w_004_388, w_004_389, w_004_390, w_004_391, w_004_392, w_004_393, w_004_394, w_004_395, w_004_396, w_004_397, w_004_398, w_004_399, w_004_400, w_004_401, w_004_402, w_004_405, w_004_406, w_004_407, w_004_408, w_004_409, w_004_410, w_004_411, w_004_413, w_004_414, w_004_415, w_004_416, w_004_418, w_004_419, w_004_420, w_004_421, w_004_423, w_004_424, w_004_425, w_004_426, w_004_427, w_004_428, w_004_429, w_004_431, w_004_432, w_004_433, w_004_434, w_004_435, w_004_436, w_004_437, w_004_438, w_004_439, w_004_440, w_004_441, w_004_443, w_004_444, w_004_445, w_004_446, w_004_447, w_004_448, w_004_449, w_004_450, w_004_451, w_004_452, w_004_453, w_004_454, w_004_455, w_004_456, w_004_457, w_004_459, w_004_460, w_004_462, w_004_463, w_004_464, w_004_465, w_004_466, w_004_468, w_004_469, w_004_470, w_004_471, w_004_472, w_004_473, w_004_474, w_004_476, w_004_477, w_004_478, w_004_479, w_004_480, w_004_482, w_004_484, w_004_486, w_004_487, w_004_488, w_004_489, w_004_490, w_004_491, w_004_492, w_004_493, w_004_495, w_004_496, w_004_497, w_004_498, w_004_499, w_004_500, w_004_501, w_004_502, w_004_503, w_004_505, w_004_506, w_004_507, w_004_508;
  wire w_005_000, w_005_001, w_005_002, w_005_003, w_005_004, w_005_005, w_005_006, w_005_007, w_005_008, w_005_009, w_005_010, w_005_011, w_005_012, w_005_013, w_005_014, w_005_015, w_005_016, w_005_017, w_005_018, w_005_019, w_005_020, w_005_021, w_005_022, w_005_023, w_005_024, w_005_025, w_005_026, w_005_027, w_005_028, w_005_029, w_005_030, w_005_031, w_005_032, w_005_033, w_005_034, w_005_035, w_005_036, w_005_037, w_005_038, w_005_039, w_005_040, w_005_041, w_005_042, w_005_043, w_005_044, w_005_046, w_005_047, w_005_048, w_005_049, w_005_050, w_005_051, w_005_052, w_005_053, w_005_054, w_005_055, w_005_056, w_005_057, w_005_058, w_005_059, w_005_060, w_005_061, w_005_062, w_005_063, w_005_064, w_005_065, w_005_066, w_005_067, w_005_068, w_005_069, w_005_070, w_005_071, w_005_072, w_005_073, w_005_074, w_005_075, w_005_076, w_005_077, w_005_078, w_005_079, w_005_080, w_005_081, w_005_083, w_005_084, w_005_085, w_005_086, w_005_087, w_005_088, w_005_089, w_005_090, w_005_091, w_005_092, w_005_093, w_005_094, w_005_095, w_005_096, w_005_097, w_005_098, w_005_099, w_005_100, w_005_101, w_005_102, w_005_103, w_005_104, w_005_105, w_005_106, w_005_107, w_005_108, w_005_109, w_005_110, w_005_111, w_005_112, w_005_113, w_005_114, w_005_115, w_005_116, w_005_117, w_005_118, w_005_119, w_005_120, w_005_121, w_005_122, w_005_123, w_005_124, w_005_125, w_005_126, w_005_127, w_005_128, w_005_129, w_005_130, w_005_131, w_005_132, w_005_133, w_005_134, w_005_135, w_005_136, w_005_137, w_005_138, w_005_139, w_005_140, w_005_141, w_005_142, w_005_143, w_005_144, w_005_145, w_005_146, w_005_147, w_005_148, w_005_149, w_005_150, w_005_151, w_005_152, w_005_153, w_005_154, w_005_155, w_005_156, w_005_157, w_005_158, w_005_159, w_005_160, w_005_161, w_005_162, w_005_163, w_005_164, w_005_165, w_005_166, w_005_167, w_005_168, w_005_169, w_005_170, w_005_171, w_005_172, w_005_173, w_005_174, w_005_175, w_005_176, w_005_177, w_005_178, w_005_180, w_005_181, w_005_182, w_005_183, w_005_184, w_005_185, w_005_186, w_005_187, w_005_188, w_005_189, w_005_190, w_005_191, w_005_192, w_005_193, w_005_194, w_005_195, w_005_196, w_005_197, w_005_198, w_005_199, w_005_200, w_005_201, w_005_202, w_005_204, w_005_205, w_005_206, w_005_207, w_005_208, w_005_209, w_005_210, w_005_211, w_005_212, w_005_213, w_005_214, w_005_215, w_005_216, w_005_218, w_005_219, w_005_220, w_005_221, w_005_223, w_005_224, w_005_225, w_005_226, w_005_227, w_005_228, w_005_229, w_005_230, w_005_231, w_005_232, w_005_233, w_005_234, w_005_235, w_005_236, w_005_237, w_005_238, w_005_239, w_005_240, w_005_242, w_005_243, w_005_244, w_005_245, w_005_246, w_005_247, w_005_248, w_005_249, w_005_250, w_005_251, w_005_252, w_005_254, w_005_255, w_005_256, w_005_257, w_005_259, w_005_260, w_005_261, w_005_262, w_005_263, w_005_266, w_005_267, w_005_268, w_005_270, w_005_271, w_005_272, w_005_273, w_005_274, w_005_275, w_005_276, w_005_277, w_005_278, w_005_279, w_005_280, w_005_281, w_005_282, w_005_283, w_005_285, w_005_286, w_005_287, w_005_288, w_005_289, w_005_290, w_005_291, w_005_292, w_005_293, w_005_294, w_005_295, w_005_296, w_005_297, w_005_298, w_005_299, w_005_300, w_005_301, w_005_302, w_005_303, w_005_304, w_005_305, w_005_306, w_005_307, w_005_308, w_005_309, w_005_310, w_005_311, w_005_312, w_005_313, w_005_314, w_005_315, w_005_316, w_005_317, w_005_318;
  wire w_006_000, w_006_001, w_006_002, w_006_003, w_006_004, w_006_005, w_006_006, w_006_007, w_006_008, w_006_009, w_006_010, w_006_011, w_006_012, w_006_013, w_006_014, w_006_015, w_006_016, w_006_017, w_006_018, w_006_019, w_006_020, w_006_021, w_006_022, w_006_023, w_006_024, w_006_025, w_006_026, w_006_027, w_006_028, w_006_029, w_006_030, w_006_031, w_006_032, w_006_033, w_006_034, w_006_035, w_006_036, w_006_037, w_006_038, w_006_039, w_006_040, w_006_041, w_006_042, w_006_043, w_006_044, w_006_045, w_006_047, w_006_048, w_006_049, w_006_051, w_006_052, w_006_053, w_006_054, w_006_055, w_006_056, w_006_057, w_006_058, w_006_059, w_006_060, w_006_061, w_006_062, w_006_063, w_006_064, w_006_065, w_006_066, w_006_067, w_006_068, w_006_069, w_006_070, w_006_071, w_006_072, w_006_073, w_006_074, w_006_075, w_006_076, w_006_077, w_006_078, w_006_079, w_006_080, w_006_081, w_006_082, w_006_083, w_006_084, w_006_085, w_006_086, w_006_087, w_006_088, w_006_089, w_006_090, w_006_091, w_006_092, w_006_093, w_006_094, w_006_095, w_006_096, w_006_097, w_006_098, w_006_099, w_006_100, w_006_101, w_006_102, w_006_103, w_006_104, w_006_105, w_006_106, w_006_107, w_006_108, w_006_109, w_006_110, w_006_111, w_006_112, w_006_113, w_006_114, w_006_115, w_006_116, w_006_117, w_006_118, w_006_119, w_006_120, w_006_121, w_006_122, w_006_123, w_006_124, w_006_125, w_006_126, w_006_127, w_006_128, w_006_129, w_006_130, w_006_131, w_006_132, w_006_133, w_006_134, w_006_135, w_006_136, w_006_137, w_006_138, w_006_139, w_006_140, w_006_141, w_006_142, w_006_143, w_006_144, w_006_145, w_006_146, w_006_147, w_006_148, w_006_149, w_006_150, w_006_151, w_006_152, w_006_153, w_006_154, w_006_155, w_006_156, w_006_157, w_006_158, w_006_159, w_006_160, w_006_161, w_006_162, w_006_163, w_006_164, w_006_165, w_006_166, w_006_167, w_006_168, w_006_169, w_006_170, w_006_171, w_006_172, w_006_173, w_006_174, w_006_175, w_006_176, w_006_177, w_006_178, w_006_179, w_006_180, w_006_181, w_006_182, w_006_183, w_006_184, w_006_185, w_006_186, w_006_187, w_006_188, w_006_189, w_006_190, w_006_191, w_006_192, w_006_193, w_006_194, w_006_195, w_006_196, w_006_197, w_006_198, w_006_199, w_006_200, w_006_201, w_006_202, w_006_203, w_006_204, w_006_205, w_006_206, w_006_207, w_006_208, w_006_209, w_006_210, w_006_211, w_006_212, w_006_213, w_006_214, w_006_215, w_006_216, w_006_217, w_006_218, w_006_219, w_006_220, w_006_221, w_006_222, w_006_223, w_006_224, w_006_225, w_006_226, w_006_227, w_006_228, w_006_229, w_006_230, w_006_231, w_006_232, w_006_233, w_006_234, w_006_235, w_006_236, w_006_237, w_006_238, w_006_239, w_006_240, w_006_241, w_006_242, w_006_243, w_006_244, w_006_245, w_006_246, w_006_247, w_006_248, w_006_249, w_006_250, w_006_251, w_006_252, w_006_254, w_006_255, w_006_256, w_006_258;
  wire w_007_000, w_007_001, w_007_002, w_007_003, w_007_004, w_007_005, w_007_006, w_007_007, w_007_008, w_007_009, w_007_010, w_007_011, w_007_012, w_007_013, w_007_014, w_007_015, w_007_016, w_007_017, w_007_018, w_007_019, w_007_020, w_007_021, w_007_022, w_007_023, w_007_025, w_007_026, w_007_027, w_007_028, w_007_029, w_007_031, w_007_032, w_007_033, w_007_034, w_007_035, w_007_036, w_007_037, w_007_038, w_007_039, w_007_040, w_007_041, w_007_042, w_007_043, w_007_044, w_007_045, w_007_046, w_007_047, w_007_049, w_007_050, w_007_051, w_007_052, w_007_053, w_007_054, w_007_055, w_007_056, w_007_057, w_007_058, w_007_059, w_007_060, w_007_061, w_007_062, w_007_063, w_007_064, w_007_065, w_007_066, w_007_067, w_007_068, w_007_069, w_007_070, w_007_071, w_007_072, w_007_073, w_007_074, w_007_076, w_007_077, w_007_078, w_007_079, w_007_080, w_007_081, w_007_082, w_007_083, w_007_084, w_007_085, w_007_086, w_007_087, w_007_088, w_007_089, w_007_090, w_007_091, w_007_092, w_007_093, w_007_094, w_007_096, w_007_097, w_007_098, w_007_099, w_007_100, w_007_101, w_007_102, w_007_103, w_007_104, w_007_105, w_007_106, w_007_107, w_007_108, w_007_109, w_007_110, w_007_111, w_007_112, w_007_113, w_007_114, w_007_115, w_007_116, w_007_117, w_007_118, w_007_119, w_007_120, w_007_121, w_007_122, w_007_123, w_007_124, w_007_125, w_007_126, w_007_127, w_007_128, w_007_129, w_007_130, w_007_131, w_007_132, w_007_134, w_007_135, w_007_136, w_007_137, w_007_138, w_007_139, w_007_140, w_007_141, w_007_142, w_007_143, w_007_144, w_007_145, w_007_146, w_007_147, w_007_148, w_007_149, w_007_150, w_007_151, w_007_152, w_007_153, w_007_154, w_007_155, w_007_156, w_007_157, w_007_158, w_007_159, w_007_160, w_007_161, w_007_162, w_007_163, w_007_164, w_007_165, w_007_166, w_007_167, w_007_168, w_007_169, w_007_170, w_007_171, w_007_172, w_007_173, w_007_175, w_007_176, w_007_177, w_007_178, w_007_179, w_007_180, w_007_181, w_007_182, w_007_183, w_007_184, w_007_185, w_007_186, w_007_187, w_007_188, w_007_189, w_007_190, w_007_191, w_007_192, w_007_193, w_007_194, w_007_195, w_007_196, w_007_197, w_007_198, w_007_199, w_007_200, w_007_201, w_007_202, w_007_203, w_007_204, w_007_205, w_007_206, w_007_207, w_007_208, w_007_209, w_007_210, w_007_211, w_007_212, w_007_213, w_007_214, w_007_215, w_007_216, w_007_217, w_007_218, w_007_219, w_007_220, w_007_221, w_007_222, w_007_223, w_007_224, w_007_225, w_007_226, w_007_227, w_007_228, w_007_230, w_007_231, w_007_232, w_007_233, w_007_234, w_007_235, w_007_236, w_007_237, w_007_238, w_007_239, w_007_240, w_007_241, w_007_244, w_007_245, w_007_246, w_007_247, w_007_248, w_007_249, w_007_250, w_007_251, w_007_252, w_007_253, w_007_254, w_007_255, w_007_256, w_007_257, w_007_258, w_007_259, w_007_260, w_007_261, w_007_262, w_007_263, w_007_264, w_007_265, w_007_266, w_007_267, w_007_268, w_007_269, w_007_270, w_007_271, w_007_272, w_007_273, w_007_274, w_007_275, w_007_276, w_007_277, w_007_278, w_007_279, w_007_280, w_007_281, w_007_282, w_007_283, w_007_284, w_007_285, w_007_286, w_007_287, w_007_288, w_007_289, w_007_291, w_007_292, w_007_293, w_007_294, w_007_295, w_007_296, w_007_297, w_007_299, w_007_300, w_007_303, w_007_304, w_007_306, w_007_307, w_007_308, w_007_309, w_007_310, w_007_312, w_007_313, w_007_314, w_007_315, w_007_316, w_007_318, w_007_319, w_007_320, w_007_321, w_007_323, w_007_324, w_007_325, w_007_327, w_007_328, w_007_330, w_007_331, w_007_332, w_007_333, w_007_334, w_007_336, w_007_337, w_007_339, w_007_340, w_007_342, w_007_343, w_007_345, w_007_346, w_007_347, w_007_348, w_007_349, w_007_350, w_007_351, w_007_353, w_007_354, w_007_356, w_007_357, w_007_359, w_007_360, w_007_361, w_007_362, w_007_363, w_007_364, w_007_365, w_007_367, w_007_368, w_007_371, w_007_372, w_007_373, w_007_374, w_007_377, w_007_378, w_007_379, w_007_380, w_007_381, w_007_382, w_007_384, w_007_385, w_007_386, w_007_387, w_007_389, w_007_390, w_007_391, w_007_392, w_007_393, w_007_394, w_007_395, w_007_396, w_007_397, w_007_398, w_007_400, w_007_403, w_007_405, w_007_407, w_007_408, w_007_410, w_007_413, w_007_414, w_007_415, w_007_416, w_007_418, w_007_419, w_007_420, w_007_421, w_007_422, w_007_423, w_007_424, w_007_425, w_007_426, w_007_427, w_007_428, w_007_429, w_007_431, w_007_432, w_007_434, w_007_436, w_007_437, w_007_438, w_007_439, w_007_440, w_007_441, w_007_443, w_007_444, w_007_445, w_007_447, w_007_448, w_007_449, w_007_450, w_007_451, w_007_452, w_007_453, w_007_454, w_007_455, w_007_456, w_007_459, w_007_460, w_007_461, w_007_462, w_007_463, w_007_464, w_007_469, w_007_470, w_007_471, w_007_472, w_007_473, w_007_474, w_007_475, w_007_477, w_007_478, w_007_480;
  wire w_008_001, w_008_003, w_008_004, w_008_005, w_008_008, w_008_009, w_008_010, w_008_011, w_008_012, w_008_013, w_008_014, w_008_015, w_008_016, w_008_017, w_008_018, w_008_019, w_008_020, w_008_021, w_008_022, w_008_023, w_008_024, w_008_025, w_008_026, w_008_027, w_008_028, w_008_029, w_008_030, w_008_031, w_008_032, w_008_033, w_008_034, w_008_035, w_008_036, w_008_037, w_008_038, w_008_039, w_008_040, w_008_041, w_008_042, w_008_043, w_008_044, w_008_045, w_008_046, w_008_047, w_008_048, w_008_049, w_008_050, w_008_051, w_008_052, w_008_053, w_008_054, w_008_055, w_008_056, w_008_059, w_008_061, w_008_062, w_008_063, w_008_064, w_008_067, w_008_068, w_008_069, w_008_071, w_008_072, w_008_073, w_008_074, w_008_076, w_008_077, w_008_078, w_008_079, w_008_082, w_008_083, w_008_084, w_008_085, w_008_088, w_008_089, w_008_090, w_008_093, w_008_094, w_008_095, w_008_096, w_008_097, w_008_099, w_008_100, w_008_103, w_008_105, w_008_107, w_008_108, w_008_110, w_008_111, w_008_112, w_008_114, w_008_115, w_008_117, w_008_118, w_008_121, w_008_122, w_008_124, w_008_125, w_008_126, w_008_127, w_008_128, w_008_129, w_008_130, w_008_131, w_008_133, w_008_134, w_008_135, w_008_136, w_008_137, w_008_138, w_008_140, w_008_142, w_008_143, w_008_145, w_008_147, w_008_149, w_008_150, w_008_152, w_008_153, w_008_156, w_008_157, w_008_159, w_008_161, w_008_162, w_008_164, w_008_167, w_008_168, w_008_169, w_008_170, w_008_171, w_008_172, w_008_173, w_008_175, w_008_178, w_008_179, w_008_180, w_008_181, w_008_182, w_008_183, w_008_184, w_008_186, w_008_188, w_008_189, w_008_190, w_008_191, w_008_192, w_008_193, w_008_194, w_008_196, w_008_198, w_008_199, w_008_200, w_008_202, w_008_205, w_008_206, w_008_207, w_008_208, w_008_209, w_008_210, w_008_211, w_008_212, w_008_213, w_008_214, w_008_215, w_008_216, w_008_217, w_008_218, w_008_220, w_008_221, w_008_222, w_008_223, w_008_225, w_008_226, w_008_227, w_008_228, w_008_230, w_008_232, w_008_236, w_008_237, w_008_239, w_008_240, w_008_241, w_008_243, w_008_244, w_008_246, w_008_247, w_008_248, w_008_249, w_008_250, w_008_252, w_008_254, w_008_255, w_008_257, w_008_258, w_008_261, w_008_262, w_008_264, w_008_266, w_008_268, w_008_269, w_008_271, w_008_272, w_008_273, w_008_274, w_008_275, w_008_277, w_008_278, w_008_281, w_008_282, w_008_283, w_008_284, w_008_285, w_008_287, w_008_288, w_008_289, w_008_290, w_008_291, w_008_292, w_008_295, w_008_298, w_008_299, w_008_300, w_008_301, w_008_302, w_008_304, w_008_307, w_008_309, w_008_310, w_008_312, w_008_314, w_008_315, w_008_316, w_008_317, w_008_318, w_008_319, w_008_320, w_008_322, w_008_325, w_008_327, w_008_329, w_008_331, w_008_332, w_008_333, w_008_334, w_008_335, w_008_336, w_008_337, w_008_338, w_008_339, w_008_341, w_008_342, w_008_343, w_008_344, w_008_345, w_008_346, w_008_347, w_008_348, w_008_349, w_008_350, w_008_351, w_008_352, w_008_353, w_008_354, w_008_355, w_008_356, w_008_357, w_008_358, w_008_360, w_008_361, w_008_362, w_008_364, w_008_366, w_008_367, w_008_370, w_008_371, w_008_374, w_008_376, w_008_377, w_008_378, w_008_381, w_008_382, w_008_383, w_008_384, w_008_386, w_008_387, w_008_388, w_008_389, w_008_390, w_008_391, w_008_394, w_008_396, w_008_397, w_008_398, w_008_399, w_008_402, w_008_403, w_008_404, w_008_405, w_008_407, w_008_408, w_008_409, w_008_411, w_008_413, w_008_414, w_008_416, w_008_417, w_008_418, w_008_419, w_008_420, w_008_421, w_008_423, w_008_424, w_008_425, w_008_426, w_008_428, w_008_429, w_008_431, w_008_432, w_008_433, w_008_434, w_008_435, w_008_436, w_008_437, w_008_439, w_008_441, w_008_442, w_008_444, w_008_446, w_008_449, w_008_453, w_008_454, w_008_457, w_008_459, w_008_460, w_008_461, w_008_463, w_008_466, w_008_467, w_008_468, w_008_469, w_008_471, w_008_472, w_008_473, w_008_474, w_008_475, w_008_477, w_008_478, w_008_479, w_008_480, w_008_482, w_008_483, w_008_484, w_008_485, w_008_486, w_008_487, w_008_488, w_008_489, w_008_490, w_008_493, w_008_494, w_008_495, w_008_496, w_008_498, w_008_499, w_008_501, w_008_502, w_008_504, w_008_505, w_008_506, w_008_509, w_008_510, w_008_511, w_008_514, w_008_515, w_008_516, w_008_517, w_008_518, w_008_519, w_008_520, w_008_521, w_008_522, w_008_523, w_008_524, w_008_525, w_008_526, w_008_528, w_008_530, w_008_533, w_008_534, w_008_535, w_008_538, w_008_539, w_008_541, w_008_543, w_008_544, w_008_545, w_008_548, w_008_550, w_008_552, w_008_553, w_008_555, w_008_556, w_008_557, w_008_558, w_008_559, w_008_560, w_008_561, w_008_562, w_008_563, w_008_565, w_008_566, w_008_567, w_008_568, w_008_569, w_008_571, w_008_572, w_008_573, w_008_574, w_008_575, w_008_576, w_008_577, w_008_580, w_008_581, w_008_582, w_008_583, w_008_584, w_008_585, w_008_587, w_008_588, w_008_589, w_008_590, w_008_591, w_008_592, w_008_594, w_008_595, w_008_598, w_008_601, w_008_602, w_008_603, w_008_604, w_008_605, w_008_608, w_008_610, w_008_611, w_008_612, w_008_613, w_008_614, w_008_615, w_008_616, w_008_619, w_008_620, w_008_621, w_008_622, w_008_623, w_008_624, w_008_625, w_008_626, w_008_628, w_008_629, w_008_636, w_008_637, w_008_638, w_008_639, w_008_640, w_008_644, w_008_645, w_008_646, w_008_647, w_008_648, w_008_650, w_008_651, w_008_653, w_008_654, w_008_656, w_008_657, w_008_658, w_008_659, w_008_661, w_008_662, w_008_663, w_008_664, w_008_665, w_008_666, w_008_668, w_008_669, w_008_674, w_008_676, w_008_677, w_008_678, w_008_679, w_008_680, w_008_681, w_008_682, w_008_683, w_008_685, w_008_686, w_008_688, w_008_692, w_008_693, w_008_694, w_008_696, w_008_697, w_008_698, w_008_699, w_008_700, w_008_701, w_008_702, w_008_703, w_008_704, w_008_707, w_008_708, w_008_709, w_008_710, w_008_711, w_008_713, w_008_714, w_008_715, w_008_718, w_008_719, w_008_720, w_008_721, w_008_722, w_008_724, w_008_725, w_008_726, w_008_727, w_008_728, w_008_729, w_008_730, w_008_733, w_008_735, w_008_737, w_008_738, w_008_740, w_008_742, w_008_743, w_008_745, w_008_746, w_008_747, w_008_748, w_008_749, w_008_750, w_008_751, w_008_753, w_008_755, w_008_757, w_008_758, w_008_760, w_008_762, w_008_763, w_008_767, w_008_768, w_008_769, w_008_770, w_008_771, w_008_772, w_008_773, w_008_777, w_008_778, w_008_779, w_008_780, w_008_781, w_008_782, w_008_783, w_008_784, w_008_786;
  wire w_009_000, w_009_001, w_009_003, w_009_004, w_009_005, w_009_006, w_009_007, w_009_009, w_009_010, w_009_011, w_009_012, w_009_013, w_009_014, w_009_015, w_009_016, w_009_017, w_009_018, w_009_019, w_009_020, w_009_021, w_009_022, w_009_023, w_009_024, w_009_025, w_009_026, w_009_027, w_009_028, w_009_029, w_009_030, w_009_031, w_009_032, w_009_033, w_009_035, w_009_036, w_009_037, w_009_038, w_009_040, w_009_041, w_009_042, w_009_043, w_009_044, w_009_045, w_009_046, w_009_047, w_009_048, w_009_049, w_009_050, w_009_051, w_009_052, w_009_053, w_009_054, w_009_055, w_009_056, w_009_058, w_009_059, w_009_060, w_009_061, w_009_062, w_009_064, w_009_065, w_009_066, w_009_068, w_009_070, w_009_071, w_009_072, w_009_073, w_009_074, w_009_075, w_009_076, w_009_077, w_009_078, w_009_079, w_009_080, w_009_081, w_009_082, w_009_083, w_009_084, w_009_085, w_009_086, w_009_087, w_009_088, w_009_089, w_009_090, w_009_091, w_009_092, w_009_093, w_009_094, w_009_095, w_009_096, w_009_097, w_009_098, w_009_099, w_009_100, w_009_101, w_009_102, w_009_103, w_009_104, w_009_105, w_009_106, w_009_107, w_009_108, w_009_109, w_009_110, w_009_111, w_009_113, w_009_114, w_009_115, w_009_116, w_009_117, w_009_118, w_009_119, w_009_120, w_009_121, w_009_122, w_009_123, w_009_124, w_009_125, w_009_126, w_009_127, w_009_128, w_009_129, w_009_130, w_009_131, w_009_132, w_009_133, w_009_134, w_009_135, w_009_136, w_009_137, w_009_138, w_009_139, w_009_140, w_009_141, w_009_142, w_009_143, w_009_144, w_009_145, w_009_146, w_009_147, w_009_149, w_009_150, w_009_151, w_009_152, w_009_153, w_009_154, w_009_155, w_009_156, w_009_158, w_009_159, w_009_160, w_009_161, w_009_162, w_009_163, w_009_164, w_009_166, w_009_167, w_009_168, w_009_169, w_009_172, w_009_173, w_009_175, w_009_176, w_009_177, w_009_180, w_009_181, w_009_182, w_009_183, w_009_184, w_009_185, w_009_186, w_009_189, w_009_190, w_009_191, w_009_193, w_009_194, w_009_196, w_009_197, w_009_198, w_009_199, w_009_200, w_009_208, w_009_209, w_009_210, w_009_211, w_009_213, w_009_214, w_009_215, w_009_216, w_009_217, w_009_219, w_009_220, w_009_221, w_009_222, w_009_223, w_009_224, w_009_226, w_009_228, w_009_229, w_009_230, w_009_231, w_009_232, w_009_233, w_009_234, w_009_235, w_009_236, w_009_237, w_009_238, w_009_239, w_009_240, w_009_241, w_009_243, w_009_244, w_009_245, w_009_246, w_009_247, w_009_248, w_009_249, w_009_250, w_009_251, w_009_253, w_009_255, w_009_258, w_009_259, w_009_260, w_009_264, w_009_265, w_009_267, w_009_268, w_009_270, w_009_271, w_009_272, w_009_273, w_009_274, w_009_279, w_009_281, w_009_283, w_009_284, w_009_288, w_009_293, w_009_294, w_009_295, w_009_296, w_009_297, w_009_300, w_009_301, w_009_302, w_009_303, w_009_305, w_009_308, w_009_310, w_009_313, w_009_314, w_009_315, w_009_316, w_009_317, w_009_318, w_009_320, w_009_321, w_009_322, w_009_325, w_009_326, w_009_328, w_009_329, w_009_330, w_009_331, w_009_333, w_009_335, w_009_336, w_009_337, w_009_338, w_009_340, w_009_341, w_009_342, w_009_343, w_009_344, w_009_345, w_009_350, w_009_351, w_009_353, w_009_354, w_009_357, w_009_359, w_009_360, w_009_361, w_009_362, w_009_363, w_009_364, w_009_365, w_009_366, w_009_368, w_009_369, w_009_370, w_009_371, w_009_372, w_009_373, w_009_374, w_009_375, w_009_376, w_009_377, w_009_378, w_009_379, w_009_380, w_009_382, w_009_383, w_009_384, w_009_388, w_009_389, w_009_390, w_009_391, w_009_392, w_009_393, w_009_394, w_009_395, w_009_396, w_009_397, w_009_398, w_009_399, w_009_402, w_009_403, w_009_404, w_009_405, w_009_406, w_009_407, w_009_408, w_009_411, w_009_412, w_009_414, w_009_415, w_009_416, w_009_417, w_009_418, w_009_420, w_009_421, w_009_422, w_009_423, w_009_424, w_009_426, w_009_427, w_009_428, w_009_430, w_009_432, w_009_433, w_009_435, w_009_438, w_009_439, w_009_440, w_009_441, w_009_442, w_009_443, w_009_444, w_009_445, w_009_446, w_009_448, w_009_449, w_009_451, w_009_452, w_009_455, w_009_456, w_009_460, w_009_462, w_009_463, w_009_464, w_009_465, w_009_468, w_009_469, w_009_470, w_009_471, w_009_472, w_009_473, w_009_476, w_009_478, w_009_479, w_009_480, w_009_481, w_009_482, w_009_483, w_009_485, w_009_486, w_009_487, w_009_488, w_009_489, w_009_490, w_009_491, w_009_492, w_009_493, w_009_497, w_009_498, w_009_499, w_009_500, w_009_501, w_009_502, w_009_503, w_009_504, w_009_505, w_009_507, w_009_508, w_009_509, w_009_510, w_009_512, w_009_513, w_009_515, w_009_516, w_009_517, w_009_520, w_009_521, w_009_522, w_009_523, w_009_524, w_009_525, w_009_527, w_009_528, w_009_529, w_009_531, w_009_532, w_009_533, w_009_536, w_009_537, w_009_539, w_009_540, w_009_541, w_009_542, w_009_543, w_009_545, w_009_546, w_009_547, w_009_549, w_009_550, w_009_551, w_009_552, w_009_553, w_009_554, w_009_555, w_009_556, w_009_557, w_009_558, w_009_560, w_009_561, w_009_562, w_009_563, w_009_564, w_009_568, w_009_570, w_009_571, w_009_572, w_009_573, w_009_574, w_009_579, w_009_581, w_009_583, w_009_584, w_009_591, w_009_594, w_009_597, w_009_598, w_009_600, w_009_601, w_009_602, w_009_603, w_009_604, w_009_606, w_009_607, w_009_609, w_009_610, w_009_611, w_009_612, w_009_614, w_009_616, w_009_619, w_009_621, w_009_623, w_009_625, w_009_626, w_009_627, w_009_628, w_009_629, w_009_631, w_009_632, w_009_633, w_009_634, w_009_635, w_009_636, w_009_637, w_009_638, w_009_642, w_009_643, w_009_644, w_009_645, w_009_646, w_009_647, w_009_648, w_009_649, w_009_650, w_009_651, w_009_652, w_009_654;
  wire w_010_000, w_010_002, w_010_003, w_010_004, w_010_005, w_010_006, w_010_008, w_010_009, w_010_010, w_010_011, w_010_012, w_010_013, w_010_014, w_010_016, w_010_017, w_010_018, w_010_020, w_010_021, w_010_027, w_010_031, w_010_032, w_010_036, w_010_039, w_010_042, w_010_043, w_010_045, w_010_049, w_010_050, w_010_051, w_010_053, w_010_054, w_010_056, w_010_057, w_010_058, w_010_059, w_010_060, w_010_061, w_010_064, w_010_067, w_010_070, w_010_073, w_010_074, w_010_076, w_010_077, w_010_078, w_010_080, w_010_083, w_010_084, w_010_085, w_010_086, w_010_087, w_010_088, w_010_089, w_010_091, w_010_094, w_010_095, w_010_097, w_010_099, w_010_102, w_010_105, w_010_106, w_010_107, w_010_108, w_010_109, w_010_113, w_010_114, w_010_117, w_010_118, w_010_119, w_010_120, w_010_121, w_010_122, w_010_123, w_010_124, w_010_125, w_010_126, w_010_127, w_010_128, w_010_129, w_010_130, w_010_131, w_010_133, w_010_134, w_010_135, w_010_136, w_010_139, w_010_140, w_010_144, w_010_145, w_010_147, w_010_148, w_010_149, w_010_151, w_010_154, w_010_155, w_010_156, w_010_157, w_010_158, w_010_159, w_010_161, w_010_162, w_010_163, w_010_164, w_010_165, w_010_166, w_010_168, w_010_169, w_010_172, w_010_174, w_010_177, w_010_178, w_010_179, w_010_181, w_010_183, w_010_185, w_010_186, w_010_187, w_010_188, w_010_190, w_010_191, w_010_192, w_010_193, w_010_194, w_010_196, w_010_197, w_010_199, w_010_201, w_010_204, w_010_205, w_010_207, w_010_209, w_010_210, w_010_211, w_010_213, w_010_216, w_010_217, w_010_218, w_010_219, w_010_220, w_010_221, w_010_222, w_010_224, w_010_225, w_010_226, w_010_227, w_010_228, w_010_229, w_010_230, w_010_232, w_010_233, w_010_235, w_010_236, w_010_238, w_010_240, w_010_241, w_010_242, w_010_243, w_010_245, w_010_248, w_010_249, w_010_250, w_010_255, w_010_258, w_010_259, w_010_260, w_010_261, w_010_263, w_010_264, w_010_265, w_010_268, w_010_269, w_010_270, w_010_272, w_010_275, w_010_276, w_010_277, w_010_278, w_010_280, w_010_282, w_010_283, w_010_285, w_010_286, w_010_288, w_010_289, w_010_290, w_010_291, w_010_295, w_010_298, w_010_300, w_010_301, w_010_303, w_010_306, w_010_308, w_010_311, w_010_312, w_010_313, w_010_314, w_010_315, w_010_317, w_010_319, w_010_321, w_010_322, w_010_326, w_010_327, w_010_328, w_010_331, w_010_335, w_010_338, w_010_339, w_010_341, w_010_342, w_010_343, w_010_347, w_010_348, w_010_349, w_010_350, w_010_351, w_010_352, w_010_353, w_010_354, w_010_355, w_010_356, w_010_357, w_010_358, w_010_359, w_010_360, w_010_361, w_010_362, w_010_364, w_010_365, w_010_368, w_010_369, w_010_370, w_010_373, w_010_375, w_010_377, w_010_381, w_010_382, w_010_383, w_010_384, w_010_385, w_010_386, w_010_387, w_010_388, w_010_395, w_010_396, w_010_397, w_010_398, w_010_399, w_010_400, w_010_403, w_010_405, w_010_406, w_010_407, w_010_408, w_010_412, w_010_413, w_010_414, w_010_415, w_010_416, w_010_417, w_010_418, w_010_419, w_010_420, w_010_421, w_010_423, w_010_425, w_010_426, w_010_427, w_010_428, w_010_429, w_010_431, w_010_432, w_010_434, w_010_437, w_010_441, w_010_442, w_010_443, w_010_444, w_010_446, w_010_447, w_010_449, w_010_450, w_010_451, w_010_452, w_010_453, w_010_454, w_010_455, w_010_456, w_010_457, w_010_458, w_010_459, w_010_460, w_010_466, w_010_467, w_010_468, w_010_471, w_010_472, w_010_476, w_010_478, w_010_479, w_010_481, w_010_482, w_010_484, w_010_486, w_010_487, w_010_488, w_010_489, w_010_491, w_010_494, w_010_496, w_010_497, w_010_498, w_010_499, w_010_500, w_010_505, w_010_506, w_010_507, w_010_510, w_010_511, w_010_513, w_010_514, w_010_515, w_010_516, w_010_517, w_010_518, w_010_519, w_010_520, w_010_522, w_010_525, w_010_526, w_010_528, w_010_529, w_010_530, w_010_531, w_010_532, w_010_533, w_010_539, w_010_540, w_010_542, w_010_544, w_010_548, w_010_550, w_010_551, w_010_553, w_010_554, w_010_556, w_010_558, w_010_559, w_010_560, w_010_561, w_010_563, w_010_564, w_010_565, w_010_566, w_010_567, w_010_568, w_010_569, w_010_570, w_010_571, w_010_576, w_010_577, w_010_579, w_010_580, w_010_581, w_010_583, w_010_584, w_010_585, w_010_586, w_010_587, w_010_588, w_010_589, w_010_591, w_010_592, w_010_593, w_010_595, w_010_596, w_010_597, w_010_598, w_010_599, w_010_603, w_010_604, w_010_606, w_010_609, w_010_610, w_010_611, w_010_612, w_010_613, w_010_614, w_010_616, w_010_618, w_010_619, w_010_622, w_010_623, w_010_625, w_010_626, w_010_627, w_010_628, w_010_631, w_010_632, w_010_633, w_010_635, w_010_638, w_010_640, w_010_641, w_010_642, w_010_644, w_010_645, w_010_646, w_010_649, w_010_653, w_010_655, w_010_656, w_010_659, w_010_660, w_010_661, w_010_663, w_010_667, w_010_668, w_010_669, w_010_670, w_010_672, w_010_673, w_010_674, w_010_675, w_010_677, w_010_678, w_010_679, w_010_680, w_010_681, w_010_682, w_010_684, w_010_685, w_010_686, w_010_688, w_010_691, w_010_692, w_010_695, w_010_697, w_010_698, w_010_700, w_010_703, w_010_705, w_010_707, w_010_709, w_010_711, w_010_712, w_010_713, w_010_714, w_010_715, w_010_716, w_010_717, w_010_718, w_010_719, w_010_720, w_010_721, w_010_722, w_010_724, w_010_726, w_010_731, w_010_732, w_010_733, w_010_735, w_010_736, w_010_737, w_010_739, w_010_742, w_010_743, w_010_745, w_010_746, w_010_747, w_010_748, w_010_749, w_010_750, w_010_751, w_010_753, w_010_754, w_010_756, w_010_757, w_010_758, w_010_759, w_010_760, w_010_763, w_010_765, w_010_766, w_010_767, w_010_768, w_010_769, w_010_770, w_010_773, w_010_775, w_010_777, w_010_779;
  wire w_011_001, w_011_002, w_011_003, w_011_004, w_011_005, w_011_006, w_011_007, w_011_009, w_011_010, w_011_011, w_011_013, w_011_014, w_011_015, w_011_016, w_011_017, w_011_018, w_011_020, w_011_021, w_011_022, w_011_023, w_011_024, w_011_025, w_011_026, w_011_027, w_011_028, w_011_030, w_011_031, w_011_032, w_011_033, w_011_035, w_011_036, w_011_037, w_011_039, w_011_041, w_011_042, w_011_043, w_011_044, w_011_045, w_011_046, w_011_047, w_011_048, w_011_049, w_011_050, w_011_051, w_011_052, w_011_054, w_011_056, w_011_057, w_011_058, w_011_059, w_011_060, w_011_061, w_011_062, w_011_063, w_011_064, w_011_066, w_011_069, w_011_070, w_011_071, w_011_072, w_011_073, w_011_075, w_011_077, w_011_078, w_011_079, w_011_080, w_011_081, w_011_082, w_011_083, w_011_084, w_011_085, w_011_086, w_011_087, w_011_088, w_011_089, w_011_090, w_011_092, w_011_093, w_011_094, w_011_095, w_011_096, w_011_097, w_011_098, w_011_099, w_011_102, w_011_103, w_011_104, w_011_108, w_011_109, w_011_110, w_011_111, w_011_112, w_011_113, w_011_114, w_011_116, w_011_117, w_011_118, w_011_119, w_011_120, w_011_121, w_011_123, w_011_124, w_011_125, w_011_126, w_011_127, w_011_128, w_011_130, w_011_131, w_011_132, w_011_133, w_011_134, w_011_135, w_011_136, w_011_137, w_011_138, w_011_139, w_011_140, w_011_141, w_011_142, w_011_143, w_011_144, w_011_146, w_011_147, w_011_148, w_011_149, w_011_150, w_011_151, w_011_152, w_011_154, w_011_155, w_011_156, w_011_157, w_011_158, w_011_159, w_011_160, w_011_162, w_011_163, w_011_164, w_011_166, w_011_167, w_011_168, w_011_169, w_011_170, w_011_172, w_011_173, w_011_174, w_011_175, w_011_176, w_011_177, w_011_179, w_011_180, w_011_181, w_011_182, w_011_187, w_011_188, w_011_189, w_011_190, w_011_191, w_011_193, w_011_194, w_011_195, w_011_196, w_011_197, w_011_198, w_011_199, w_011_201, w_011_202, w_011_203, w_011_204, w_011_205, w_011_206, w_011_208, w_011_209, w_011_210, w_011_211, w_011_213, w_011_214, w_011_215, w_011_216, w_011_217, w_011_219, w_011_220, w_011_222, w_011_224, w_011_227, w_011_228, w_011_229, w_011_231, w_011_232, w_011_233, w_011_235, w_011_236, w_011_237, w_011_239, w_011_240, w_011_242, w_011_243, w_011_244, w_011_248, w_011_249, w_011_251, w_011_253, w_011_257, w_011_260, w_011_262, w_011_263, w_011_265, w_011_267, w_011_268, w_011_269, w_011_270, w_011_271, w_011_273, w_011_276, w_011_278, w_011_279, w_011_280, w_011_281, w_011_284, w_011_286, w_011_288, w_011_289, w_011_290, w_011_291, w_011_295, w_011_298, w_011_300, w_011_301, w_011_302, w_011_303, w_011_306, w_011_308, w_011_309, w_011_310, w_011_312, w_011_315, w_011_317, w_011_319, w_011_320, w_011_321, w_011_322, w_011_324, w_011_325, w_011_328, w_011_329, w_011_330, w_011_332, w_011_333, w_011_334, w_011_336, w_011_337, w_011_338, w_011_339, w_011_341, w_011_342, w_011_343, w_011_344, w_011_345, w_011_347, w_011_350, w_011_351, w_011_352, w_011_353, w_011_356, w_011_357, w_011_359, w_011_360, w_011_361, w_011_364, w_011_365, w_011_366, w_011_367, w_011_368, w_011_371, w_011_372, w_011_373, w_011_374, w_011_378, w_011_379, w_011_383, w_011_384, w_011_385, w_011_387, w_011_390, w_011_391, w_011_392, w_011_393, w_011_396, w_011_397, w_011_398, w_011_401, w_011_405, w_011_406, w_011_407, w_011_409, w_011_410, w_011_411, w_011_414, w_011_416, w_011_419, w_011_420, w_011_421, w_011_424, w_011_426, w_011_427, w_011_428, w_011_430, w_011_431, w_011_433, w_011_435, w_011_437, w_011_438, w_011_439, w_011_440, w_011_441, w_011_443, w_011_444, w_011_446, w_011_450, w_011_455, w_011_457, w_011_458, w_011_459, w_011_460, w_011_461, w_011_462, w_011_463, w_011_465, w_011_466, w_011_467, w_011_468, w_011_469, w_011_471, w_011_472, w_011_473, w_011_474, w_011_477, w_011_480, w_011_481, w_011_486, w_011_489, w_011_490, w_011_491, w_011_492, w_011_494, w_011_500, w_011_502, w_011_503, w_011_504, w_011_508, w_011_510, w_011_511, w_011_512, w_011_514, w_011_515, w_011_517, w_011_519, w_011_520, w_011_521, w_011_523, w_011_525, w_011_527, w_011_529, w_011_530, w_011_531, w_011_532, w_011_533, w_011_538, w_011_539, w_011_540, w_011_541, w_011_542, w_011_543, w_011_544, w_011_545, w_011_546, w_011_548, w_011_549, w_011_550, w_011_551, w_011_554, w_011_555, w_011_556, w_011_557, w_011_558, w_011_559, w_011_560, w_011_561, w_011_562, w_011_563, w_011_564, w_011_565, w_011_566, w_011_567, w_011_568, w_011_569, w_011_570, w_011_571, w_011_572, w_011_575, w_011_576, w_011_579, w_011_582, w_011_583, w_011_586, w_011_587, w_011_589, w_011_591, w_011_592, w_011_594, w_011_596, w_011_597, w_011_599, w_011_603, w_011_605, w_011_606, w_011_607, w_011_611, w_011_615, w_011_616, w_011_617, w_011_618, w_011_620, w_011_622, w_011_624, w_011_626, w_011_629, w_011_630, w_011_631, w_011_632, w_011_633, w_011_634, w_011_635, w_011_637, w_011_639, w_011_641, w_011_642;
  wire w_012_000, w_012_001, w_012_002, w_012_003, w_012_004, w_012_005, w_012_006, w_012_007, w_012_008, w_012_009, w_012_010, w_012_011, w_012_012, w_012_013, w_012_015, w_012_016, w_012_017, w_012_018, w_012_019, w_012_020, w_012_021, w_012_022, w_012_023, w_012_024, w_012_025, w_012_026, w_012_027, w_012_028, w_012_029, w_012_030, w_012_031, w_012_032, w_012_033, w_012_034, w_012_035, w_012_036, w_012_037, w_012_038, w_012_039, w_012_040, w_012_041, w_012_042, w_012_043, w_012_044, w_012_045, w_012_046, w_012_047, w_012_048, w_012_049, w_012_050, w_012_051, w_012_052, w_012_053, w_012_054, w_012_055, w_012_056, w_012_057, w_012_058, w_012_059, w_012_060, w_012_061, w_012_062, w_012_063, w_012_065, w_012_066, w_012_067, w_012_068, w_012_069, w_012_070, w_012_071, w_012_072, w_012_073, w_012_074, w_012_075, w_012_076, w_012_077, w_012_078, w_012_079, w_012_080, w_012_081, w_012_082, w_012_083, w_012_084, w_012_086, w_012_087, w_012_088, w_012_089, w_012_090, w_012_091, w_012_092, w_012_093, w_012_094, w_012_095, w_012_096, w_012_098, w_012_099, w_012_101, w_012_102, w_012_103, w_012_104, w_012_105, w_012_106, w_012_107, w_012_108, w_012_109, w_012_110, w_012_111, w_012_112, w_012_113, w_012_114, w_012_115, w_012_116, w_012_118, w_012_119, w_012_120, w_012_121, w_012_122, w_012_123, w_012_124, w_012_125, w_012_126, w_012_127, w_012_129, w_012_130, w_012_131, w_012_132, w_012_134, w_012_135, w_012_136, w_012_137, w_012_138, w_012_140, w_012_141, w_012_142, w_012_143, w_012_145, w_012_147, w_012_149, w_012_150, w_012_151, w_012_152, w_012_153, w_012_154, w_012_155, w_012_157, w_012_158, w_012_162, w_012_163, w_012_164, w_012_165, w_012_167, w_012_168, w_012_169, w_012_170, w_012_171, w_012_172, w_012_174, w_012_175, w_012_176, w_012_177, w_012_178, w_012_179, w_012_181, w_012_182, w_012_183, w_012_185, w_012_187, w_012_188, w_012_189, w_012_190, w_012_191, w_012_192, w_012_193, w_012_194, w_012_198, w_012_199, w_012_200, w_012_201, w_012_202, w_012_203, w_012_204, w_012_205, w_012_206, w_012_207, w_012_208, w_012_209, w_012_210, w_012_211, w_012_212, w_012_213, w_012_214, w_012_215, w_012_216, w_012_217, w_012_219, w_012_221, w_012_223, w_012_224, w_012_225, w_012_226, w_012_227, w_012_228, w_012_229, w_012_230, w_012_231, w_012_232, w_012_233, w_012_234, w_012_235, w_012_236, w_012_237, w_012_238, w_012_239, w_012_240, w_012_241, w_012_242, w_012_243, w_012_244, w_012_245, w_012_246, w_012_247, w_012_249, w_012_250, w_012_252, w_012_253, w_012_254, w_012_255, w_012_256, w_012_257, w_012_258, w_012_259, w_012_260, w_012_261, w_012_262, w_012_263, w_012_264, w_012_267, w_012_268, w_012_269, w_012_270, w_012_271, w_012_272, w_012_273, w_012_274, w_012_275, w_012_276, w_012_277, w_012_278, w_012_279, w_012_281, w_012_282, w_012_285, w_012_286, w_012_287, w_012_288, w_012_289, w_012_290, w_012_291, w_012_292, w_012_293, w_012_294, w_012_295, w_012_296, w_012_297, w_012_298, w_012_299, w_012_300, w_012_301, w_012_302, w_012_303, w_012_304, w_012_305, w_012_306, w_012_308, w_012_309, w_012_310, w_012_311, w_012_312, w_012_313, w_012_314, w_012_315, w_012_316, w_012_317, w_012_319, w_012_320, w_012_321, w_012_322, w_012_323, w_012_324, w_012_325, w_012_327, w_012_328, w_012_330, w_012_331, w_012_332, w_012_333, w_012_335, w_012_336, w_012_337, w_012_338, w_012_340, w_012_342, w_012_344, w_012_345, w_012_346, w_012_347, w_012_348, w_012_350;
  wire w_013_000, w_013_001, w_013_002, w_013_003, w_013_004, w_013_005, w_013_006, w_013_008, w_013_009, w_013_010, w_013_011, w_013_012, w_013_013, w_013_015, w_013_016, w_013_017, w_013_020, w_013_021, w_013_022, w_013_023, w_013_024, w_013_025, w_013_026, w_013_027, w_013_028, w_013_029, w_013_030, w_013_031, w_013_032, w_013_034, w_013_035, w_013_036, w_013_037, w_013_040, w_013_041, w_013_042, w_013_043, w_013_044, w_013_046, w_013_047, w_013_048, w_013_049, w_013_050, w_013_053, w_013_054, w_013_055, w_013_059, w_013_060, w_013_061, w_013_062, w_013_063, w_013_064, w_013_065, w_013_066, w_013_067, w_013_068, w_013_069, w_013_070, w_013_071, w_013_072, w_013_073, w_013_074, w_013_075, w_013_076, w_013_077, w_013_078, w_013_079, w_013_080, w_013_081, w_013_083, w_013_086, w_013_087, w_013_088, w_013_089, w_013_090, w_013_091, w_013_092, w_013_093, w_013_095, w_013_096, w_013_097, w_013_098, w_013_099, w_013_100, w_013_102, w_013_103, w_013_104, w_013_105, w_013_106, w_013_107, w_013_108, w_013_109, w_013_110, w_013_111, w_013_112, w_013_114, w_013_115, w_013_116, w_013_117, w_013_118, w_013_121, w_013_122, w_013_123, w_013_124, w_013_125, w_013_126, w_013_127, w_013_128, w_013_129, w_013_130, w_013_131, w_013_132, w_013_133, w_013_134, w_013_135, w_013_136, w_013_137, w_013_138, w_013_139, w_013_140, w_013_141, w_013_142, w_013_144, w_013_145, w_013_146, w_013_147, w_013_148, w_013_150, w_013_151, w_013_153, w_013_154, w_013_155, w_013_156, w_013_157, w_013_158, w_013_159, w_013_160, w_013_161, w_013_162, w_013_163, w_013_164, w_013_165, w_013_166, w_013_168, w_013_169, w_013_170, w_013_171, w_013_172, w_013_174, w_013_175, w_013_176, w_013_178, w_013_179, w_013_180, w_013_181, w_013_183, w_013_184, w_013_185, w_013_186, w_013_188, w_013_189, w_013_190, w_013_191, w_013_194, w_013_195, w_013_197, w_013_199, w_013_200, w_013_201, w_013_202, w_013_203, w_013_204, w_013_205, w_013_206, w_013_207, w_013_208, w_013_209, w_013_210, w_013_211, w_013_214, w_013_215, w_013_217, w_013_218, w_013_219, w_013_220, w_013_222, w_013_224, w_013_229, w_013_230, w_013_232, w_013_235, w_013_236, w_013_237, w_013_239, w_013_242, w_013_243, w_013_246, w_013_249, w_013_251, w_013_256, w_013_257, w_013_258, w_013_259, w_013_260, w_013_263, w_013_265, w_013_266, w_013_269, w_013_270, w_013_272, w_013_274, w_013_275, w_013_278, w_013_279, w_013_284, w_013_286, w_013_288, w_013_290, w_013_292, w_013_293, w_013_295, w_013_296, w_013_297, w_013_301, w_013_302, w_013_303, w_013_305, w_013_306, w_013_307, w_013_309, w_013_311, w_013_313, w_013_316, w_013_317, w_013_318, w_013_320, w_013_321, w_013_322, w_013_323, w_013_326, w_013_327, w_013_329, w_013_330, w_013_331, w_013_332, w_013_334, w_013_339, w_013_340, w_013_344, w_013_346, w_013_348, w_013_349, w_013_352, w_013_353, w_013_357, w_013_358, w_013_359, w_013_361, w_013_363, w_013_367, w_013_369, w_013_370, w_013_371, w_013_372, w_013_373, w_013_374, w_013_376, w_013_379, w_013_380, w_013_382, w_013_385, w_013_386, w_013_391, w_013_392, w_013_394, w_013_396, w_013_397, w_013_399, w_013_400, w_013_401, w_013_403, w_013_404, w_013_407, w_013_408, w_013_409, w_013_411, w_013_412, w_013_413, w_013_414, w_013_415, w_013_416, w_013_418, w_013_419, w_013_422, w_013_426, w_013_428, w_013_429, w_013_431, w_013_432, w_013_436, w_013_437, w_013_439, w_013_442, w_013_443, w_013_444, w_013_445, w_013_446, w_013_447, w_013_448, w_013_452, w_013_453, w_013_455, w_013_458, w_013_461, w_013_462, w_013_463, w_013_464, w_013_466, w_013_467, w_013_468, w_013_469, w_013_470, w_013_471, w_013_478, w_013_479, w_013_484, w_013_489, w_013_494, w_013_496, w_013_501, w_013_506, w_013_507, w_013_509, w_013_510, w_013_511, w_013_514, w_013_515, w_013_517, w_013_518, w_013_519, w_013_520, w_013_521, w_013_522, w_013_523, w_013_524, w_013_526, w_013_527, w_013_528, w_013_529, w_013_530, w_013_534, w_013_536, w_013_538, w_013_539, w_013_540, w_013_541, w_013_542, w_013_543, w_013_544, w_013_545, w_013_546, w_013_548, w_013_551, w_013_552, w_013_555, w_013_556, w_013_558, w_013_559, w_013_560, w_013_561, w_013_562, w_013_563, w_013_564, w_013_565, w_013_570, w_013_571, w_013_572, w_013_573, w_013_574, w_013_575, w_013_576, w_013_578, w_013_582, w_013_583, w_013_585, w_013_586, w_013_587, w_013_588, w_013_589, w_013_590, w_013_591, w_013_592, w_013_593, w_013_594, w_013_595, w_013_596;
  wire w_014_000, w_014_001, w_014_002, w_014_003, w_014_004, w_014_005, w_014_007, w_014_008, w_014_009, w_014_010, w_014_011, w_014_012, w_014_013, w_014_014, w_014_015, w_014_016, w_014_017, w_014_018, w_014_019, w_014_021, w_014_022, w_014_023, w_014_024, w_014_025, w_014_026, w_014_027, w_014_028, w_014_029, w_014_030, w_014_031, w_014_032, w_014_034, w_014_035, w_014_036, w_014_037, w_014_039, w_014_040, w_014_041, w_014_042, w_014_043, w_014_044, w_014_045, w_014_046, w_014_047, w_014_048, w_014_049, w_014_050, w_014_052, w_014_053, w_014_054, w_014_055, w_014_056, w_014_057, w_014_058, w_014_059, w_014_060, w_014_061, w_014_062, w_014_064, w_014_066, w_014_067, w_014_068, w_014_069, w_014_070, w_014_071, w_014_072, w_014_073, w_014_074, w_014_075, w_014_076, w_014_077, w_014_080, w_014_081, w_014_082, w_014_083, w_014_084, w_014_085, w_014_088, w_014_089, w_014_090, w_014_092, w_014_093, w_014_094, w_014_095, w_014_096, w_014_097, w_014_099, w_014_100, w_014_101, w_014_102, w_014_103, w_014_104, w_014_105, w_014_106, w_014_108, w_014_109, w_014_110, w_014_111, w_014_112, w_014_113, w_014_114, w_014_115, w_014_116, w_014_117, w_014_119, w_014_120, w_014_121, w_014_122, w_014_123, w_014_124, w_014_125, w_014_126, w_014_127, w_014_129, w_014_130, w_014_131, w_014_132, w_014_133, w_014_134, w_014_135, w_014_136, w_014_137, w_014_138, w_014_140, w_014_141, w_014_142, w_014_143, w_014_144, w_014_145, w_014_146, w_014_147, w_014_148, w_014_149, w_014_150, w_014_151, w_014_152, w_014_153, w_014_155, w_014_156, w_014_157, w_014_158, w_014_159, w_014_160, w_014_161, w_014_162, w_014_163, w_014_164, w_014_165, w_014_166, w_014_167, w_014_168, w_014_169, w_014_171, w_014_172, w_014_173, w_014_174, w_014_175, w_014_176, w_014_177, w_014_178, w_014_179, w_014_180, w_014_181, w_014_182, w_014_183, w_014_184, w_014_185, w_014_186, w_014_187, w_014_188, w_014_189, w_014_190, w_014_191, w_014_192, w_014_193, w_014_194, w_014_195, w_014_196, w_014_197, w_014_198, w_014_201, w_014_202, w_014_203, w_014_205, w_014_206, w_014_209, w_014_210, w_014_211, w_014_212, w_014_214, w_014_215, w_014_216, w_014_217, w_014_218, w_014_219, w_014_220, w_014_221, w_014_222, w_014_224, w_014_225, w_014_226, w_014_228, w_014_229, w_014_231, w_014_233, w_014_234, w_014_235, w_014_236, w_014_237, w_014_238, w_014_240, w_014_241, w_014_242, w_014_243, w_014_245, w_014_246, w_014_247, w_014_248, w_014_249, w_014_250, w_014_252, w_014_253, w_014_254, w_014_256, w_014_257, w_014_258, w_014_259, w_014_260, w_014_261, w_014_264, w_014_265, w_014_266, w_014_267, w_014_268, w_014_269, w_014_271, w_014_272, w_014_273, w_014_274, w_014_276, w_014_277, w_014_279, w_014_280, w_014_281, w_014_282, w_014_284, w_014_285, w_014_286, w_014_287, w_014_288, w_014_289, w_014_290, w_014_291, w_014_292, w_014_294, w_014_295;
  wire w_015_001, w_015_003, w_015_004, w_015_005, w_015_006, w_015_007, w_015_008, w_015_010, w_015_011, w_015_013, w_015_014, w_015_015, w_015_016, w_015_017, w_015_019, w_015_020, w_015_022, w_015_023, w_015_024, w_015_026, w_015_027, w_015_029, w_015_033, w_015_036, w_015_038, w_015_040, w_015_041, w_015_042, w_015_043, w_015_044, w_015_045, w_015_046, w_015_047, w_015_048, w_015_049, w_015_051, w_015_052, w_015_054, w_015_055, w_015_056, w_015_057, w_015_058, w_015_059, w_015_060, w_015_061, w_015_062, w_015_065, w_015_067, w_015_068, w_015_069, w_015_070, w_015_071, w_015_072, w_015_073, w_015_079, w_015_080, w_015_081, w_015_082, w_015_083, w_015_084, w_015_086, w_015_087, w_015_088, w_015_089, w_015_090, w_015_091, w_015_092, w_015_093, w_015_095, w_015_096, w_015_097, w_015_099, w_015_100, w_015_102, w_015_103, w_015_104, w_015_105, w_015_106, w_015_107, w_015_108, w_015_110, w_015_111, w_015_112, w_015_113, w_015_114, w_015_115, w_015_116, w_015_117, w_015_118, w_015_119, w_015_120, w_015_121, w_015_123, w_015_124, w_015_126, w_015_127, w_015_128, w_015_129, w_015_131, w_015_132, w_015_133, w_015_134, w_015_135, w_015_136, w_015_137, w_015_139, w_015_142, w_015_143, w_015_144, w_015_146, w_015_149, w_015_151, w_015_152, w_015_155, w_015_158, w_015_160, w_015_161, w_015_162, w_015_163, w_015_164, w_015_165, w_015_166, w_015_167, w_015_168, w_015_170, w_015_172, w_015_174, w_015_177, w_015_178, w_015_180, w_015_183, w_015_186, w_015_187, w_015_188, w_015_190, w_015_191, w_015_192, w_015_194, w_015_196, w_015_197, w_015_198, w_015_200, w_015_201, w_015_202, w_015_204, w_015_205, w_015_208, w_015_209, w_015_210, w_015_212, w_015_214, w_015_215, w_015_220, w_015_222, w_015_223, w_015_224, w_015_229, w_015_230, w_015_232, w_015_234, w_015_235, w_015_236, w_015_240, w_015_246, w_015_248, w_015_249, w_015_252, w_015_253, w_015_254, w_015_256, w_015_257, w_015_258, w_015_259, w_015_260, w_015_261, w_015_263, w_015_265, w_015_266, w_015_267, w_015_269, w_015_271, w_015_272, w_015_275, w_015_276, w_015_277, w_015_278, w_015_280, w_015_281, w_015_283, w_015_286, w_015_287, w_015_288, w_015_290, w_015_295, w_015_296, w_015_299, w_015_301, w_015_302, w_015_308, w_015_309, w_015_314, w_015_315, w_015_317, w_015_318, w_015_319, w_015_322, w_015_323, w_015_325, w_015_328, w_015_332, w_015_333, w_015_335, w_015_336, w_015_339, w_015_340, w_015_343, w_015_344, w_015_346, w_015_347, w_015_348, w_015_351, w_015_353, w_015_354, w_015_355, w_015_357, w_015_360, w_015_363, w_015_366, w_015_369, w_015_370, w_015_371, w_015_372, w_015_373, w_015_374, w_015_376, w_015_377, w_015_379, w_015_382, w_015_384, w_015_385, w_015_386, w_015_387, w_015_389, w_015_390, w_015_392, w_015_393, w_015_394, w_015_396, w_015_399, w_015_400, w_015_401, w_015_402, w_015_405, w_015_407, w_015_408, w_015_413, w_015_416, w_015_417, w_015_418, w_015_421, w_015_423, w_015_426, w_015_428, w_015_429, w_015_430, w_015_431, w_015_432, w_015_433, w_015_434, w_015_435, w_015_436, w_015_439, w_015_440, w_015_441, w_015_442, w_015_443, w_015_445, w_015_447, w_015_448, w_015_449, w_015_458, w_015_459, w_015_461, w_015_463, w_015_464, w_015_467, w_015_468, w_015_469, w_015_471, w_015_474, w_015_476, w_015_477, w_015_478, w_015_479, w_015_480, w_015_481, w_015_484, w_015_490, w_015_491, w_015_497, w_015_498, w_015_499, w_015_501, w_015_502, w_015_504, w_015_506, w_015_511, w_015_513, w_015_516, w_015_517, w_015_521, w_015_523, w_015_524, w_015_526, w_015_527, w_015_529, w_015_530, w_015_534, w_015_538, w_015_543, w_015_544, w_015_546, w_015_547, w_015_548, w_015_550, w_015_552, w_015_555, w_015_556, w_015_557, w_015_558, w_015_559, w_015_561, w_015_562, w_015_565, w_015_566, w_015_568, w_015_570, w_015_577, w_015_579, w_015_580, w_015_582, w_015_584, w_015_585, w_015_589, w_015_590, w_015_591, w_015_596, w_015_598, w_015_600, w_015_603, w_015_604, w_015_605, w_015_606, w_015_607, w_015_608, w_015_612, w_015_613, w_015_614, w_015_615, w_015_616, w_015_618, w_015_619, w_015_620, w_015_624, w_015_625, w_015_629, w_015_632, w_015_633, w_015_636, w_015_637, w_015_641, w_015_642, w_015_644, w_015_647, w_015_648, w_015_649, w_015_650, w_015_651, w_015_652, w_015_653, w_015_654, w_015_658, w_015_660, w_015_662, w_015_663, w_015_664, w_015_665, w_015_668, w_015_669, w_015_671, w_015_673, w_015_675, w_015_676, w_015_677;
  wire w_016_000, w_016_001, w_016_002, w_016_003, w_016_004, w_016_005, w_016_006, w_016_007, w_016_008;
  wire w_017_001, w_017_002, w_017_003, w_017_004, w_017_005, w_017_006, w_017_007, w_017_008, w_017_009, w_017_010, w_017_012, w_017_013, w_017_014, w_017_015, w_017_016, w_017_017, w_017_018, w_017_019, w_017_020, w_017_022, w_017_023, w_017_024, w_017_025, w_017_026, w_017_027, w_017_028, w_017_029, w_017_030, w_017_031, w_017_032, w_017_033, w_017_034, w_017_035, w_017_036, w_017_037, w_017_038, w_017_040, w_017_042, w_017_043, w_017_045, w_017_047, w_017_048, w_017_050, w_017_051, w_017_052, w_017_053, w_017_054, w_017_055, w_017_056, w_017_057, w_017_059, w_017_060, w_017_063, w_017_064, w_017_065, w_017_066, w_017_068, w_017_069, w_017_070, w_017_071, w_017_072, w_017_073, w_017_075, w_017_078, w_017_080, w_017_082, w_017_085, w_017_086, w_017_087, w_017_088, w_017_089, w_017_091, w_017_092, w_017_093, w_017_094, w_017_095, w_017_096, w_017_097, w_017_098, w_017_099, w_017_100, w_017_101, w_017_102, w_017_103, w_017_104, w_017_107, w_017_108, w_017_111, w_017_112, w_017_114, w_017_115, w_017_116, w_017_118, w_017_119, w_017_120, w_017_121, w_017_122, w_017_123, w_017_124, w_017_125, w_017_126, w_017_127, w_017_128, w_017_130, w_017_131, w_017_132, w_017_133, w_017_134, w_017_135, w_017_138, w_017_140, w_017_141, w_017_142, w_017_144, w_017_146, w_017_151, w_017_154, w_017_156, w_017_157, w_017_159, w_017_162, w_017_164, w_017_165, w_017_166, w_017_168, w_017_171, w_017_174, w_017_176, w_017_177, w_017_178, w_017_179, w_017_184, w_017_186, w_017_187, w_017_189, w_017_190, w_017_191, w_017_193, w_017_194, w_017_197, w_017_200, w_017_201, w_017_206, w_017_207, w_017_211, w_017_214, w_017_215, w_017_218, w_017_222, w_017_224, w_017_226, w_017_227, w_017_228, w_017_229, w_017_232, w_017_234, w_017_235, w_017_236, w_017_238, w_017_240, w_017_242, w_017_243, w_017_245, w_017_246, w_017_247, w_017_248, w_017_249, w_017_251, w_017_252, w_017_256, w_017_257, w_017_258, w_017_260, w_017_262, w_017_263, w_017_264, w_017_267, w_017_269, w_017_270, w_017_271, w_017_272, w_017_274, w_017_279, w_017_280, w_017_283, w_017_286, w_017_288, w_017_291, w_017_292, w_017_293, w_017_294, w_017_295, w_017_297, w_017_298, w_017_305, w_017_306, w_017_309, w_017_312, w_017_314, w_017_315, w_017_318, w_017_319, w_017_321, w_017_322, w_017_323, w_017_325, w_017_329, w_017_333, w_017_336, w_017_337, w_017_338, w_017_341, w_017_343, w_017_344, w_017_345, w_017_347, w_017_349, w_017_352, w_017_356, w_017_357, w_017_359, w_017_360, w_017_364, w_017_365, w_017_366, w_017_367, w_017_368, w_017_370, w_017_371, w_017_372, w_017_373, w_017_374, w_017_375, w_017_376, w_017_379, w_017_380, w_017_381, w_017_385, w_017_386, w_017_390, w_017_392, w_017_394, w_017_399, w_017_402, w_017_403, w_017_404, w_017_406, w_017_407, w_017_408, w_017_409, w_017_410, w_017_412, w_017_415, w_017_416, w_017_419, w_017_421, w_017_422, w_017_424, w_017_425, w_017_426, w_017_428, w_017_429, w_017_430, w_017_433, w_017_434, w_017_435, w_017_436, w_017_437, w_017_438, w_017_439, w_017_443, w_017_447, w_017_449, w_017_451, w_017_453, w_017_458, w_017_460, w_017_461, w_017_462, w_017_463, w_017_464, w_017_467, w_017_468, w_017_470, w_017_471, w_017_475, w_017_477, w_017_479, w_017_480, w_017_482, w_017_483, w_017_484, w_017_485, w_017_487, w_017_492, w_017_495, w_017_496, w_017_497, w_017_498, w_017_499, w_017_501, w_017_502, w_017_506, w_017_508, w_017_512, w_017_513, w_017_515, w_017_517, w_017_518, w_017_522, w_017_523, w_017_524, w_017_525, w_017_529, w_017_531, w_017_532, w_017_536, w_017_538, w_017_540, w_017_541, w_017_543, w_017_546, w_017_549, w_017_552, w_017_553, w_017_555, w_017_559, w_017_560, w_017_561, w_017_562, w_017_564, w_017_565, w_017_567, w_017_569, w_017_572, w_017_575, w_017_576, w_017_578, w_017_579, w_017_581, w_017_587, w_017_589, w_017_590, w_017_591, w_017_592, w_017_594, w_017_596, w_017_597, w_017_598, w_017_599, w_017_601, w_017_603, w_017_606, w_017_607, w_017_609, w_017_611, w_017_612, w_017_613, w_017_616, w_017_620, w_017_623, w_017_625, w_017_626, w_017_629, w_017_631, w_017_636, w_017_639, w_017_640, w_017_648, w_017_649, w_017_650, w_017_651, w_017_653, w_017_655, w_017_657, w_017_659, w_017_660, w_017_662, w_017_663, w_017_664, w_017_667, w_017_669, w_017_670;
  wire w_018_000, w_018_001, w_018_002, w_018_003, w_018_004, w_018_005, w_018_006, w_018_007, w_018_008, w_018_009, w_018_010, w_018_011, w_018_012, w_018_013, w_018_014, w_018_015, w_018_016, w_018_017, w_018_018, w_018_019, w_018_020, w_018_021, w_018_022, w_018_023, w_018_024, w_018_025, w_018_026, w_018_027, w_018_028, w_018_029, w_018_030, w_018_031, w_018_032, w_018_033, w_018_034, w_018_035, w_018_036, w_018_037, w_018_038, w_018_039, w_018_040, w_018_041, w_018_042, w_018_043, w_018_044;
  wire w_019_000, w_019_001, w_019_002, w_019_003, w_019_004, w_019_005, w_019_006, w_019_007, w_019_008, w_019_009, w_019_010, w_019_011, w_019_012, w_019_013, w_019_014, w_019_015, w_019_016, w_019_017, w_019_018, w_019_019, w_019_020;
  wire w_020_000, w_020_001, w_020_002, w_020_003, w_020_004, w_020_005, w_020_006, w_020_007, w_020_008, w_020_009, w_020_010, w_020_011, w_020_012, w_020_013, w_020_015, w_020_016, w_020_018, w_020_019, w_020_020, w_020_021, w_020_022, w_020_023, w_020_024, w_020_025, w_020_027, w_020_028, w_020_029, w_020_030, w_020_031, w_020_032, w_020_033, w_020_034, w_020_035, w_020_036, w_020_037, w_020_038, w_020_039, w_020_042, w_020_043, w_020_044, w_020_045, w_020_049, w_020_050, w_020_051, w_020_054, w_020_055, w_020_057, w_020_058, w_020_059, w_020_062, w_020_063, w_020_064, w_020_065, w_020_067, w_020_068, w_020_069, w_020_071, w_020_072, w_020_074, w_020_075, w_020_076, w_020_077, w_020_078, w_020_080, w_020_083, w_020_084, w_020_086, w_020_087, w_020_088, w_020_090, w_020_091, w_020_092, w_020_094, w_020_095, w_020_096, w_020_098, w_020_099, w_020_100, w_020_102, w_020_103, w_020_105, w_020_107, w_020_108, w_020_109, w_020_110, w_020_114, w_020_115, w_020_116, w_020_118, w_020_119, w_020_122, w_020_123, w_020_124, w_020_125, w_020_126, w_020_129, w_020_130, w_020_131, w_020_132, w_020_134, w_020_135, w_020_136, w_020_138, w_020_139, w_020_140, w_020_142, w_020_144, w_020_146, w_020_147, w_020_148, w_020_149, w_020_151, w_020_152, w_020_153, w_020_154, w_020_155, w_020_157, w_020_158, w_020_160, w_020_161, w_020_162, w_020_163, w_020_164, w_020_165, w_020_166, w_020_167, w_020_169, w_020_170, w_020_171, w_020_172, w_020_173, w_020_175, w_020_177, w_020_179, w_020_180, w_020_181, w_020_183, w_020_184, w_020_186, w_020_188, w_020_189, w_020_192, w_020_193, w_020_196, w_020_198, w_020_199, w_020_203, w_020_205, w_020_208, w_020_209, w_020_210, w_020_216, w_020_217, w_020_221, w_020_225, w_020_226, w_020_230, w_020_232, w_020_236, w_020_240, w_020_244, w_020_246, w_020_247, w_020_248, w_020_250, w_020_251, w_020_252, w_020_255, w_020_257, w_020_259, w_020_260, w_020_264, w_020_266, w_020_267, w_020_269, w_020_271, w_020_272, w_020_277, w_020_278, w_020_280, w_020_281, w_020_283, w_020_285, w_020_287, w_020_288, w_020_290, w_020_291, w_020_296, w_020_297, w_020_300, w_020_301, w_020_305, w_020_306, w_020_307, w_020_309, w_020_311, w_020_314, w_020_315, w_020_319, w_020_320, w_020_322, w_020_327, w_020_329, w_020_331, w_020_334, w_020_335, w_020_339, w_020_340, w_020_341, w_020_342, w_020_347, w_020_348, w_020_350, w_020_355, w_020_356, w_020_359, w_020_361, w_020_363, w_020_364, w_020_370, w_020_372, w_020_374, w_020_378, w_020_379, w_020_380, w_020_381, w_020_383, w_020_386, w_020_387, w_020_389, w_020_391, w_020_393, w_020_394, w_020_395, w_020_396, w_020_398, w_020_399, w_020_400, w_020_403, w_020_404, w_020_406, w_020_407, w_020_408, w_020_409, w_020_410, w_020_411, w_020_412, w_020_416, w_020_417, w_020_420, w_020_423, w_020_425, w_020_426, w_020_427, w_020_428, w_020_429, w_020_430, w_020_433, w_020_436, w_020_438, w_020_441, w_020_442, w_020_445, w_020_446, w_020_447, w_020_448, w_020_450, w_020_451, w_020_452, w_020_453, w_020_455, w_020_457, w_020_460, w_020_461, w_020_462, w_020_463, w_020_465, w_020_466, w_020_472, w_020_473, w_020_474, w_020_475, w_020_476, w_020_479, w_020_482, w_020_483, w_020_484, w_020_489, w_020_490, w_020_494, w_020_495, w_020_498, w_020_500, w_020_501, w_020_502, w_020_506, w_020_508, w_020_511, w_020_512, w_020_513, w_020_514, w_020_515, w_020_516, w_020_517, w_020_518, w_020_519, w_020_520, w_020_521, w_020_525, w_020_527, w_020_529, w_020_530, w_020_536, w_020_539, w_020_543, w_020_545, w_020_546, w_020_547, w_020_549, w_020_550, w_020_551, w_020_554, w_020_561, w_020_562, w_020_564, w_020_565, w_020_568, w_020_569, w_020_571, w_020_576, w_020_577, w_020_584, w_020_586, w_020_588, w_020_590, w_020_591, w_020_592, w_020_595, w_020_598, w_020_599, w_020_602, w_020_603, w_020_604, w_020_605, w_020_606, w_020_607, w_020_609, w_020_610, w_020_615, w_020_617, w_020_618, w_020_619, w_020_620, w_020_622, w_020_624, w_020_625, w_020_626, w_020_627, w_020_628, w_020_629, w_020_631;
  wire w_021_000, w_021_001, w_021_003, w_021_004, w_021_005, w_021_006, w_021_007, w_021_009, w_021_010, w_021_011, w_021_013, w_021_014, w_021_015, w_021_016, w_021_017, w_021_018, w_021_021, w_021_022, w_021_023, w_021_024, w_021_025, w_021_026, w_021_027, w_021_028, w_021_029, w_021_032, w_021_033, w_021_034, w_021_035, w_021_036, w_021_037, w_021_039, w_021_040, w_021_041, w_021_042, w_021_043, w_021_044, w_021_045, w_021_047, w_021_048, w_021_050, w_021_051, w_021_054, w_021_055, w_021_056, w_021_059, w_021_060, w_021_061, w_021_062, w_021_064, w_021_066, w_021_067, w_021_068, w_021_069, w_021_071, w_021_072, w_021_073, w_021_074, w_021_077, w_021_078, w_021_079, w_021_080, w_021_081, w_021_082, w_021_083, w_021_084, w_021_085, w_021_086, w_021_088, w_021_089, w_021_090, w_021_091, w_021_092, w_021_093, w_021_094, w_021_095, w_021_096, w_021_097, w_021_098, w_021_099, w_021_100, w_021_101, w_021_102, w_021_103, w_021_104, w_021_105, w_021_106, w_021_108, w_021_110, w_021_111, w_021_112, w_021_113, w_021_114, w_021_115, w_021_116, w_021_117, w_021_118, w_021_119, w_021_121, w_021_122, w_021_123, w_021_124, w_021_125, w_021_126, w_021_127, w_021_128, w_021_130, w_021_131, w_021_136, w_021_137, w_021_138, w_021_139, w_021_140, w_021_141, w_021_142, w_021_143, w_021_144, w_021_145, w_021_146, w_021_147, w_021_148, w_021_149, w_021_150, w_021_152, w_021_153, w_021_154, w_021_155, w_021_158, w_021_160, w_021_161, w_021_162, w_021_163, w_021_164, w_021_165, w_021_166, w_021_167, w_021_168, w_021_169, w_021_170, w_021_171, w_021_172, w_021_174, w_021_175, w_021_176, w_021_177, w_021_179, w_021_180, w_021_181, w_021_182, w_021_183, w_021_184, w_021_187, w_021_188, w_021_189, w_021_190, w_021_191, w_021_192, w_021_193, w_021_194, w_021_195, w_021_196, w_021_199, w_021_200, w_021_201, w_021_202, w_021_203, w_021_204, w_021_205, w_021_207, w_021_208, w_021_209, w_021_210, w_021_211, w_021_212, w_021_213, w_021_214, w_021_215, w_021_216, w_021_217, w_021_218, w_021_219, w_021_220, w_021_221, w_021_222, w_021_223, w_021_224, w_021_225, w_021_226, w_021_227, w_021_230, w_021_231, w_021_232, w_021_233, w_021_234, w_021_235, w_021_236, w_021_237, w_021_238, w_021_239, w_021_240, w_021_241, w_021_242, w_021_243, w_021_244, w_021_246, w_021_247, w_021_248, w_021_249, w_021_250, w_021_251, w_021_255, w_021_256, w_021_257, w_021_259, w_021_261, w_021_262, w_021_263, w_021_264, w_021_265, w_021_266, w_021_267, w_021_270, w_021_271, w_021_272, w_021_273, w_021_274;
  wire w_022_000, w_022_001, w_022_003, w_022_005, w_022_006, w_022_009, w_022_010, w_022_011, w_022_012, w_022_013, w_022_017, w_022_020, w_022_021, w_022_023, w_022_024, w_022_026, w_022_029, w_022_030, w_022_031, w_022_032, w_022_033, w_022_034, w_022_035, w_022_036, w_022_037, w_022_038, w_022_039, w_022_041, w_022_042, w_022_043, w_022_044, w_022_045, w_022_048, w_022_050, w_022_051, w_022_052, w_022_053, w_022_054, w_022_055, w_022_056, w_022_058, w_022_059, w_022_061, w_022_062, w_022_064, w_022_065, w_022_066, w_022_068, w_022_071, w_022_074, w_022_076, w_022_077, w_022_079, w_022_080, w_022_081, w_022_082, w_022_083, w_022_084, w_022_086, w_022_087, w_022_088, w_022_089, w_022_090, w_022_093, w_022_094, w_022_097, w_022_098, w_022_100, w_022_102, w_022_103, w_022_104, w_022_111, w_022_112, w_022_114, w_022_115, w_022_117, w_022_118, w_022_119, w_022_120, w_022_123, w_022_124, w_022_125, w_022_126, w_022_128, w_022_129, w_022_130, w_022_131, w_022_132, w_022_134, w_022_135, w_022_136, w_022_137, w_022_138, w_022_140, w_022_141, w_022_142, w_022_144, w_022_145, w_022_148, w_022_149, w_022_150, w_022_151, w_022_152, w_022_153, w_022_154, w_022_155, w_022_158, w_022_160, w_022_161, w_022_163, w_022_164, w_022_165, w_022_167, w_022_168, w_022_170, w_022_172, w_022_173, w_022_174, w_022_175, w_022_177, w_022_181, w_022_183, w_022_185, w_022_186, w_022_187, w_022_188, w_022_193, w_022_194, w_022_195, w_022_196, w_022_198, w_022_199, w_022_200, w_022_201, w_022_202, w_022_204, w_022_205, w_022_206, w_022_207, w_022_210, w_022_211, w_022_213, w_022_214, w_022_219, w_022_220, w_022_221, w_022_226, w_022_227, w_022_229, w_022_231, w_022_232, w_022_234, w_022_235, w_022_236, w_022_237, w_022_238, w_022_239, w_022_240, w_022_241, w_022_243, w_022_245, w_022_247, w_022_248, w_022_249, w_022_251, w_022_252, w_022_253, w_022_255, w_022_256, w_022_258, w_022_259, w_022_261, w_022_262, w_022_263, w_022_264, w_022_265, w_022_266, w_022_267, w_022_268, w_022_269, w_022_270, w_022_271, w_022_272, w_022_276, w_022_277, w_022_279, w_022_280, w_022_281, w_022_282, w_022_283, w_022_287, w_022_288, w_022_290, w_022_291, w_022_293, w_022_294, w_022_295, w_022_296, w_022_297, w_022_298, w_022_300, w_022_303, w_022_304, w_022_305, w_022_307, w_022_309, w_022_310, w_022_311, w_022_313, w_022_315, w_022_316, w_022_319, w_022_320, w_022_321, w_022_322, w_022_323, w_022_328, w_022_330, w_022_331, w_022_332, w_022_333, w_022_334, w_022_336, w_022_337, w_022_341, w_022_342, w_022_343, w_022_344, w_022_345, w_022_347, w_022_348, w_022_349, w_022_351, w_022_352, w_022_353, w_022_355, w_022_356, w_022_357, w_022_360, w_022_361, w_022_362, w_022_364, w_022_365, w_022_366, w_022_367, w_022_368, w_022_369, w_022_370, w_022_373, w_022_376, w_022_378, w_022_380, w_022_381, w_022_382, w_022_383, w_022_384, w_022_385, w_022_386, w_022_388, w_022_389, w_022_390, w_022_392, w_022_393, w_022_395, w_022_397, w_022_399, w_022_401, w_022_404, w_022_407, w_022_408;
  wire w_023_000, w_023_002, w_023_003, w_023_005, w_023_006, w_023_007, w_023_008, w_023_009, w_023_011, w_023_012, w_023_013, w_023_015, w_023_016, w_023_017, w_023_018, w_023_019, w_023_020, w_023_021, w_023_023, w_023_024, w_023_025, w_023_026, w_023_027, w_023_028, w_023_029, w_023_031, w_023_032, w_023_033, w_023_034, w_023_035, w_023_037, w_023_038, w_023_039, w_023_040, w_023_041, w_023_042, w_023_043, w_023_044, w_023_045, w_023_046, w_023_047, w_023_048, w_023_049, w_023_051, w_023_052, w_023_053, w_023_054, w_023_055, w_023_056, w_023_058, w_023_059, w_023_060, w_023_062, w_023_063, w_023_064, w_023_065, w_023_066, w_023_067, w_023_068, w_023_069, w_023_070, w_023_071, w_023_073, w_023_074, w_023_075, w_023_076, w_023_077, w_023_078, w_023_079, w_023_080, w_023_081, w_023_082, w_023_083, w_023_084, w_023_086, w_023_087, w_023_088, w_023_090, w_023_091, w_023_092, w_023_093, w_023_095, w_023_096, w_023_098, w_023_099, w_023_100, w_023_101, w_023_102, w_023_103, w_023_104, w_023_105, w_023_106, w_023_107, w_023_108, w_023_109, w_023_110, w_023_111, w_023_112, w_023_113, w_023_114, w_023_115, w_023_116, w_023_117, w_023_120, w_023_121, w_023_122, w_023_123, w_023_124, w_023_125, w_023_128, w_023_129, w_023_130, w_023_131, w_023_132, w_023_134, w_023_135, w_023_136, w_023_137, w_023_138, w_023_139, w_023_141, w_023_142, w_023_143, w_023_144, w_023_145, w_023_146, w_023_147, w_023_148, w_023_149, w_023_150, w_023_151, w_023_152, w_023_153, w_023_154, w_023_155, w_023_156, w_023_157, w_023_158, w_023_159, w_023_160, w_023_161, w_023_162, w_023_164, w_023_165, w_023_166, w_023_169, w_023_170, w_023_171, w_023_172, w_023_173, w_023_175, w_023_176, w_023_178, w_023_179, w_023_181, w_023_183, w_023_184, w_023_186, w_023_188, w_023_189, w_023_191, w_023_192, w_023_193, w_023_194, w_023_195, w_023_196, w_023_197, w_023_198, w_023_199, w_023_200, w_023_201, w_023_202, w_023_203, w_023_205, w_023_206, w_023_207, w_023_208, w_023_210, w_023_212, w_023_213, w_023_214, w_023_215, w_023_216, w_023_217;
  wire w_024_000, w_024_003, w_024_004, w_024_005, w_024_007, w_024_008, w_024_009, w_024_010, w_024_013, w_024_015, w_024_016, w_024_017, w_024_018, w_024_020, w_024_022, w_024_024, w_024_025, w_024_026, w_024_027, w_024_028, w_024_029, w_024_030, w_024_032, w_024_034, w_024_035, w_024_036, w_024_039, w_024_040, w_024_041, w_024_042, w_024_044, w_024_045, w_024_048, w_024_049, w_024_051, w_024_054, w_024_055, w_024_056, w_024_057, w_024_059, w_024_060, w_024_061, w_024_062, w_024_064, w_024_065, w_024_068, w_024_070, w_024_071, w_024_073, w_024_077, w_024_079, w_024_081, w_024_082, w_024_083, w_024_086, w_024_088, w_024_089, w_024_090, w_024_092, w_024_093, w_024_095, w_024_096, w_024_097, w_024_098, w_024_099, w_024_101, w_024_102, w_024_103, w_024_105, w_024_107, w_024_108, w_024_109, w_024_110, w_024_115, w_024_116, w_024_117, w_024_118, w_024_119, w_024_120, w_024_121, w_024_122, w_024_123, w_024_125, w_024_126, w_024_127, w_024_128, w_024_129, w_024_130, w_024_133, w_024_137, w_024_139, w_024_141, w_024_142, w_024_143, w_024_144, w_024_145, w_024_146, w_024_151, w_024_155, w_024_157, w_024_164, w_024_166, w_024_171, w_024_172, w_024_173, w_024_175, w_024_176, w_024_178, w_024_180, w_024_181, w_024_182, w_024_183, w_024_184, w_024_186, w_024_187, w_024_188, w_024_189, w_024_190, w_024_191, w_024_192, w_024_193, w_024_194, w_024_195, w_024_197, w_024_200, w_024_202, w_024_205, w_024_206, w_024_207, w_024_208, w_024_209, w_024_210, w_024_211, w_024_212, w_024_213, w_024_214, w_024_215, w_024_216, w_024_218, w_024_219, w_024_221, w_024_222, w_024_223, w_024_224, w_024_225, w_024_227, w_024_229, w_024_230, w_024_231, w_024_243, w_024_244, w_024_247, w_024_253, w_024_254, w_024_257, w_024_258, w_024_260, w_024_262, w_024_263, w_024_265, w_024_268, w_024_272, w_024_273, w_024_275, w_024_276, w_024_277, w_024_280, w_024_283, w_024_284, w_024_286, w_024_292, w_024_295, w_024_299, w_024_300, w_024_301, w_024_305, w_024_307, w_024_311, w_024_312, w_024_313, w_024_316, w_024_317, w_024_319, w_024_324, w_024_326, w_024_327, w_024_329, w_024_339, w_024_342, w_024_346, w_024_347, w_024_354, w_024_355, w_024_358, w_024_359, w_024_361, w_024_365, w_024_367, w_024_369, w_024_371, w_024_372, w_024_373, w_024_377, w_024_378, w_024_386, w_024_387, w_024_388, w_024_389, w_024_391, w_024_392, w_024_395, w_024_399, w_024_401, w_024_404, w_024_411, w_024_413, w_024_418, w_024_419, w_024_421, w_024_422, w_024_424, w_024_426, w_024_430, w_024_433, w_024_434, w_024_435, w_024_436, w_024_439, w_024_441, w_024_444, w_024_445, w_024_447, w_024_452, w_024_456, w_024_457, w_024_461, w_024_464, w_024_473, w_024_477, w_024_478, w_024_481, w_024_482, w_024_483, w_024_489, w_024_491, w_024_492, w_024_493, w_024_496, w_024_499, w_024_503, w_024_506, w_024_507, w_024_509, w_024_510, w_024_513, w_024_516, w_024_517, w_024_518, w_024_521, w_024_523, w_024_524, w_024_525, w_024_528, w_024_530, w_024_534, w_024_535, w_024_537, w_024_541, w_024_542, w_024_545, w_024_549, w_024_551, w_024_557, w_024_558, w_024_559, w_024_563, w_024_565, w_024_566, w_024_569, w_024_571, w_024_574, w_024_577, w_024_579, w_024_581, w_024_582, w_024_583, w_024_584, w_024_585, w_024_586, w_024_587, w_024_589, w_024_591, w_024_592, w_024_593, w_024_594, w_024_595, w_024_596, w_024_597, w_024_599;
  wire w_025_000, w_025_001, w_025_002, w_025_003, w_025_004, w_025_005, w_025_006, w_025_007, w_025_008, w_025_009, w_025_010, w_025_011, w_025_012, w_025_013, w_025_015, w_025_016, w_025_018, w_025_019, w_025_021, w_025_023, w_025_024, w_025_025, w_025_026, w_025_027, w_025_028, w_025_029, w_025_032, w_025_034, w_025_035, w_025_036, w_025_037, w_025_038, w_025_039, w_025_040, w_025_042, w_025_043, w_025_044, w_025_048, w_025_049, w_025_050, w_025_051, w_025_053, w_025_054, w_025_055, w_025_056, w_025_057, w_025_059, w_025_060, w_025_061, w_025_062, w_025_063, w_025_064, w_025_066, w_025_067, w_025_069, w_025_072, w_025_073, w_025_074, w_025_075, w_025_076, w_025_077, w_025_078, w_025_079, w_025_080, w_025_081, w_025_082, w_025_083, w_025_084, w_025_086, w_025_088, w_025_089, w_025_092, w_025_093, w_025_094, w_025_095, w_025_096, w_025_097, w_025_098, w_025_099, w_025_100, w_025_101, w_025_102, w_025_103, w_025_104, w_025_105, w_025_106, w_025_108, w_025_110, w_025_111, w_025_112, w_025_113, w_025_114, w_025_115, w_025_116, w_025_117, w_025_118, w_025_119, w_025_120, w_025_121, w_025_122, w_025_123, w_025_124, w_025_125, w_025_126, w_025_127, w_025_130, w_025_131, w_025_132, w_025_133, w_025_134, w_025_135, w_025_137, w_025_138, w_025_139, w_025_140, w_025_141, w_025_142, w_025_143, w_025_145, w_025_147, w_025_148, w_025_149, w_025_151, w_025_152, w_025_154, w_025_155, w_025_157, w_025_158, w_025_160, w_025_161, w_025_162, w_025_163, w_025_164, w_025_165, w_025_166, w_025_167, w_025_168, w_025_169, w_025_170, w_025_171, w_025_172, w_025_173, w_025_174, w_025_176, w_025_177, w_025_178, w_025_179, w_025_180, w_025_181, w_025_182, w_025_184, w_025_186, w_025_187, w_025_188, w_025_189, w_025_191, w_025_192, w_025_194, w_025_199, w_025_201, w_025_202, w_025_204, w_025_205, w_025_207, w_025_209, w_025_210, w_025_211, w_025_216, w_025_217, w_025_218, w_025_219, w_025_221, w_025_222, w_025_223, w_025_227, w_025_228, w_025_229, w_025_231, w_025_233, w_025_234, w_025_235, w_025_236, w_025_239, w_025_240, w_025_241, w_025_242, w_025_243, w_025_247, w_025_249, w_025_251, w_025_253, w_025_257, w_025_258, w_025_261, w_025_263, w_025_264, w_025_265, w_025_269, w_025_271, w_025_272, w_025_277, w_025_279, w_025_280, w_025_281, w_025_282, w_025_283, w_025_287, w_025_288, w_025_290, w_025_291, w_025_294, w_025_296, w_025_297, w_025_303, w_025_304, w_025_305, w_025_306, w_025_307, w_025_308;
  wire w_026_000, w_026_002, w_026_004, w_026_005, w_026_006, w_026_007, w_026_008, w_026_009, w_026_010, w_026_012, w_026_013, w_026_015, w_026_018, w_026_023, w_026_025, w_026_026, w_026_027, w_026_028, w_026_033, w_026_038, w_026_039, w_026_042, w_026_044, w_026_045, w_026_048, w_026_049, w_026_050, w_026_051, w_026_055, w_026_056, w_026_058, w_026_059, w_026_060, w_026_061, w_026_064, w_026_067, w_026_068, w_026_070, w_026_071, w_026_072, w_026_074, w_026_076, w_026_077, w_026_082, w_026_088, w_026_090, w_026_092, w_026_093, w_026_098, w_026_105, w_026_107, w_026_109, w_026_110, w_026_112, w_026_113, w_026_114, w_026_115, w_026_117, w_026_118, w_026_121, w_026_122, w_026_123, w_026_125, w_026_126, w_026_127, w_026_128, w_026_130, w_026_132, w_026_136, w_026_139, w_026_140, w_026_144, w_026_145, w_026_146, w_026_149, w_026_152, w_026_154, w_026_160, w_026_161, w_026_163, w_026_169, w_026_172, w_026_173, w_026_174, w_026_178, w_026_179, w_026_181, w_026_182, w_026_184, w_026_187, w_026_188, w_026_189, w_026_191, w_026_192, w_026_193, w_026_196, w_026_198, w_026_201, w_026_211, w_026_216, w_026_217, w_026_223, w_026_224, w_026_225, w_026_226, w_026_227, w_026_229, w_026_231, w_026_234, w_026_237, w_026_238, w_026_239, w_026_250, w_026_257, w_026_261, w_026_267, w_026_268, w_026_273, w_026_274, w_026_275, w_026_283, w_026_286, w_026_287, w_026_288, w_026_289, w_026_290, w_026_291, w_026_294, w_026_295, w_026_296, w_026_297, w_026_298, w_026_299, w_026_304, w_026_305, w_026_310, w_026_311, w_026_315, w_026_317, w_026_321, w_026_322, w_026_326, w_026_328, w_026_331, w_026_332, w_026_333, w_026_343, w_026_344, w_026_346, w_026_348, w_026_351, w_026_354, w_026_357, w_026_358, w_026_361, w_026_364, w_026_366, w_026_371, w_026_380, w_026_381, w_026_382, w_026_383, w_026_393, w_026_394, w_026_395, w_026_396, w_026_400, w_026_404, w_026_410, w_026_411, w_026_413, w_026_415, w_026_420, w_026_424, w_026_427, w_026_430, w_026_431, w_026_433, w_026_439, w_026_441, w_026_442, w_026_447, w_026_448, w_026_449, w_026_451, w_026_453, w_026_455, w_026_457, w_026_459, w_026_466, w_026_471, w_026_477, w_026_480, w_026_483, w_026_488, w_026_489, w_026_490, w_026_491, w_026_493, w_026_494, w_026_499, w_026_500, w_026_502, w_026_506, w_026_507, w_026_508, w_026_513, w_026_514, w_026_515, w_026_517, w_026_519, w_026_520, w_026_523, w_026_527, w_026_530, w_026_531, w_026_532, w_026_534, w_026_535, w_026_536, w_026_538, w_026_539, w_026_541, w_026_544, w_026_548, w_026_549, w_026_550, w_026_551, w_026_555, w_026_561, w_026_564, w_026_566, w_026_570, w_026_572, w_026_579, w_026_580, w_026_585, w_026_591, w_026_593, w_026_595, w_026_597, w_026_598, w_026_600, w_026_604, w_026_605, w_026_606, w_026_608, w_026_613, w_026_614, w_026_617, w_026_620, w_026_621, w_026_630, w_026_632, w_026_635, w_026_642, w_026_643, w_026_645, w_026_648, w_026_649, w_026_655, w_026_657, w_026_660, w_026_661, w_026_662, w_026_663, w_026_665, w_026_668, w_026_669, w_026_670, w_026_675, w_026_681, w_026_683, w_026_684, w_026_687, w_026_692, w_026_693, w_026_694, w_026_695, w_026_698, w_026_699, w_026_701, w_026_702, w_026_703, w_026_705, w_026_706, w_026_708, w_026_709, w_026_711, w_026_712, w_026_718, w_026_720;
  wire w_027_000, w_027_001, w_027_002, w_027_004, w_027_006, w_027_007, w_027_008, w_027_009, w_027_011, w_027_012, w_027_014, w_027_015, w_027_016, w_027_018, w_027_019, w_027_020, w_027_023, w_027_024, w_027_026, w_027_027, w_027_028, w_027_030, w_027_031, w_027_032, w_027_033, w_027_034, w_027_035, w_027_036, w_027_037, w_027_039, w_027_040, w_027_041, w_027_042, w_027_043, w_027_044, w_027_045, w_027_046, w_027_047, w_027_048, w_027_049, w_027_050, w_027_051, w_027_053, w_027_054, w_027_055, w_027_056, w_027_057, w_027_058, w_027_059, w_027_060, w_027_061, w_027_062, w_027_063, w_027_064, w_027_065, w_027_066, w_027_067, w_027_068, w_027_070, w_027_071, w_027_072, w_027_073, w_027_074, w_027_075, w_027_076, w_027_077, w_027_078, w_027_079, w_027_080, w_027_081, w_027_082, w_027_083, w_027_084, w_027_086, w_027_088, w_027_089, w_027_090, w_027_091, w_027_092, w_027_093, w_027_094, w_027_095, w_027_096, w_027_097, w_027_098, w_027_099, w_027_101, w_027_102, w_027_103, w_027_104, w_027_105, w_027_107, w_027_109, w_027_110, w_027_111, w_027_112, w_027_113, w_027_114, w_027_115, w_027_116, w_027_117, w_027_118, w_027_119, w_027_120, w_027_121, w_027_122, w_027_123, w_027_124, w_027_125, w_027_126, w_027_127, w_027_129, w_027_130, w_027_131, w_027_132, w_027_134, w_027_135, w_027_136, w_027_138, w_027_139, w_027_140, w_027_141, w_027_142, w_027_143, w_027_145, w_027_146, w_027_148, w_027_149, w_027_150, w_027_151, w_027_153, w_027_155, w_027_156, w_027_157, w_027_158, w_027_159, w_027_160, w_027_161, w_027_162, w_027_163, w_027_164, w_027_165, w_027_166, w_027_167, w_027_168, w_027_169, w_027_170, w_027_171, w_027_173, w_027_175, w_027_176, w_027_177, w_027_178, w_027_179, w_027_180, w_027_181, w_027_182, w_027_183, w_027_184, w_027_185, w_027_187, w_027_188, w_027_189, w_027_191, w_027_192, w_027_194, w_027_195, w_027_197, w_027_198, w_027_199, w_027_202, w_027_204;
  wire w_028_000, w_028_001, w_028_003, w_028_005, w_028_006, w_028_008, w_028_011, w_028_012, w_028_013, w_028_014, w_028_018, w_028_021, w_028_022, w_028_025, w_028_026, w_028_027, w_028_028, w_028_029, w_028_030, w_028_033, w_028_034, w_028_035, w_028_036, w_028_037, w_028_038, w_028_039, w_028_040, w_028_041, w_028_042, w_028_044, w_028_045, w_028_050, w_028_052, w_028_053, w_028_056, w_028_057, w_028_058, w_028_060, w_028_064, w_028_065, w_028_068, w_028_069, w_028_070, w_028_072, w_028_074, w_028_076, w_028_077, w_028_078, w_028_079, w_028_080, w_028_084, w_028_085, w_028_086, w_028_087, w_028_088, w_028_089, w_028_090, w_028_091, w_028_094, w_028_096, w_028_097, w_028_098, w_028_099, w_028_101, w_028_102, w_028_104, w_028_105, w_028_106, w_028_107, w_028_109, w_028_110, w_028_111, w_028_113, w_028_115, w_028_117, w_028_118, w_028_119, w_028_120, w_028_121, w_028_122, w_028_123, w_028_125, w_028_126, w_028_127, w_028_128, w_028_129, w_028_130, w_028_131, w_028_132, w_028_133, w_028_134, w_028_135, w_028_136, w_028_137, w_028_139, w_028_140, w_028_141, w_028_142, w_028_143, w_028_144, w_028_145, w_028_147, w_028_149, w_028_150, w_028_151, w_028_152, w_028_154, w_028_156, w_028_160, w_028_162, w_028_163, w_028_165, w_028_170, w_028_171, w_028_173, w_028_175, w_028_177, w_028_178, w_028_181, w_028_182, w_028_183, w_028_184, w_028_185, w_028_186, w_028_187, w_028_190, w_028_191, w_028_196, w_028_197, w_028_198, w_028_200, w_028_201, w_028_202, w_028_203, w_028_204, w_028_205, w_028_206, w_028_208, w_028_209, w_028_215, w_028_216, w_028_222, w_028_224, w_028_226, w_028_228, w_028_231, w_028_232, w_028_234, w_028_240, w_028_244, w_028_245, w_028_248, w_028_251, w_028_252, w_028_254, w_028_255, w_028_256, w_028_258, w_028_260, w_028_262, w_028_263, w_028_264, w_028_267, w_028_268, w_028_270, w_028_274, w_028_275, w_028_277, w_028_279, w_028_283, w_028_284, w_028_287, w_028_296, w_028_299, w_028_300, w_028_301, w_028_302, w_028_304, w_028_310, w_028_313, w_028_317, w_028_321, w_028_324, w_028_325, w_028_326, w_028_335, w_028_336, w_028_340, w_028_345, w_028_350, w_028_354, w_028_361, w_028_362, w_028_366, w_028_368, w_028_374, w_028_376, w_028_380, w_028_390, w_028_392, w_028_393, w_028_397, w_028_400, w_028_402, w_028_405, w_028_408, w_028_409, w_028_411, w_028_413, w_028_415, w_028_416, w_028_425, w_028_427, w_028_433, w_028_436, w_028_437, w_028_438, w_028_440, w_028_441, w_028_446, w_028_449, w_028_456, w_028_458, w_028_462, w_028_463, w_028_464, w_028_465, w_028_470, w_028_473, w_028_474, w_028_475, w_028_479, w_028_483, w_028_488, w_028_489, w_028_490, w_028_491, w_028_497, w_028_499, w_028_503, w_028_505, w_028_512, w_028_517, w_028_521, w_028_522, w_028_523, w_028_526, w_028_527, w_028_528, w_028_536, w_028_541, w_028_542, w_028_543, w_028_547, w_028_550, w_028_551, w_028_554, w_028_559, w_028_560, w_028_564, w_028_565, w_028_567, w_028_569, w_028_574, w_028_575, w_028_578, w_028_586, w_028_588, w_028_589, w_028_590, w_028_591, w_028_592, w_028_593, w_028_594, w_028_595, w_028_596, w_028_597, w_028_599, w_028_601, w_028_602, w_028_603, w_028_604, w_028_605, w_028_607;
  wire w_029_000, w_029_001, w_029_002, w_029_003, w_029_004, w_029_005, w_029_006, w_029_007, w_029_008, w_029_009, w_029_010, w_029_011, w_029_012, w_029_013, w_029_014, w_029_015, w_029_016, w_029_017, w_029_018, w_029_019, w_029_020, w_029_021, w_029_022, w_029_023, w_029_024, w_029_025, w_029_026, w_029_027, w_029_028, w_029_029, w_029_031, w_029_032, w_029_033, w_029_035, w_029_036, w_029_037, w_029_038, w_029_039, w_029_041, w_029_042, w_029_043, w_029_044, w_029_045, w_029_046, w_029_047, w_029_048, w_029_049, w_029_050, w_029_051, w_029_052, w_029_053, w_029_054, w_029_055, w_029_056, w_029_057, w_029_058, w_029_059, w_029_060, w_029_061, w_029_062, w_029_063, w_029_064, w_029_065, w_029_066, w_029_067, w_029_068, w_029_069, w_029_070, w_029_071, w_029_072, w_029_073, w_029_074, w_029_075, w_029_076, w_029_077, w_029_078, w_029_079, w_029_080, w_029_081, w_029_082, w_029_083, w_029_085, w_029_086, w_029_087, w_029_088, w_029_089, w_029_090, w_029_091, w_029_092, w_029_093, w_029_094, w_029_095, w_029_096, w_029_097, w_029_098, w_029_099, w_029_100, w_029_101, w_029_102, w_029_103, w_029_104, w_029_105, w_029_106, w_029_107, w_029_108, w_029_109, w_029_110, w_029_111, w_029_112, w_029_113, w_029_114, w_029_115, w_029_116, w_029_117;
  wire w_030_004, w_030_006, w_030_007, w_030_008, w_030_009, w_030_011, w_030_012, w_030_013, w_030_015, w_030_016, w_030_017, w_030_020, w_030_021, w_030_022, w_030_024, w_030_031, w_030_033, w_030_035, w_030_036, w_030_037, w_030_040, w_030_041, w_030_044, w_030_047, w_030_048, w_030_049, w_030_050, w_030_051, w_030_052, w_030_053, w_030_055, w_030_056, w_030_057, w_030_061, w_030_064, w_030_067, w_030_069, w_030_070, w_030_071, w_030_073, w_030_074, w_030_076, w_030_077, w_030_078, w_030_080, w_030_083, w_030_086, w_030_088, w_030_089, w_030_090, w_030_091, w_030_097, w_030_099, w_030_100, w_030_101, w_030_102, w_030_104, w_030_105, w_030_106, w_030_107, w_030_108, w_030_112, w_030_113, w_030_117, w_030_119, w_030_121, w_030_123, w_030_125, w_030_132, w_030_134, w_030_136, w_030_137, w_030_138, w_030_143, w_030_144, w_030_145, w_030_146, w_030_148, w_030_149, w_030_151, w_030_152, w_030_155, w_030_157, w_030_159, w_030_161, w_030_162, w_030_163, w_030_167, w_030_168, w_030_171, w_030_172, w_030_174, w_030_177, w_030_178, w_030_179, w_030_180, w_030_183, w_030_184, w_030_185, w_030_188, w_030_191, w_030_192, w_030_194, w_030_196, w_030_198, w_030_199, w_030_200, w_030_201, w_030_202, w_030_203, w_030_204, w_030_205, w_030_207, w_030_208, w_030_210, w_030_212, w_030_213, w_030_214, w_030_215, w_030_219, w_030_220, w_030_222, w_030_223, w_030_224, w_030_225, w_030_226, w_030_227, w_030_228, w_030_229, w_030_231, w_030_235, w_030_236, w_030_239, w_030_240, w_030_241, w_030_242, w_030_243, w_030_244, w_030_247, w_030_248, w_030_249, w_030_250, w_030_251, w_030_252, w_030_257, w_030_258, w_030_259, w_030_261, w_030_262, w_030_263, w_030_264, w_030_265, w_030_267, w_030_268, w_030_269, w_030_270, w_030_273, w_030_274, w_030_275, w_030_276, w_030_278, w_030_279, w_030_280, w_030_284, w_030_287, w_030_288, w_030_290, w_030_291, w_030_292, w_030_293, w_030_295, w_030_296, w_030_298, w_030_300, w_030_301, w_030_302, w_030_305, w_030_307, w_030_308, w_030_309, w_030_311, w_030_312, w_030_313, w_030_315, w_030_316, w_030_317, w_030_318, w_030_319, w_030_320, w_030_324, w_030_325, w_030_326, w_030_327, w_030_328, w_030_330, w_030_331, w_030_332, w_030_337, w_030_338, w_030_339, w_030_340, w_030_341, w_030_345, w_030_346, w_030_348, w_030_349, w_030_350, w_030_352, w_030_353, w_030_354, w_030_355, w_030_358, w_030_359, w_030_360, w_030_364, w_030_365, w_030_367, w_030_369, w_030_370, w_030_372, w_030_374, w_030_375, w_030_377, w_030_378, w_030_379, w_030_382, w_030_385, w_030_391, w_030_392, w_030_393, w_030_396, w_030_399, w_030_408, w_030_409, w_030_410, w_030_411, w_030_413, w_030_414, w_030_417, w_030_419;
  wire w_031_001, w_031_002, w_031_008, w_031_009, w_031_011, w_031_012, w_031_014, w_031_015, w_031_016, w_031_017, w_031_020, w_031_021, w_031_026, w_031_027, w_031_030, w_031_032, w_031_033, w_031_034, w_031_040, w_031_043, w_031_049, w_031_050, w_031_054, w_031_055, w_031_058, w_031_059, w_031_065, w_031_066, w_031_068, w_031_069, w_031_070, w_031_072, w_031_074, w_031_076, w_031_081, w_031_082, w_031_083, w_031_086, w_031_088, w_031_090, w_031_092, w_031_093, w_031_095, w_031_097, w_031_100, w_031_101, w_031_102, w_031_103, w_031_105, w_031_107, w_031_111, w_031_112, w_031_116, w_031_118, w_031_119, w_031_120, w_031_121, w_031_122, w_031_124, w_031_125, w_031_126, w_031_127, w_031_128, w_031_129, w_031_130, w_031_131, w_031_133, w_031_134, w_031_136, w_031_138, w_031_143, w_031_144, w_031_145, w_031_147, w_031_148, w_031_150, w_031_151, w_031_153, w_031_154, w_031_155, w_031_156, w_031_160, w_031_161, w_031_162, w_031_163, w_031_165, w_031_168, w_031_171, w_031_174, w_031_175, w_031_176, w_031_177, w_031_178, w_031_179, w_031_182, w_031_186, w_031_188, w_031_193, w_031_195, w_031_202, w_031_204, w_031_205, w_031_206, w_031_213, w_031_214, w_031_218, w_031_223, w_031_231, w_031_234, w_031_235, w_031_236, w_031_239, w_031_251, w_031_253, w_031_256, w_031_259, w_031_260, w_031_265, w_031_268, w_031_271, w_031_272, w_031_273, w_031_276, w_031_277, w_031_281, w_031_287, w_031_290, w_031_295, w_031_297, w_031_302, w_031_308, w_031_309, w_031_315, w_031_319, w_031_330, w_031_336, w_031_340, w_031_343, w_031_346, w_031_356, w_031_362, w_031_366, w_031_367, w_031_370, w_031_375, w_031_377, w_031_380, w_031_382, w_031_386, w_031_387, w_031_389, w_031_390, w_031_392, w_031_410, w_031_413, w_031_415, w_031_417, w_031_419, w_031_420, w_031_422, w_031_423, w_031_425, w_031_434, w_031_437, w_031_439, w_031_440, w_031_442, w_031_444, w_031_445, w_031_446, w_031_453, w_031_456, w_031_457, w_031_460, w_031_462, w_031_463, w_031_465, w_031_466, w_031_467, w_031_469, w_031_470, w_031_471, w_031_472, w_031_476, w_031_482, w_031_483, w_031_487, w_031_488, w_031_489, w_031_490, w_031_494, w_031_495, w_031_497, w_031_498, w_031_499, w_031_501, w_031_508, w_031_509, w_031_511, w_031_514, w_031_518, w_031_520, w_031_528, w_031_531, w_031_539, w_031_540, w_031_541, w_031_543, w_031_546, w_031_548, w_031_553, w_031_555, w_031_556, w_031_557, w_031_558, w_031_561, w_031_566, w_031_570, w_031_571, w_031_574, w_031_581, w_031_582, w_031_588, w_031_590, w_031_593, w_031_595, w_031_596, w_031_599, w_031_601, w_031_602, w_031_604, w_031_605, w_031_610, w_031_611, w_031_612, w_031_613, w_031_614, w_031_615, w_031_616, w_031_618, w_031_620, w_031_621, w_031_622, w_031_623, w_031_624, w_031_625, w_031_626, w_031_627, w_031_628, w_031_629, w_031_631;
  wire w_032_000, w_032_011, w_032_013, w_032_019, w_032_021, w_032_022, w_032_025, w_032_028, w_032_030, w_032_031, w_032_033, w_032_037, w_032_039, w_032_041, w_032_042, w_032_043, w_032_044, w_032_045, w_032_046, w_032_049, w_032_051, w_032_052, w_032_053, w_032_057, w_032_060, w_032_064, w_032_065, w_032_066, w_032_067, w_032_068, w_032_072, w_032_073, w_032_074, w_032_076, w_032_077, w_032_078, w_032_083, w_032_084, w_032_085, w_032_086, w_032_088, w_032_089, w_032_090, w_032_091, w_032_092, w_032_095, w_032_097, w_032_098, w_032_099, w_032_102, w_032_103, w_032_105, w_032_106, w_032_108, w_032_109, w_032_110, w_032_114, w_032_115, w_032_116, w_032_118, w_032_120, w_032_121, w_032_122, w_032_123, w_032_124, w_032_129, w_032_132, w_032_133, w_032_134, w_032_136, w_032_137, w_032_138, w_032_143, w_032_144, w_032_148, w_032_149, w_032_150, w_032_151, w_032_152, w_032_153, w_032_154, w_032_158, w_032_160, w_032_163, w_032_165, w_032_167, w_032_168, w_032_169, w_032_172, w_032_173, w_032_174, w_032_175, w_032_177, w_032_178, w_032_180, w_032_183, w_032_184, w_032_185, w_032_186, w_032_187, w_032_189, w_032_191, w_032_192, w_032_193, w_032_194, w_032_195, w_032_197, w_032_204, w_032_207, w_032_208, w_032_209, w_032_210, w_032_211, w_032_213, w_032_219, w_032_221, w_032_225, w_032_226, w_032_228, w_032_229, w_032_232, w_032_234, w_032_239, w_032_240, w_032_243, w_032_247, w_032_249, w_032_254, w_032_257, w_032_259, w_032_261, w_032_264, w_032_269, w_032_273, w_032_275, w_032_279, w_032_280, w_032_281, w_032_283, w_032_285, w_032_287, w_032_290, w_032_293, w_032_294, w_032_295, w_032_297, w_032_298, w_032_300, w_032_307, w_032_309, w_032_310, w_032_312, w_032_313, w_032_321, w_032_322, w_032_325, w_032_328, w_032_330, w_032_331, w_032_342, w_032_345, w_032_346, w_032_348, w_032_350, w_032_352, w_032_355, w_032_357, w_032_359, w_032_360, w_032_363, w_032_364, w_032_368, w_032_376, w_032_377, w_032_379, w_032_389, w_032_391, w_032_395, w_032_398, w_032_399, w_032_404, w_032_409, w_032_410, w_032_411, w_032_414, w_032_418, w_032_425, w_032_429, w_032_430, w_032_433, w_032_434, w_032_437, w_032_438, w_032_442, w_032_443, w_032_444, w_032_445, w_032_446, w_032_448, w_032_449, w_032_451, w_032_457, w_032_462, w_032_464, w_032_465, w_032_466, w_032_471, w_032_477, w_032_478, w_032_490, w_032_491, w_032_493, w_032_496, w_032_497, w_032_499, w_032_502, w_032_504, w_032_507, w_032_508, w_032_509, w_032_510, w_032_512, w_032_514, w_032_515, w_032_520, w_032_521, w_032_524, w_032_525, w_032_526, w_032_533, w_032_537, w_032_540, w_032_541, w_032_545, w_032_546, w_032_552, w_032_553, w_032_559, w_032_562, w_032_568, w_032_569, w_032_570, w_032_574, w_032_575, w_032_579, w_032_583, w_032_588, w_032_594, w_032_596, w_032_597, w_032_599, w_032_603, w_032_604, w_032_605, w_032_606, w_032_607, w_032_609;
  wire w_033_001, w_033_002, w_033_008, w_033_009, w_033_011, w_033_012, w_033_014, w_033_015, w_033_016, w_033_017, w_033_019, w_033_021, w_033_022, w_033_024, w_033_026, w_033_029, w_033_053, w_033_057, w_033_059, w_033_061, w_033_062, w_033_065, w_033_068, w_033_076, w_033_082, w_033_084, w_033_085, w_033_086, w_033_087, w_033_091, w_033_094, w_033_095, w_033_100, w_033_109, w_033_111, w_033_114, w_033_116, w_033_119, w_033_121, w_033_123, w_033_127, w_033_129, w_033_132, w_033_142, w_033_143, w_033_148, w_033_149, w_033_157, w_033_159, w_033_160, w_033_161, w_033_162, w_033_163, w_033_171, w_033_172, w_033_181, w_033_182, w_033_183, w_033_184, w_033_191, w_033_194, w_033_197, w_033_200, w_033_201, w_033_207, w_033_208, w_033_209, w_033_216, w_033_217, w_033_220, w_033_224, w_033_231, w_033_235, w_033_236, w_033_238, w_033_241, w_033_244, w_033_249, w_033_250, w_033_251, w_033_253, w_033_256, w_033_259, w_033_263, w_033_269, w_033_272, w_033_275, w_033_278, w_033_282, w_033_289, w_033_291, w_033_293, w_033_297, w_033_309, w_033_310, w_033_312, w_033_313, w_033_318, w_033_319, w_033_321, w_033_322, w_033_323, w_033_328, w_033_329, w_033_330, w_033_331, w_033_335, w_033_336, w_033_339, w_033_340, w_033_341, w_033_354, w_033_355, w_033_358, w_033_363, w_033_365, w_033_366, w_033_369, w_033_372, w_033_377, w_033_378, w_033_379, w_033_380, w_033_382, w_033_391, w_033_392, w_033_396, w_033_404, w_033_406, w_033_407, w_033_414, w_033_419, w_033_426, w_033_427, w_033_428, w_033_436, w_033_437, w_033_442, w_033_447, w_033_449, w_033_451, w_033_452, w_033_453, w_033_462, w_033_468, w_033_475, w_033_486, w_033_487, w_033_488, w_033_492, w_033_493, w_033_494, w_033_505, w_033_506, w_033_509, w_033_510, w_033_511, w_033_512, w_033_513, w_033_515, w_033_516, w_033_517, w_033_522, w_033_530, w_033_534, w_033_535, w_033_537, w_033_539, w_033_541, w_033_545, w_033_546, w_033_551, w_033_555, w_033_557, w_033_558, w_033_560, w_033_566, w_033_568, w_033_569, w_033_574, w_033_580, w_033_583, w_033_587, w_033_590, w_033_604, w_033_605, w_033_608, w_033_613, w_033_614, w_033_617, w_033_618, w_033_619, w_033_622, w_033_629, w_033_630, w_033_631, w_033_637, w_033_638, w_033_639, w_033_646, w_033_647, w_033_653, w_033_656, w_033_658, w_033_660, w_033_670, w_033_671, w_033_675, w_033_685, w_033_689, w_033_692, w_033_695, w_033_698, w_033_703, w_033_705, w_033_710, w_033_711, w_033_715, w_033_718, w_033_719, w_033_722, w_033_724, w_033_725, w_033_726, w_033_727, w_033_730, w_033_735, w_033_740, w_033_745, w_033_748, w_033_751, w_033_753, w_033_756, w_033_762, w_033_766, w_033_769, w_033_770, w_033_771, w_033_775, w_033_779, w_033_783;
  wire w_034_000, w_034_001, w_034_002, w_034_003, w_034_004, w_034_005, w_034_006, w_034_007, w_034_008, w_034_009, w_034_010, w_034_011, w_034_012, w_034_013, w_034_015, w_034_016, w_034_017, w_034_018, w_034_019, w_034_020, w_034_021, w_034_022, w_034_023, w_034_024, w_034_025, w_034_026, w_034_027, w_034_028, w_034_029, w_034_030, w_034_031, w_034_032, w_034_033, w_034_034, w_034_035, w_034_036, w_034_037, w_034_038, w_034_039, w_034_040, w_034_041, w_034_042, w_034_043, w_034_044, w_034_045, w_034_046, w_034_047, w_034_048, w_034_049, w_034_050, w_034_051, w_034_052, w_034_053, w_034_054, w_034_055, w_034_056, w_034_057, w_034_058, w_034_059, w_034_060, w_034_061, w_034_062, w_034_063, w_034_064, w_034_065, w_034_066, w_034_067, w_034_068, w_034_069, w_034_070, w_034_071, w_034_072, w_034_073, w_034_074, w_034_075;
  wire w_035_000, w_035_001, w_035_002, w_035_003, w_035_004, w_035_005, w_035_006, w_035_007, w_035_008, w_035_009, w_035_010, w_035_012, w_035_013, w_035_014, w_035_015, w_035_016, w_035_017, w_035_018, w_035_019, w_035_020, w_035_021, w_035_022, w_035_023, w_035_024, w_035_025, w_035_027, w_035_028, w_035_029, w_035_030, w_035_031, w_035_032, w_035_034, w_035_035, w_035_036, w_035_037, w_035_039, w_035_040, w_035_042, w_035_043, w_035_044, w_035_045, w_035_046, w_035_047, w_035_048, w_035_049, w_035_050, w_035_051, w_035_052, w_035_053, w_035_054, w_035_055, w_035_056, w_035_057, w_035_059, w_035_060, w_035_061, w_035_062, w_035_063, w_035_064, w_035_065, w_035_066, w_035_067, w_035_068, w_035_069, w_035_070, w_035_072, w_035_073, w_035_074, w_035_076, w_035_077, w_035_078, w_035_080, w_035_081, w_035_082, w_035_083, w_035_084, w_035_085, w_035_087, w_035_088, w_035_090, w_035_091, w_035_092, w_035_093, w_035_094, w_035_095, w_035_096, w_035_097, w_035_098, w_035_099, w_035_100, w_035_101, w_035_102, w_035_103, w_035_104, w_035_105, w_035_106, w_035_107, w_035_108, w_035_110, w_035_111, w_035_112, w_035_114, w_035_115, w_035_116, w_035_117, w_035_118, w_035_119, w_035_120, w_035_121, w_035_122, w_035_124, w_035_125, w_035_126, w_035_127;
  wire w_036_002, w_036_004, w_036_006, w_036_009, w_036_010, w_036_011, w_036_012, w_036_014, w_036_018, w_036_019, w_036_020, w_036_022, w_036_023, w_036_024, w_036_026, w_036_028, w_036_029, w_036_032, w_036_033, w_036_034, w_036_035, w_036_037, w_036_039, w_036_042, w_036_043, w_036_044, w_036_046, w_036_047, w_036_049, w_036_050, w_036_052, w_036_053, w_036_058, w_036_059, w_036_060, w_036_062, w_036_063, w_036_064, w_036_066, w_036_068, w_036_071, w_036_072, w_036_073, w_036_074, w_036_075, w_036_076, w_036_078, w_036_079, w_036_080, w_036_082, w_036_083, w_036_084, w_036_085, w_036_087, w_036_088, w_036_090, w_036_091, w_036_093, w_036_094, w_036_096, w_036_097, w_036_099, w_036_101, w_036_103, w_036_109, w_036_110, w_036_112, w_036_114, w_036_117, w_036_118, w_036_120, w_036_121, w_036_123, w_036_125, w_036_126, w_036_128, w_036_129, w_036_131, w_036_132, w_036_134, w_036_136, w_036_138, w_036_139, w_036_140, w_036_141, w_036_144, w_036_146, w_036_148, w_036_151, w_036_153, w_036_154, w_036_156, w_036_157, w_036_158, w_036_160, w_036_161, w_036_162, w_036_163, w_036_164, w_036_165, w_036_166, w_036_170, w_036_173, w_036_175, w_036_177, w_036_178, w_036_179, w_036_180, w_036_182, w_036_186, w_036_188, w_036_190, w_036_191, w_036_192, w_036_194, w_036_197, w_036_200, w_036_201, w_036_206, w_036_207, w_036_211, w_036_215, w_036_217, w_036_221, w_036_224, w_036_227, w_036_229, w_036_231, w_036_232, w_036_235, w_036_237, w_036_239, w_036_240, w_036_241, w_036_242, w_036_243, w_036_244, w_036_245, w_036_247, w_036_251, w_036_255, w_036_256, w_036_257, w_036_258, w_036_259, w_036_261, w_036_262, w_036_265, w_036_266, w_036_267, w_036_269, w_036_271, w_036_272, w_036_273, w_036_274, w_036_276, w_036_277, w_036_278, w_036_281, w_036_282, w_036_283, w_036_284, w_036_286, w_036_289, w_036_291, w_036_294, w_036_295, w_036_296, w_036_297, w_036_298, w_036_299, w_036_302, w_036_304, w_036_305, w_036_307, w_036_309, w_036_310, w_036_311, w_036_312, w_036_313, w_036_314, w_036_318, w_036_319, w_036_322, w_036_323, w_036_324, w_036_327, w_036_328, w_036_330, w_036_335, w_036_336, w_036_348, w_036_349, w_036_350, w_036_354, w_036_357, w_036_359, w_036_368, w_036_376, w_036_386, w_036_393, w_036_395, w_036_400, w_036_404, w_036_408, w_036_412, w_036_430, w_036_432, w_036_440, w_036_444, w_036_447, w_036_449, w_036_455, w_036_459, w_036_461;
  wire w_037_001, w_037_002, w_037_003, w_037_008, w_037_010, w_037_011, w_037_013, w_037_015, w_037_017, w_037_020, w_037_021, w_037_022, w_037_023, w_037_024, w_037_026, w_037_028, w_037_030, w_037_031, w_037_032, w_037_033, w_037_034, w_037_036, w_037_041, w_037_042, w_037_044, w_037_045, w_037_047, w_037_048, w_037_049, w_037_050, w_037_051, w_037_055, w_037_059, w_037_060, w_037_062, w_037_063, w_037_064, w_037_066, w_037_068, w_037_070, w_037_071, w_037_073, w_037_074, w_037_075, w_037_076, w_037_077, w_037_081, w_037_082, w_037_083, w_037_085, w_037_086, w_037_087, w_037_088, w_037_089, w_037_093, w_037_095, w_037_096, w_037_097, w_037_100, w_037_101, w_037_103, w_037_104, w_037_105, w_037_110, w_037_115, w_037_117, w_037_119, w_037_120, w_037_122, w_037_123, w_037_124, w_037_129, w_037_130, w_037_131, w_037_132, w_037_133, w_037_140, w_037_141, w_037_146, w_037_147, w_037_149, w_037_150, w_037_152, w_037_153, w_037_154, w_037_155, w_037_157, w_037_158, w_037_162, w_037_164, w_037_166, w_037_168, w_037_169, w_037_172, w_037_173, w_037_177, w_037_185, w_037_186, w_037_188, w_037_189, w_037_195, w_037_198, w_037_200, w_037_201, w_037_203, w_037_206, w_037_207, w_037_208, w_037_210, w_037_211, w_037_212, w_037_217, w_037_218, w_037_221, w_037_223, w_037_225, w_037_228, w_037_229, w_037_231, w_037_232, w_037_233, w_037_234, w_037_235, w_037_236, w_037_242, w_037_245, w_037_246, w_037_248, w_037_249, w_037_251, w_037_253, w_037_257, w_037_258, w_037_261, w_037_262, w_037_263, w_037_266, w_037_267, w_037_268, w_037_273, w_037_277, w_037_278, w_037_279, w_037_280, w_037_285, w_037_286, w_037_287, w_037_293, w_037_295, w_037_300, w_037_301, w_037_302, w_037_303, w_037_305, w_037_308, w_037_309, w_037_310, w_037_312, w_037_313, w_037_314, w_037_315, w_037_316, w_037_318, w_037_319, w_037_320, w_037_323, w_037_330, w_037_332, w_037_333, w_037_336, w_037_338, w_037_339, w_037_343, w_037_345, w_037_346, w_037_349, w_037_350, w_037_351;
  wire w_038_000, w_038_002, w_038_005, w_038_011, w_038_012, w_038_016, w_038_018, w_038_019, w_038_020, w_038_021, w_038_022, w_038_024, w_038_025, w_038_032, w_038_033, w_038_043, w_038_044, w_038_047, w_038_051, w_038_052, w_038_053, w_038_054, w_038_055, w_038_059, w_038_061, w_038_064, w_038_065, w_038_066, w_038_067, w_038_068, w_038_070, w_038_074, w_038_076, w_038_077, w_038_079, w_038_082, w_038_085, w_038_087, w_038_090, w_038_093, w_038_095, w_038_096, w_038_097, w_038_099, w_038_100, w_038_103, w_038_106, w_038_108, w_038_111, w_038_115, w_038_116, w_038_117, w_038_120, w_038_121, w_038_123, w_038_132, w_038_134, w_038_135, w_038_138, w_038_140, w_038_142, w_038_143, w_038_144, w_038_146, w_038_147, w_038_148, w_038_149, w_038_150, w_038_151, w_038_152, w_038_157, w_038_160, w_038_162, w_038_163, w_038_164, w_038_169, w_038_173, w_038_176, w_038_178, w_038_182, w_038_185, w_038_188, w_038_193, w_038_196, w_038_200, w_038_203, w_038_211, w_038_225, w_038_234, w_038_240, w_038_247, w_038_255, w_038_256, w_038_260, w_038_265, w_038_268, w_038_275, w_038_285, w_038_288, w_038_290, w_038_297, w_038_298, w_038_299, w_038_302, w_038_303, w_038_304, w_038_308, w_038_311, w_038_315, w_038_317, w_038_321, w_038_322, w_038_325, w_038_331, w_038_333, w_038_337, w_038_340, w_038_358, w_038_359, w_038_365, w_038_368, w_038_370, w_038_377, w_038_383, w_038_385, w_038_386, w_038_396, w_038_397, w_038_402, w_038_405, w_038_415, w_038_418, w_038_423, w_038_429, w_038_431, w_038_434, w_038_435, w_038_447, w_038_454, w_038_455, w_038_456, w_038_457, w_038_458, w_038_462, w_038_465, w_038_467, w_038_468, w_038_469, w_038_471, w_038_472, w_038_484, w_038_486, w_038_489, w_038_491, w_038_495, w_038_496, w_038_498, w_038_499, w_038_501, w_038_503, w_038_504, w_038_505, w_038_508, w_038_512, w_038_515, w_038_516, w_038_521, w_038_526, w_038_531, w_038_532, w_038_538, w_038_542, w_038_546, w_038_548, w_038_549, w_038_550, w_038_551, w_038_559, w_038_565, w_038_567, w_038_575, w_038_588, w_038_589, w_038_590, w_038_591, w_038_597, w_038_598, w_038_600, w_038_601, w_038_602, w_038_604, w_038_606, w_038_610, w_038_618, w_038_624, w_038_625, w_038_626, w_038_627, w_038_628, w_038_629, w_038_630, w_038_631, w_038_632;
  wire w_039_003, w_039_005, w_039_007, w_039_010, w_039_014, w_039_016, w_039_024, w_039_029, w_039_030, w_039_032, w_039_033, w_039_035, w_039_037, w_039_039, w_039_040, w_039_043, w_039_046, w_039_050, w_039_051, w_039_052, w_039_054, w_039_055, w_039_057, w_039_061, w_039_063, w_039_064, w_039_066, w_039_068, w_039_069, w_039_072, w_039_073, w_039_076, w_039_078, w_039_079, w_039_082, w_039_085, w_039_088, w_039_089, w_039_092, w_039_093, w_039_095, w_039_099, w_039_103, w_039_104, w_039_108, w_039_111, w_039_117, w_039_119, w_039_121, w_039_127, w_039_141, w_039_143, w_039_145, w_039_148, w_039_152, w_039_155, w_039_158, w_039_160, w_039_161, w_039_167, w_039_170, w_039_173, w_039_175, w_039_182, w_039_185, w_039_187, w_039_197, w_039_203, w_039_206, w_039_208, w_039_213, w_039_214, w_039_218, w_039_219, w_039_221, w_039_228, w_039_231, w_039_240, w_039_242, w_039_256, w_039_258, w_039_260, w_039_263, w_039_264, w_039_267, w_039_278, w_039_280, w_039_289, w_039_295, w_039_300, w_039_301, w_039_302, w_039_306, w_039_309, w_039_317, w_039_318, w_039_324, w_039_327, w_039_329, w_039_348, w_039_351, w_039_352, w_039_360, w_039_361, w_039_367, w_039_368, w_039_370, w_039_371, w_039_372, w_039_373, w_039_374, w_039_377, w_039_380, w_039_383, w_039_395, w_039_396, w_039_401, w_039_404, w_039_406, w_039_413, w_039_415, w_039_421, w_039_422, w_039_424, w_039_425, w_039_427, w_039_428, w_039_429, w_039_432, w_039_440, w_039_446, w_039_448, w_039_459, w_039_466, w_039_470, w_039_471, w_039_478, w_039_492, w_039_493, w_039_495, w_039_505, w_039_506, w_039_510, w_039_513, w_039_515, w_039_518, w_039_519, w_039_522, w_039_524, w_039_527, w_039_528, w_039_530, w_039_534, w_039_536, w_039_537, w_039_538, w_039_539, w_039_543, w_039_544, w_039_550, w_039_552, w_039_553, w_039_559, w_039_561, w_039_567, w_039_569, w_039_571, w_039_578, w_039_580, w_039_581, w_039_586, w_039_588, w_039_598, w_039_599, w_039_600, w_039_602, w_039_604, w_039_606, w_039_609, w_039_612, w_039_616, w_039_620, w_039_621, w_039_625, w_039_634, w_039_646, w_039_648, w_039_650, w_039_652, w_039_656, w_039_657, w_039_658, w_039_667, w_039_668, w_039_676, w_039_680, w_039_681, w_039_697, w_039_699, w_039_706, w_039_708, w_039_710, w_039_713, w_039_714, w_039_718, w_039_719;
  wire w_040_000, w_040_004, w_040_005, w_040_008, w_040_012, w_040_013, w_040_014, w_040_015, w_040_017, w_040_019, w_040_021, w_040_027, w_040_031, w_040_032, w_040_039, w_040_040, w_040_043, w_040_044, w_040_045, w_040_047, w_040_049, w_040_050, w_040_051, w_040_053, w_040_054, w_040_063, w_040_065, w_040_067, w_040_068, w_040_070, w_040_071, w_040_072, w_040_077, w_040_080, w_040_083, w_040_086, w_040_088, w_040_090, w_040_091, w_040_096, w_040_098, w_040_099, w_040_101, w_040_102, w_040_106, w_040_119, w_040_120, w_040_123, w_040_129, w_040_132, w_040_133, w_040_139, w_040_146, w_040_147, w_040_149, w_040_163, w_040_164, w_040_166, w_040_174, w_040_180, w_040_184, w_040_193, w_040_196, w_040_210, w_040_219, w_040_221, w_040_225, w_040_228, w_040_234, w_040_235, w_040_238, w_040_241, w_040_243, w_040_246, w_040_252, w_040_254, w_040_257, w_040_268, w_040_278, w_040_281, w_040_283, w_040_286, w_040_288, w_040_294, w_040_295, w_040_298, w_040_299, w_040_304, w_040_309, w_040_311, w_040_312, w_040_316, w_040_317, w_040_318, w_040_322, w_040_324, w_040_325, w_040_327, w_040_328, w_040_340, w_040_343, w_040_346, w_040_348, w_040_353, w_040_356, w_040_357, w_040_358, w_040_360, w_040_361, w_040_366, w_040_367, w_040_371, w_040_373, w_040_382, w_040_386, w_040_393, w_040_395, w_040_404, w_040_405, w_040_409, w_040_415, w_040_423, w_040_425, w_040_427, w_040_428, w_040_430, w_040_432, w_040_433, w_040_439, w_040_440, w_040_441, w_040_442, w_040_449, w_040_462, w_040_463, w_040_464, w_040_468, w_040_469, w_040_475, w_040_478, w_040_479, w_040_480, w_040_481, w_040_482, w_040_484, w_040_486, w_040_488, w_040_493, w_040_497, w_040_501, w_040_505, w_040_509, w_040_514, w_040_515, w_040_519, w_040_520, w_040_521, w_040_524, w_040_539, w_040_542, w_040_549, w_040_551, w_040_553, w_040_554, w_040_555, w_040_558, w_040_565, w_040_568, w_040_571, w_040_582, w_040_583, w_040_592, w_040_594, w_040_599, w_040_601, w_040_607, w_040_609, w_040_611, w_040_614, w_040_616, w_040_617, w_040_623, w_040_630, w_040_632, w_040_639, w_040_644, w_040_646, w_040_660, w_040_663, w_040_667, w_040_670, w_040_682, w_040_689, w_040_691, w_040_692, w_040_693, w_040_698, w_040_699, w_040_704, w_040_705, w_040_713, w_040_719, w_040_720, w_040_721, w_040_722, w_040_723, w_040_724, w_040_725, w_040_726, w_040_727, w_040_728, w_040_729, w_040_730;
  wire w_041_007, w_041_010, w_041_011, w_041_013, w_041_016, w_041_023, w_041_024, w_041_026, w_041_029, w_041_032, w_041_035, w_041_036, w_041_037, w_041_038, w_041_041, w_041_046, w_041_048, w_041_051, w_041_052, w_041_053, w_041_054, w_041_055, w_041_057, w_041_060, w_041_062, w_041_070, w_041_073, w_041_077, w_041_079, w_041_081, w_041_083, w_041_086, w_041_088, w_041_090, w_041_097, w_041_100, w_041_102, w_041_104, w_041_106, w_041_110, w_041_113, w_041_116, w_041_117, w_041_128, w_041_131, w_041_138, w_041_154, w_041_160, w_041_166, w_041_172, w_041_178, w_041_181, w_041_185, w_041_189, w_041_194, w_041_197, w_041_206, w_041_212, w_041_220, w_041_226, w_041_228, w_041_231, w_041_234, w_041_241, w_041_243, w_041_244, w_041_246, w_041_248, w_041_257, w_041_263, w_041_275, w_041_276, w_041_279, w_041_282, w_041_288, w_041_293, w_041_298, w_041_300, w_041_304, w_041_305, w_041_306, w_041_315, w_041_326, w_041_334, w_041_336, w_041_337, w_041_338, w_041_339, w_041_340, w_041_342, w_041_345, w_041_346, w_041_349, w_041_354, w_041_355, w_041_359, w_041_378, w_041_380, w_041_389, w_041_392, w_041_397, w_041_399, w_041_403, w_041_408, w_041_409, w_041_412, w_041_414, w_041_429, w_041_432, w_041_433, w_041_434, w_041_439, w_041_441, w_041_444, w_041_446, w_041_453, w_041_457, w_041_460, w_041_463, w_041_476, w_041_482, w_041_485, w_041_488, w_041_489, w_041_491, w_041_494, w_041_496, w_041_497, w_041_499, w_041_504, w_041_507, w_041_510, w_041_511, w_041_512, w_041_513, w_041_515, w_041_524, w_041_525, w_041_528, w_041_529, w_041_531, w_041_532, w_041_535, w_041_537, w_041_541, w_041_548, w_041_549, w_041_561, w_041_576, w_041_579, w_041_581, w_041_583, w_041_587, w_041_589, w_041_593, w_041_594, w_041_604, w_041_606, w_041_610, w_041_614, w_041_618, w_041_623, w_041_625, w_041_627, w_041_628, w_041_630, w_041_632, w_041_647, w_041_659, w_041_661, w_041_663, w_041_664, w_041_665, w_041_668, w_041_670, w_041_673, w_041_676, w_041_683, w_041_685, w_041_692, w_041_698, w_041_713, w_041_714, w_041_721;
  wire w_042_000, w_042_001, w_042_002, w_042_005, w_042_006, w_042_008, w_042_010, w_042_012, w_042_013, w_042_018, w_042_023, w_042_024, w_042_025, w_042_026, w_042_034, w_042_035, w_042_036, w_042_038, w_042_039, w_042_041, w_042_043, w_042_044, w_042_045, w_042_050, w_042_052, w_042_056, w_042_057, w_042_059, w_042_061, w_042_062, w_042_066, w_042_071, w_042_072, w_042_076, w_042_077, w_042_081, w_042_082, w_042_084, w_042_090, w_042_092, w_042_094, w_042_095, w_042_099, w_042_101, w_042_102, w_042_103, w_042_104, w_042_109, w_042_110, w_042_111, w_042_112, w_042_113, w_042_116, w_042_117, w_042_121, w_042_123, w_042_124, w_042_125, w_042_126, w_042_127, w_042_130, w_042_132, w_042_133, w_042_134, w_042_135, w_042_138, w_042_139, w_042_144, w_042_146, w_042_147, w_042_148, w_042_150, w_042_152, w_042_155, w_042_156, w_042_157, w_042_158, w_042_159, w_042_162, w_042_165, w_042_169, w_042_171, w_042_172, w_042_178, w_042_180, w_042_181, w_042_182, w_042_184, w_042_185, w_042_186, w_042_191, w_042_192, w_042_194, w_042_195, w_042_197, w_042_198, w_042_199, w_042_201, w_042_203, w_042_206, w_042_209, w_042_215, w_042_217, w_042_219, w_042_220, w_042_222, w_042_226, w_042_227, w_042_229, w_042_232, w_042_233, w_042_237, w_042_252, w_042_255, w_042_257, w_042_258, w_042_260, w_042_261, w_042_264, w_042_265, w_042_267, w_042_268, w_042_271, w_042_272, w_042_275, w_042_276, w_042_278, w_042_279, w_042_281, w_042_282, w_042_286, w_042_288, w_042_290, w_042_292, w_042_293, w_042_295, w_042_297, w_042_298, w_042_304, w_042_305, w_042_307, w_042_309, w_042_310, w_042_311, w_042_312, w_042_316, w_042_317, w_042_318, w_042_319, w_042_320, w_042_321, w_042_323, w_042_325, w_042_327, w_042_328, w_042_331, w_042_332, w_042_334, w_042_339, w_042_340, w_042_343, w_042_346, w_042_356, w_042_358, w_042_359, w_042_362, w_042_367, w_042_368, w_042_369, w_042_377, w_042_384, w_042_385, w_042_389, w_042_401, w_042_402, w_042_404, w_042_406, w_042_409, w_042_413, w_042_414, w_042_415, w_042_422, w_042_423, w_042_427, w_042_428, w_042_432, w_042_433, w_042_437, w_042_443, w_042_451, w_042_453, w_042_455, w_042_456;
  wire w_043_000, w_043_001, w_043_002, w_043_003, w_043_004, w_043_005, w_043_006, w_043_007, w_043_008, w_043_009, w_043_010, w_043_011, w_043_012, w_043_013, w_043_014, w_043_015, w_043_016, w_043_017, w_043_018, w_043_019, w_043_020, w_043_021, w_043_022, w_043_023, w_043_024, w_043_025, w_043_026, w_043_027, w_043_028, w_043_029, w_043_030, w_043_031, w_043_032, w_043_033, w_043_034, w_043_035, w_043_036, w_043_037, w_043_038, w_043_039, w_043_040, w_043_041, w_043_042, w_043_043, w_043_044, w_043_045, w_043_046, w_043_047;
  wire w_044_000, w_044_002, w_044_013, w_044_014, w_044_019, w_044_021, w_044_022, w_044_026, w_044_027, w_044_029, w_044_030, w_044_033, w_044_036, w_044_040, w_044_041, w_044_046, w_044_048, w_044_050, w_044_054, w_044_055, w_044_058, w_044_062, w_044_070, w_044_072, w_044_080, w_044_082, w_044_093, w_044_098, w_044_100, w_044_109, w_044_110, w_044_115, w_044_119, w_044_122, w_044_127, w_044_128, w_044_137, w_044_139, w_044_154, w_044_158, w_044_159, w_044_160, w_044_165, w_044_169, w_044_175, w_044_180, w_044_181, w_044_191, w_044_195, w_044_197, w_044_199, w_044_201, w_044_206, w_044_209, w_044_219, w_044_223, w_044_225, w_044_229, w_044_243, w_044_248, w_044_261, w_044_267, w_044_268, w_044_273, w_044_276, w_044_284, w_044_286, w_044_289, w_044_290, w_044_292, w_044_293, w_044_295, w_044_296, w_044_301, w_044_303, w_044_306, w_044_312, w_044_322, w_044_331, w_044_332, w_044_335, w_044_338, w_044_341, w_044_344, w_044_347, w_044_348, w_044_366, w_044_367, w_044_371, w_044_373, w_044_375, w_044_377, w_044_384, w_044_390, w_044_395, w_044_398, w_044_402, w_044_403, w_044_405, w_044_407, w_044_414, w_044_418, w_044_419, w_044_424, w_044_435, w_044_447, w_044_449, w_044_450, w_044_452, w_044_454, w_044_457, w_044_458, w_044_459, w_044_460, w_044_461, w_044_465, w_044_473, w_044_475, w_044_487, w_044_496, w_044_497, w_044_499, w_044_500, w_044_502, w_044_507, w_044_510, w_044_514, w_044_518, w_044_521, w_044_532, w_044_534, w_044_535, w_044_540, w_044_544, w_044_559, w_044_562, w_044_563, w_044_564, w_044_569, w_044_571, w_044_573, w_044_574, w_044_577, w_044_583, w_044_587, w_044_588, w_044_589, w_044_598, w_044_599, w_044_603, w_044_608, w_044_610, w_044_611, w_044_616, w_044_628, w_044_632, w_044_643, w_044_646, w_044_650, w_044_652, w_044_653, w_044_657, w_044_658, w_044_662, w_044_663, w_044_666, w_044_670, w_044_673, w_044_675, w_044_681, w_044_684, w_044_686, w_044_687, w_044_689, w_044_690, w_044_691, w_044_694, w_044_705, w_044_710, w_044_712, w_044_713, w_044_719, w_044_721, w_044_722, w_044_723, w_044_740, w_044_743, w_044_746;
  wire w_045_000, w_045_001, w_045_002, w_045_003, w_045_005, w_045_006, w_045_007, w_045_009, w_045_012, w_045_013, w_045_014, w_045_016, w_045_017, w_045_020, w_045_023, w_045_024, w_045_026, w_045_029, w_045_034, w_045_038, w_045_039, w_045_041, w_045_043, w_045_044, w_045_047, w_045_048, w_045_049, w_045_050, w_045_052, w_045_055, w_045_057, w_045_060, w_045_063, w_045_067, w_045_068, w_045_069, w_045_071, w_045_074, w_045_075, w_045_083, w_045_084, w_045_088, w_045_091, w_045_092, w_045_100, w_045_102, w_045_105, w_045_106, w_045_108, w_045_109, w_045_117, w_045_118, w_045_124, w_045_126, w_045_129, w_045_130, w_045_131, w_045_138, w_045_139, w_045_144, w_045_148, w_045_149, w_045_151, w_045_157, w_045_158, w_045_160, w_045_161, w_045_166, w_045_167, w_045_168, w_045_169, w_045_170, w_045_172, w_045_174, w_045_176, w_045_177, w_045_180, w_045_181, w_045_182, w_045_186, w_045_189, w_045_191, w_045_196, w_045_197, w_045_198, w_045_199, w_045_204, w_045_205, w_045_206, w_045_210, w_045_212, w_045_215, w_045_219, w_045_220, w_045_224, w_045_225, w_045_226, w_045_227, w_045_228, w_045_230, w_045_231, w_045_235, w_045_239, w_045_242, w_045_245, w_045_255, w_045_258, w_045_259, w_045_260, w_045_264, w_045_265, w_045_266, w_045_267, w_045_268, w_045_269, w_045_270, w_045_271, w_045_272, w_045_274, w_045_276, w_045_277, w_045_280, w_045_282, w_045_283, w_045_284, w_045_286, w_045_287, w_045_289, w_045_290, w_045_291, w_045_292, w_045_293, w_045_294, w_045_296, w_045_300, w_045_304, w_045_305, w_045_307, w_045_308, w_045_310, w_045_311, w_045_314, w_045_315, w_045_317, w_045_319, w_045_321, w_045_323, w_045_326, w_045_327, w_045_330, w_045_331, w_045_332, w_045_333, w_045_334, w_045_335, w_045_336, w_045_337, w_045_338, w_045_344, w_045_345, w_045_348, w_045_353, w_045_358, w_045_359, w_045_361, w_045_362, w_045_366, w_045_367, w_045_368, w_045_369, w_045_375, w_045_378, w_045_379, w_045_381, w_045_386, w_045_388, w_045_389, w_045_390, w_045_400, w_045_401, w_045_405, w_045_407, w_045_410, w_045_411, w_045_412, w_045_413, w_045_414, w_045_418, w_045_419, w_045_420, w_045_421, w_045_422, w_045_423, w_045_424, w_045_425, w_045_426, w_045_427, w_045_429;
  wire w_046_002, w_046_009, w_046_010, w_046_013, w_046_015, w_046_023, w_046_024, w_046_025, w_046_028, w_046_029, w_046_031, w_046_033, w_046_037, w_046_039, w_046_041, w_046_042, w_046_047, w_046_050, w_046_052, w_046_057, w_046_058, w_046_059, w_046_061, w_046_062, w_046_068, w_046_073, w_046_074, w_046_082, w_046_085, w_046_092, w_046_096, w_046_097, w_046_099, w_046_100, w_046_101, w_046_104, w_046_106, w_046_110, w_046_118, w_046_120, w_046_121, w_046_127, w_046_129, w_046_132, w_046_137, w_046_143, w_046_164, w_046_168, w_046_171, w_046_172, w_046_174, w_046_176, w_046_184, w_046_189, w_046_194, w_046_196, w_046_197, w_046_201, w_046_209, w_046_210, w_046_211, w_046_222, w_046_229, w_046_230, w_046_232, w_046_234, w_046_236, w_046_238, w_046_240, w_046_246, w_046_247, w_046_248, w_046_250, w_046_255, w_046_261, w_046_263, w_046_264, w_046_267, w_046_270, w_046_272, w_046_279, w_046_284, w_046_288, w_046_292, w_046_294, w_046_297, w_046_298, w_046_299, w_046_300, w_046_302, w_046_303, w_046_304, w_046_314, w_046_318, w_046_319, w_046_323, w_046_330, w_046_334, w_046_336, w_046_338, w_046_339, w_046_341, w_046_346, w_046_351, w_046_356, w_046_360, w_046_372, w_046_373, w_046_377, w_046_387, w_046_389, w_046_390, w_046_394, w_046_397, w_046_401, w_046_414, w_046_422, w_046_425, w_046_427, w_046_429, w_046_432, w_046_435, w_046_436, w_046_443, w_046_447, w_046_450, w_046_452, w_046_456, w_046_459, w_046_463, w_046_467, w_046_472, w_046_477, w_046_478, w_046_480, w_046_483, w_046_484, w_046_494, w_046_496, w_046_509, w_046_515, w_046_516, w_046_517, w_046_525, w_046_526, w_046_532, w_046_545, w_046_551, w_046_561, w_046_562, w_046_564, w_046_571, w_046_575, w_046_576, w_046_580, w_046_583, w_046_593, w_046_598, w_046_599, w_046_604, w_046_606, w_046_608, w_046_609, w_046_611, w_046_612, w_046_616, w_046_619, w_046_620, w_046_625, w_046_627, w_046_630, w_046_631, w_046_632, w_046_637, w_046_646, w_046_647, w_046_655, w_046_659, w_046_660, w_046_662, w_046_677, w_046_686, w_046_698, w_046_699, w_046_702, w_046_704, w_046_712;
  wire w_047_001, w_047_002, w_047_005, w_047_006, w_047_007, w_047_008, w_047_013, w_047_014, w_047_018, w_047_021, w_047_023, w_047_024, w_047_031, w_047_032, w_047_033, w_047_038, w_047_040, w_047_042, w_047_045, w_047_047, w_047_049, w_047_050, w_047_051, w_047_054, w_047_065, w_047_070, w_047_072, w_047_073, w_047_077, w_047_080, w_047_087, w_047_088, w_047_090, w_047_099, w_047_105, w_047_106, w_047_107, w_047_113, w_047_115, w_047_116, w_047_118, w_047_119, w_047_121, w_047_124, w_047_125, w_047_126, w_047_129, w_047_132, w_047_134, w_047_136, w_047_137, w_047_139, w_047_140, w_047_141, w_047_142, w_047_147, w_047_148, w_047_152, w_047_154, w_047_155, w_047_158, w_047_174, w_047_177, w_047_185, w_047_188, w_047_191, w_047_192, w_047_197, w_047_199, w_047_201, w_047_205, w_047_206, w_047_207, w_047_208, w_047_209, w_047_210, w_047_211, w_047_214, w_047_215, w_047_219, w_047_220, w_047_221, w_047_224, w_047_225, w_047_229, w_047_230, w_047_232, w_047_237, w_047_238, w_047_239, w_047_245, w_047_246, w_047_248, w_047_249, w_047_251, w_047_254, w_047_255, w_047_256, w_047_263, w_047_265, w_047_267, w_047_268, w_047_270, w_047_273, w_047_275, w_047_276, w_047_277, w_047_279, w_047_280, w_047_283, w_047_287, w_047_288, w_047_290, w_047_291, w_047_294, w_047_295, w_047_298, w_047_299, w_047_305, w_047_306, w_047_307, w_047_309, w_047_311, w_047_317, w_047_318, w_047_320, w_047_323, w_047_325, w_047_327, w_047_329, w_047_330, w_047_340, w_047_341, w_047_342, w_047_350, w_047_359, w_047_360, w_047_362, w_047_367, w_047_370, w_047_379, w_047_383, w_047_390, w_047_394, w_047_396, w_047_399, w_047_404, w_047_407, w_047_413, w_047_419, w_047_420, w_047_422, w_047_428, w_047_436, w_047_443, w_047_454, w_047_458, w_047_465, w_047_469;
  wire w_048_000, w_048_001, w_048_002, w_048_003, w_048_004, w_048_005, w_048_006, w_048_007, w_048_008, w_048_009, w_048_010, w_048_011, w_048_012, w_048_013, w_048_014, w_048_015, w_048_016, w_048_017, w_048_018, w_048_019;
  wire w_049_002, w_049_003, w_049_004, w_049_005, w_049_006, w_049_009, w_049_011, w_049_012, w_049_016, w_049_017, w_049_018, w_049_019, w_049_020, w_049_021, w_049_022, w_049_023, w_049_024, w_049_025, w_049_026, w_049_029, w_049_033, w_049_035, w_049_036, w_049_041, w_049_045, w_049_047, w_049_049, w_049_060, w_049_065, w_049_066, w_049_070, w_049_074, w_049_076, w_049_079, w_049_081, w_049_083, w_049_093, w_049_095, w_049_101, w_049_104, w_049_107, w_049_110, w_049_111, w_049_112, w_049_116, w_049_119, w_049_120, w_049_121, w_049_124, w_049_130, w_049_131, w_049_134, w_049_135, w_049_140, w_049_144, w_049_153, w_049_154, w_049_161, w_049_162, w_049_164, w_049_165, w_049_166, w_049_168, w_049_171, w_049_172, w_049_174, w_049_175, w_049_177, w_049_178, w_049_179, w_049_182, w_049_184, w_049_187, w_049_189, w_049_190, w_049_192, w_049_200, w_049_202, w_049_204, w_049_207, w_049_209, w_049_210, w_049_217, w_049_220, w_049_222, w_049_223, w_049_231, w_049_232, w_049_233, w_049_236, w_049_237, w_049_238, w_049_239, w_049_240, w_049_246, w_049_249, w_049_252, w_049_253, w_049_254, w_049_256, w_049_259, w_049_260, w_049_263, w_049_267, w_049_268, w_049_269, w_049_271, w_049_272, w_049_277, w_049_278, w_049_279, w_049_280, w_049_281, w_049_282, w_049_285, w_049_288, w_049_290, w_049_292, w_049_294, w_049_299, w_049_303, w_049_304, w_049_305, w_049_309, w_049_312, w_049_313, w_049_320, w_049_322, w_049_324, w_049_334, w_049_335, w_049_337, w_049_338, w_049_341, w_049_342, w_049_347, w_049_348, w_049_358, w_049_362, w_049_363, w_049_372, w_049_373, w_049_386, w_049_389, w_049_397, w_049_411;
  wire w_050_004, w_050_007, w_050_008, w_050_009, w_050_010, w_050_011, w_050_012, w_050_016, w_050_017, w_050_021, w_050_024, w_050_027, w_050_030, w_050_031, w_050_032, w_050_034, w_050_035, w_050_036, w_050_037, w_050_041, w_050_042, w_050_045, w_050_046, w_050_047, w_050_048, w_050_050, w_050_054, w_050_056, w_050_058, w_050_062, w_050_064, w_050_069, w_050_071, w_050_072, w_050_079, w_050_080, w_050_082, w_050_085, w_050_091, w_050_093, w_050_099, w_050_101, w_050_103, w_050_105, w_050_106, w_050_110, w_050_112, w_050_117, w_050_119, w_050_120, w_050_121, w_050_123, w_050_127, w_050_130, w_050_131, w_050_133, w_050_135, w_050_136, w_050_138, w_050_141, w_050_148, w_050_149, w_050_152, w_050_161, w_050_164, w_050_175, w_050_177, w_050_186, w_050_199, w_050_205, w_050_207, w_050_211, w_050_222, w_050_226, w_050_234, w_050_236, w_050_237, w_050_238, w_050_242, w_050_247, w_050_257, w_050_259, w_050_263, w_050_264, w_050_266, w_050_267, w_050_271, w_050_274, w_050_280, w_050_292, w_050_295, w_050_305, w_050_306, w_050_309, w_050_312, w_050_317, w_050_322, w_050_323, w_050_333, w_050_334, w_050_344, w_050_348, w_050_359, w_050_363, w_050_365, w_050_367, w_050_373, w_050_376, w_050_377, w_050_384, w_050_385, w_050_386, w_050_388, w_050_392, w_050_398, w_050_399, w_050_401, w_050_404, w_050_405, w_050_406, w_050_407, w_050_408, w_050_412, w_050_415, w_050_416, w_050_417, w_050_427, w_050_435, w_050_437, w_050_440, w_050_446, w_050_454, w_050_460, w_050_461, w_050_470, w_050_475, w_050_479, w_050_480, w_050_488, w_050_493, w_050_500, w_050_510, w_050_514, w_050_520, w_050_526, w_050_532, w_050_533, w_050_534, w_050_537, w_050_543, w_050_546, w_050_570, w_050_571, w_050_573, w_050_578, w_050_584, w_050_589, w_050_593, w_050_597, w_050_602, w_050_610, w_050_611, w_050_612, w_050_621, w_050_626, w_050_627, w_050_630, w_050_646;
  wire w_051_003, w_051_005, w_051_006, w_051_008, w_051_009, w_051_011, w_051_013, w_051_014, w_051_017, w_051_019, w_051_021, w_051_023, w_051_024, w_051_025, w_051_027, w_051_028, w_051_031, w_051_033, w_051_036, w_051_037, w_051_041, w_051_044, w_051_045, w_051_051, w_051_052, w_051_053, w_051_055, w_051_061, w_051_062, w_051_063, w_051_067, w_051_069, w_051_073, w_051_074, w_051_075, w_051_078, w_051_080, w_051_081, w_051_084, w_051_090, w_051_092, w_051_094, w_051_095, w_051_096, w_051_098, w_051_103, w_051_105, w_051_106, w_051_107, w_051_113, w_051_115, w_051_117, w_051_120, w_051_121, w_051_126, w_051_136, w_051_137, w_051_138, w_051_140, w_051_141, w_051_147, w_051_148, w_051_150, w_051_157, w_051_159, w_051_162, w_051_165, w_051_166, w_051_167, w_051_170, w_051_171, w_051_172, w_051_173, w_051_181, w_051_183, w_051_185, w_051_186, w_051_188, w_051_189, w_051_195, w_051_196, w_051_199, w_051_200, w_051_203, w_051_204, w_051_206, w_051_208, w_051_210, w_051_215, w_051_218, w_051_222, w_051_225, w_051_226, w_051_230, w_051_231, w_051_232, w_051_233, w_051_235, w_051_237, w_051_242, w_051_243, w_051_244, w_051_246, w_051_248, w_051_249, w_051_250, w_051_256, w_051_260, w_051_262, w_051_263, w_051_265, w_051_268, w_051_275, w_051_279, w_051_282, w_051_286, w_051_291, w_051_298, w_051_301, w_051_303, w_051_307, w_051_308, w_051_309, w_051_312, w_051_313, w_051_317, w_051_318, w_051_319, w_051_320, w_051_322, w_051_323, w_051_326, w_051_330, w_051_333, w_051_337, w_051_340, w_051_342, w_051_343, w_051_346, w_051_348, w_051_349, w_051_351, w_051_353, w_051_354, w_051_358, w_051_366, w_051_367, w_051_369, w_051_370, w_051_372, w_051_378, w_051_380, w_051_381, w_051_395, w_051_398, w_051_406;
  wire w_052_000, w_052_001, w_052_002, w_052_003, w_052_004, w_052_005, w_052_006, w_052_007, w_052_008, w_052_009, w_052_011, w_052_012, w_052_013, w_052_014, w_052_015, w_052_017, w_052_018, w_052_019, w_052_020, w_052_021, w_052_022, w_052_023, w_052_024, w_052_025, w_052_026, w_052_027, w_052_028, w_052_029, w_052_030, w_052_031, w_052_032, w_052_033, w_052_034, w_052_035, w_052_036, w_052_037, w_052_038, w_052_039, w_052_040, w_052_041, w_052_042, w_052_043, w_052_044, w_052_045, w_052_046;
  wire w_053_000, w_053_001, w_053_004, w_053_005, w_053_006, w_053_007, w_053_009, w_053_010, w_053_013, w_053_014, w_053_015, w_053_017, w_053_018, w_053_020, w_053_021, w_053_023, w_053_024, w_053_025, w_053_026, w_053_028, w_053_029, w_053_031, w_053_033, w_053_034, w_053_035, w_053_037, w_053_038, w_053_040, w_053_041, w_053_042, w_053_044, w_053_046, w_053_047, w_053_048, w_053_049, w_053_050, w_053_051, w_053_053, w_053_054, w_053_055, w_053_056, w_053_058, w_053_060, w_053_061, w_053_062, w_053_065, w_053_066, w_053_067, w_053_069, w_053_070, w_053_071, w_053_072, w_053_073, w_053_074, w_053_075, w_053_076, w_053_077, w_053_078, w_053_079, w_053_080, w_053_081, w_053_082, w_053_083, w_053_085, w_053_086, w_053_087, w_053_088, w_053_089, w_053_090, w_053_091, w_053_092, w_053_093, w_053_094, w_053_095, w_053_096, w_053_097, w_053_098, w_053_099, w_053_101, w_053_102, w_053_103, w_053_105, w_053_106, w_053_108, w_053_109, w_053_110, w_053_111, w_053_112, w_053_113, w_053_114, w_053_115, w_053_116, w_053_119, w_053_120, w_053_126, w_053_129, w_053_131, w_053_132, w_053_134, w_053_135, w_053_136, w_053_137, w_053_139, w_053_140, w_053_143, w_053_144, w_053_149, w_053_151, w_053_152, w_053_153, w_053_154, w_053_155, w_053_156, w_053_158, w_053_161;
  wire w_054_001, w_054_003, w_054_004, w_054_009, w_054_013, w_054_020, w_054_021, w_054_024, w_054_026, w_054_029, w_054_033, w_054_035, w_054_041, w_054_043, w_054_049, w_054_051, w_054_055, w_054_058, w_054_061, w_054_066, w_054_068, w_054_071, w_054_073, w_054_074, w_054_077, w_054_078, w_054_081, w_054_082, w_054_084, w_054_085, w_054_088, w_054_089, w_054_095, w_054_096, w_054_098, w_054_102, w_054_104, w_054_106, w_054_109, w_054_114, w_054_116, w_054_122, w_054_126, w_054_131, w_054_133, w_054_137, w_054_138, w_054_141, w_054_144, w_054_145, w_054_146, w_054_148, w_054_149, w_054_150, w_054_151, w_054_155, w_054_157, w_054_161, w_054_162, w_054_164, w_054_166, w_054_167, w_054_169, w_054_170, w_054_173, w_054_176, w_054_178, w_054_184, w_054_186, w_054_190, w_054_194, w_054_199, w_054_203, w_054_214, w_054_228, w_054_230, w_054_231, w_054_234, w_054_239, w_054_240, w_054_252, w_054_256, w_054_258, w_054_262, w_054_274, w_054_276, w_054_279, w_054_283, w_054_284, w_054_305, w_054_310, w_054_314, w_054_319, w_054_323, w_054_332, w_054_344, w_054_346, w_054_347, w_054_365, w_054_394, w_054_410, w_054_412, w_054_415, w_054_417, w_054_425, w_054_431, w_054_439, w_054_440, w_054_456, w_054_463, w_054_466, w_054_467, w_054_472, w_054_486, w_054_490, w_054_494, w_054_502, w_054_508, w_054_510, w_054_515, w_054_521, w_054_533, w_054_534, w_054_542, w_054_545, w_054_549, w_054_557, w_054_569, w_054_581, w_054_588, w_054_590;
  wire w_055_000, w_055_006, w_055_007, w_055_014, w_055_015, w_055_018, w_055_022, w_055_023, w_055_027, w_055_029, w_055_030, w_055_033, w_055_034, w_055_035, w_055_036, w_055_038, w_055_039, w_055_040, w_055_041, w_055_042, w_055_043, w_055_045, w_055_046, w_055_047, w_055_049, w_055_051, w_055_052, w_055_053, w_055_057, w_055_058, w_055_059, w_055_061, w_055_064, w_055_066, w_055_068, w_055_072, w_055_074, w_055_076, w_055_077, w_055_078, w_055_080, w_055_082, w_055_084, w_055_085, w_055_088, w_055_089, w_055_090, w_055_091, w_055_094, w_055_095, w_055_096, w_055_097, w_055_103, w_055_104, w_055_106, w_055_108, w_055_110, w_055_114, w_055_116, w_055_122, w_055_123, w_055_124, w_055_127, w_055_129, w_055_131, w_055_132, w_055_133, w_055_137, w_055_138, w_055_139, w_055_140, w_055_142, w_055_145, w_055_154, w_055_155, w_055_156, w_055_161, w_055_164, w_055_165, w_055_168, w_055_174, w_055_180, w_055_181, w_055_183, w_055_185, w_055_187, w_055_191, w_055_192, w_055_197, w_055_200, w_055_202, w_055_204, w_055_207, w_055_213, w_055_215, w_055_219, w_055_220, w_055_225, w_055_226, w_055_227, w_055_234, w_055_236, w_055_239, w_055_240, w_055_241, w_055_242, w_055_243, w_055_254, w_055_255, w_055_257, w_055_258, w_055_259, w_055_262, w_055_265, w_055_266, w_055_267, w_055_276, w_055_279, w_055_282, w_055_285, w_055_286, w_055_287, w_055_290, w_055_294, w_055_297, w_055_298, w_055_302, w_055_307, w_055_309, w_055_312, w_055_313, w_055_316, w_055_324, w_055_330, w_055_337, w_055_339, w_055_344, w_055_345;
  wire w_056_007, w_056_008, w_056_009, w_056_012, w_056_016, w_056_017, w_056_020, w_056_022, w_056_030, w_056_033, w_056_035, w_056_037, w_056_038, w_056_039, w_056_044, w_056_046, w_056_048, w_056_049, w_056_051, w_056_057, w_056_058, w_056_069, w_056_070, w_056_071, w_056_081, w_056_082, w_056_084, w_056_088, w_056_089, w_056_090, w_056_094, w_056_106, w_056_108, w_056_119, w_056_120, w_056_123, w_056_129, w_056_141, w_056_145, w_056_154, w_056_172, w_056_176, w_056_184, w_056_200, w_056_214, w_056_224, w_056_229, w_056_231, w_056_232, w_056_235, w_056_238, w_056_241, w_056_242, w_056_244, w_056_249, w_056_250, w_056_252, w_056_254, w_056_255, w_056_267, w_056_280, w_056_289, w_056_303, w_056_314, w_056_317, w_056_323, w_056_332, w_056_348, w_056_357, w_056_365, w_056_369, w_056_371, w_056_383, w_056_390, w_056_400, w_056_412, w_056_427, w_056_434, w_056_438, w_056_457, w_056_462, w_056_463, w_056_465, w_056_466, w_056_476, w_056_487, w_056_490, w_056_491, w_056_493, w_056_499, w_056_500, w_056_501, w_056_505, w_056_507, w_056_509, w_056_520, w_056_523, w_056_525, w_056_528, w_056_532, w_056_540, w_056_545, w_056_551, w_056_554, w_056_557, w_056_567, w_056_579, w_056_586, w_056_596, w_056_597, w_056_609, w_056_610, w_056_615, w_056_620, w_056_622, w_056_623, w_056_627, w_056_629, w_056_633, w_056_642, w_056_645, w_056_655, w_056_661, w_056_663, w_056_665, w_056_675, w_056_686, w_056_692, w_056_702, w_056_703, w_056_709, w_056_710, w_056_713, w_056_721, w_056_723, w_056_724, w_056_736;
  wire w_057_000, w_057_001, w_057_002, w_057_004, w_057_006, w_057_007, w_057_008, w_057_010, w_057_013, w_057_018, w_057_019, w_057_022, w_057_023, w_057_025, w_057_028, w_057_029, w_057_032, w_057_036, w_057_047, w_057_049, w_057_052, w_057_053, w_057_055, w_057_056, w_057_057, w_057_058, w_057_060, w_057_061, w_057_062, w_057_063, w_057_066, w_057_068, w_057_070, w_057_073, w_057_076, w_057_078, w_057_081, w_057_082, w_057_083, w_057_084, w_057_085, w_057_086, w_057_087, w_057_088, w_057_092, w_057_094, w_057_095, w_057_097, w_057_099, w_057_100, w_057_101, w_057_102, w_057_105, w_057_107, w_057_112, w_057_114, w_057_117, w_057_121, w_057_123, w_057_124, w_057_126, w_057_131, w_057_135, w_057_137, w_057_140, w_057_141, w_057_143, w_057_144, w_057_145, w_057_146, w_057_147, w_057_150, w_057_155, w_057_156, w_057_160, w_057_171, w_057_174, w_057_175, w_057_182, w_057_185, w_057_187, w_057_194, w_057_200, w_057_203, w_057_210, w_057_213, w_057_215, w_057_220, w_057_228, w_057_229, w_057_230, w_057_235, w_057_236, w_057_237, w_057_239, w_057_241, w_057_243, w_057_246, w_057_250, w_057_254, w_057_257, w_057_258, w_057_262, w_057_268, w_057_271, w_057_273, w_057_274, w_057_279, w_057_281, w_057_285, w_057_289, w_057_291, w_057_293, w_057_296, w_057_307, w_057_313;
  wire w_058_005, w_058_017, w_058_022, w_058_025, w_058_029, w_058_030, w_058_032, w_058_033, w_058_037, w_058_050, w_058_056, w_058_060, w_058_061, w_058_065, w_058_070, w_058_073, w_058_074, w_058_075, w_058_081, w_058_082, w_058_085, w_058_086, w_058_088, w_058_090, w_058_092, w_058_095, w_058_104, w_058_105, w_058_111, w_058_112, w_058_119, w_058_123, w_058_132, w_058_134, w_058_135, w_058_136, w_058_140, w_058_148, w_058_156, w_058_159, w_058_161, w_058_162, w_058_164, w_058_171, w_058_174, w_058_179, w_058_182, w_058_193, w_058_195, w_058_206, w_058_208, w_058_210, w_058_216, w_058_224, w_058_229, w_058_235, w_058_238, w_058_251, w_058_253, w_058_254, w_058_255, w_058_256, w_058_258, w_058_271, w_058_274, w_058_280, w_058_282, w_058_287, w_058_292, w_058_295, w_058_304, w_058_306, w_058_310, w_058_316, w_058_321, w_058_327, w_058_330, w_058_332, w_058_335, w_058_341, w_058_344, w_058_352, w_058_359, w_058_366, w_058_368, w_058_376, w_058_379, w_058_383, w_058_402, w_058_404, w_058_416, w_058_420, w_058_423, w_058_425, w_058_427, w_058_428, w_058_442, w_058_447, w_058_453, w_058_454, w_058_457, w_058_459, w_058_467, w_058_469, w_058_472, w_058_477, w_058_478, w_058_479, w_058_484, w_058_485, w_058_493, w_058_498, w_058_503, w_058_504, w_058_505, w_058_513, w_058_515, w_058_522, w_058_527, w_058_534, w_058_536, w_058_538, w_058_540, w_058_541, w_058_550, w_058_555, w_058_559, w_058_562, w_058_568, w_058_570, w_058_581, w_058_589, w_058_590, w_058_593, w_058_594, w_058_596, w_058_597, w_058_602, w_058_607, w_058_635, w_058_638, w_058_645, w_058_647, w_058_655, w_058_656, w_058_658, w_058_660, w_058_664, w_058_673, w_058_681, w_058_683, w_058_696, w_058_699;
  wire w_059_001, w_059_002, w_059_003, w_059_005, w_059_012, w_059_017, w_059_026, w_059_029, w_059_032, w_059_043, w_059_045, w_059_049, w_059_052, w_059_055, w_059_056, w_059_057, w_059_060, w_059_061, w_059_066, w_059_084, w_059_089, w_059_090, w_059_094, w_059_101, w_059_103, w_059_111, w_059_114, w_059_125, w_059_131, w_059_135, w_059_140, w_059_146, w_059_147, w_059_150, w_059_157, w_059_159, w_059_162, w_059_165, w_059_166, w_059_167, w_059_168, w_059_170, w_059_173, w_059_174, w_059_178, w_059_181, w_059_183, w_059_184, w_059_186, w_059_196, w_059_200, w_059_201, w_059_202, w_059_209, w_059_213, w_059_218, w_059_220, w_059_233, w_059_236, w_059_239, w_059_242, w_059_248, w_059_249, w_059_255, w_059_258, w_059_260, w_059_278, w_059_286, w_059_288, w_059_301, w_059_309, w_059_313, w_059_315, w_059_321, w_059_328, w_059_337, w_059_340, w_059_348, w_059_354, w_059_355, w_059_364, w_059_392, w_059_396, w_059_405, w_059_413, w_059_423, w_059_425, w_059_430, w_059_431, w_059_432, w_059_439, w_059_444, w_059_455, w_059_459, w_059_462, w_059_479, w_059_482, w_059_489, w_059_500, w_059_501, w_059_507, w_059_508, w_059_512, w_059_517, w_059_521, w_059_522, w_059_533, w_059_538, w_059_550, w_059_552, w_059_553, w_059_554, w_059_555, w_059_559, w_059_567, w_059_578, w_059_587, w_059_588, w_059_589, w_059_596, w_059_600, w_059_612, w_059_616, w_059_633, w_059_636, w_059_637, w_059_639, w_059_647, w_059_660, w_059_667, w_059_683, w_059_695, w_059_698, w_059_702, w_059_708, w_059_722, w_059_724, w_059_727, w_059_730, w_059_734;
  wire w_060_003, w_060_009, w_060_012, w_060_016, w_060_017, w_060_019, w_060_020, w_060_024, w_060_025, w_060_026, w_060_027, w_060_030, w_060_033, w_060_036, w_060_037, w_060_038, w_060_039, w_060_045, w_060_049, w_060_050, w_060_053, w_060_058, w_060_071, w_060_073, w_060_075, w_060_080, w_060_081, w_060_085, w_060_086, w_060_088, w_060_097, w_060_098, w_060_109, w_060_112, w_060_114, w_060_116, w_060_118, w_060_119, w_060_122, w_060_123, w_060_125, w_060_126, w_060_131, w_060_141, w_060_148, w_060_155, w_060_160, w_060_161, w_060_164, w_060_167, w_060_168, w_060_169, w_060_171, w_060_176, w_060_189, w_060_190, w_060_194, w_060_198, w_060_204, w_060_208, w_060_209, w_060_212, w_060_216, w_060_222, w_060_224, w_060_225, w_060_246, w_060_254, w_060_257, w_060_259, w_060_261, w_060_262, w_060_265, w_060_266, w_060_268, w_060_272, w_060_277, w_060_278, w_060_284, w_060_285, w_060_288, w_060_289, w_060_290, w_060_291, w_060_294, w_060_296, w_060_299, w_060_300, w_060_305, w_060_308, w_060_310, w_060_313, w_060_323, w_060_324, w_060_326, w_060_330, w_060_331, w_060_332, w_060_333, w_060_336, w_060_338, w_060_341, w_060_343, w_060_344, w_060_354, w_060_355, w_060_359, w_060_365, w_060_366, w_060_372, w_060_381, w_060_387, w_060_395;
  wire w_061_002, w_061_003, w_061_004, w_061_005, w_061_012, w_061_023, w_061_027, w_061_028, w_061_029, w_061_033, w_061_042, w_061_046, w_061_047, w_061_050, w_061_051, w_061_052, w_061_056, w_061_057, w_061_058, w_061_059, w_061_061, w_061_062, w_061_063, w_061_064, w_061_065, w_061_066, w_061_073, w_061_082, w_061_084, w_061_088, w_061_089, w_061_099, w_061_100, w_061_101, w_061_103, w_061_105, w_061_106, w_061_122, w_061_123, w_061_125, w_061_126, w_061_142, w_061_143, w_061_146, w_061_147, w_061_148, w_061_157, w_061_158, w_061_160, w_061_161, w_061_162, w_061_168, w_061_172, w_061_175, w_061_178, w_061_179, w_061_182, w_061_184, w_061_188, w_061_192, w_061_194, w_061_196, w_061_198, w_061_199, w_061_200, w_061_205, w_061_213, w_061_217, w_061_219, w_061_221, w_061_227, w_061_230, w_061_240, w_061_241, w_061_242, w_061_253, w_061_255, w_061_256, w_061_257, w_061_260, w_061_264, w_061_266, w_061_270, w_061_271, w_061_276, w_061_277, w_061_283, w_061_285, w_061_287, w_061_294, w_061_296, w_061_298, w_061_300, w_061_301, w_061_302, w_061_305, w_061_306, w_061_307, w_061_311, w_061_313, w_061_314, w_061_323, w_061_326, w_061_338, w_061_343, w_061_356, w_061_357, w_061_365, w_061_374, w_061_380, w_061_383, w_061_388, w_061_405, w_061_407, w_061_408, w_061_426, w_061_434, w_061_437, w_061_440, w_061_443, w_061_452, w_061_464, w_061_465, w_061_467, w_061_472, w_061_473, w_061_477, w_061_486, w_061_487, w_061_488, w_061_489;
  wire w_062_000, w_062_003, w_062_009, w_062_013, w_062_017, w_062_027, w_062_030, w_062_057, w_062_058, w_062_060, w_062_081, w_062_083, w_062_088, w_062_089, w_062_093, w_062_096, w_062_099, w_062_100, w_062_116, w_062_125, w_062_128, w_062_131, w_062_132, w_062_134, w_062_135, w_062_138, w_062_140, w_062_144, w_062_149, w_062_151, w_062_157, w_062_159, w_062_162, w_062_164, w_062_168, w_062_173, w_062_177, w_062_178, w_062_185, w_062_194, w_062_206, w_062_208, w_062_211, w_062_220, w_062_224, w_062_229, w_062_239, w_062_241, w_062_245, w_062_249, w_062_250, w_062_251, w_062_253, w_062_259, w_062_264, w_062_268, w_062_273, w_062_280, w_062_282, w_062_305, w_062_307, w_062_308, w_062_311, w_062_313, w_062_316, w_062_329, w_062_330, w_062_338, w_062_342, w_062_349, w_062_352, w_062_355, w_062_362, w_062_370, w_062_371, w_062_377, w_062_378, w_062_380, w_062_384, w_062_390, w_062_401, w_062_406, w_062_430, w_062_435, w_062_440, w_062_455, w_062_458, w_062_465, w_062_473, w_062_483, w_062_484, w_062_503, w_062_508, w_062_511, w_062_512, w_062_513, w_062_516, w_062_517, w_062_518, w_062_526, w_062_535, w_062_539, w_062_540, w_062_544, w_062_546, w_062_549, w_062_554, w_062_586, w_062_591, w_062_593, w_062_598, w_062_606, w_062_607, w_062_612, w_062_628, w_062_633, w_062_643, w_062_653, w_062_661, w_062_666, w_062_670, w_062_672, w_062_673, w_062_677, w_062_689, w_062_696, w_062_697, w_062_704, w_062_718, w_062_731, w_062_732, w_062_734, w_062_739, w_062_745, w_062_761, w_062_768, w_062_772, w_062_776, w_062_784, w_062_785, w_062_796;
  wire w_063_002, w_063_003, w_063_004, w_063_005, w_063_006, w_063_008, w_063_009, w_063_010, w_063_014, w_063_018, w_063_019, w_063_024, w_063_025, w_063_026, w_063_027, w_063_029, w_063_034, w_063_035, w_063_036, w_063_045, w_063_047, w_063_050, w_063_052, w_063_058, w_063_059, w_063_062, w_063_063, w_063_064, w_063_066, w_063_072, w_063_073, w_063_076, w_063_082, w_063_083, w_063_084, w_063_085, w_063_086, w_063_088, w_063_089, w_063_090, w_063_093, w_063_094, w_063_101, w_063_104, w_063_107, w_063_108, w_063_109, w_063_110, w_063_111, w_063_113, w_063_114, w_063_115, w_063_120, w_063_121, w_063_123, w_063_128, w_063_133, w_063_139, w_063_142, w_063_149, w_063_153, w_063_155, w_063_156, w_063_160, w_063_166, w_063_173, w_063_175, w_063_176, w_063_177, w_063_178, w_063_179, w_063_180, w_063_181, w_063_183, w_063_188, w_063_190, w_063_193, w_063_194, w_063_197, w_063_198, w_063_208, w_063_212, w_063_213, w_063_216, w_063_218, w_063_219, w_063_222, w_063_223, w_063_224, w_063_225, w_063_226, w_063_227, w_063_228, w_063_229, w_063_233, w_063_238, w_063_244, w_063_245, w_063_250, w_063_251, w_063_252, w_063_262, w_063_267, w_063_268, w_063_269, w_063_274, w_063_290, w_063_297, w_063_301, w_063_302, w_063_304, w_063_317, w_063_319, w_063_326, w_063_341, w_063_361, w_063_366, w_063_374, w_063_376, w_063_383, w_063_387, w_063_388, w_063_397, w_063_400, w_063_402, w_063_410, w_063_415, w_063_417, w_063_418, w_063_421, w_063_424, w_063_432, w_063_438, w_063_445, w_063_450, w_063_456, w_063_469, w_063_470, w_063_483, w_063_503, w_063_504, w_063_509, w_063_514, w_063_519, w_063_524, w_063_527, w_063_528, w_063_545, w_063_547;
  wire w_064_004, w_064_005, w_064_009, w_064_010, w_064_012, w_064_014, w_064_018, w_064_020, w_064_027, w_064_029, w_064_032, w_064_034, w_064_036, w_064_038, w_064_044, w_064_049, w_064_052, w_064_055, w_064_056, w_064_058, w_064_059, w_064_061, w_064_064, w_064_066, w_064_069, w_064_070, w_064_072, w_064_074, w_064_077, w_064_078, w_064_080, w_064_081, w_064_082, w_064_086, w_064_087, w_064_093, w_064_094, w_064_097, w_064_100, w_064_103, w_064_106, w_064_107, w_064_111, w_064_112, w_064_114, w_064_115, w_064_118, w_064_121, w_064_125, w_064_127, w_064_130, w_064_133, w_064_134, w_064_135, w_064_136, w_064_140, w_064_142, w_064_143, w_064_150, w_064_153, w_064_154, w_064_155, w_064_165, w_064_166, w_064_170, w_064_174, w_064_180, w_064_182, w_064_184, w_064_194, w_064_197, w_064_202, w_064_205, w_064_207, w_064_214, w_064_215, w_064_226, w_064_228, w_064_229, w_064_233, w_064_235, w_064_237, w_064_241, w_064_253, w_064_255, w_064_256, w_064_265, w_064_267, w_064_271, w_064_279, w_064_280, w_064_285, w_064_286, w_064_289, w_064_297, w_064_306, w_064_308, w_064_310, w_064_311, w_064_312, w_064_315, w_064_324, w_064_327, w_064_328, w_064_329, w_064_330, w_064_335, w_064_338, w_064_339, w_064_345;
  wire w_065_000, w_065_010, w_065_012, w_065_015, w_065_016, w_065_026, w_065_028, w_065_031, w_065_032, w_065_038, w_065_040, w_065_043, w_065_046, w_065_056, w_065_058, w_065_059, w_065_060, w_065_063, w_065_066, w_065_069, w_065_074, w_065_075, w_065_084, w_065_086, w_065_087, w_065_095, w_065_097, w_065_098, w_065_107, w_065_117, w_065_126, w_065_132, w_065_136, w_065_144, w_065_152, w_065_165, w_065_172, w_065_174, w_065_181, w_065_185, w_065_214, w_065_218, w_065_228, w_065_244, w_065_246, w_065_248, w_065_250, w_065_253, w_065_256, w_065_259, w_065_263, w_065_270, w_065_272, w_065_275, w_065_280, w_065_285, w_065_295, w_065_296, w_065_304, w_065_307, w_065_311, w_065_316, w_065_320, w_065_327, w_065_333, w_065_338, w_065_342, w_065_343, w_065_344, w_065_348, w_065_359, w_065_361, w_065_363, w_065_372, w_065_381, w_065_386, w_065_387, w_065_389, w_065_393, w_065_407, w_065_411, w_065_425, w_065_426, w_065_449, w_065_453, w_065_474, w_065_496, w_065_499, w_065_507, w_065_512, w_065_515, w_065_517, w_065_522, w_065_537, w_065_542, w_065_543, w_065_547, w_065_555, w_065_557, w_065_558, w_065_563, w_065_565, w_065_569, w_065_572, w_065_576, w_065_582, w_065_590, w_065_593, w_065_603, w_065_606, w_065_609, w_065_641, w_065_646, w_065_654, w_065_658, w_065_666, w_065_668, w_065_673, w_065_687;
  wire w_066_004, w_066_007, w_066_011, w_066_013, w_066_017, w_066_023, w_066_025, w_066_029, w_066_035, w_066_040, w_066_045, w_066_052, w_066_058, w_066_061, w_066_063, w_066_064, w_066_072, w_066_080, w_066_084, w_066_089, w_066_093, w_066_095, w_066_099, w_066_101, w_066_103, w_066_104, w_066_110, w_066_111, w_066_112, w_066_115, w_066_118, w_066_119, w_066_123, w_066_125, w_066_126, w_066_134, w_066_135, w_066_141, w_066_147, w_066_154, w_066_170, w_066_181, w_066_182, w_066_185, w_066_191, w_066_202, w_066_216, w_066_224, w_066_234, w_066_240, w_066_243, w_066_246, w_066_273, w_066_276, w_066_281, w_066_290, w_066_293, w_066_315, w_066_319, w_066_327, w_066_335, w_066_341, w_066_343, w_066_348, w_066_349, w_066_356, w_066_370, w_066_372, w_066_376, w_066_378, w_066_385, w_066_402, w_066_403, w_066_404, w_066_405, w_066_406, w_066_416, w_066_421, w_066_433, w_066_454, w_066_463, w_066_473, w_066_476, w_066_482, w_066_489, w_066_493, w_066_503, w_066_512, w_066_516, w_066_518, w_066_531, w_066_542, w_066_544, w_066_555, w_066_556, w_066_558, w_066_559, w_066_572, w_066_578, w_066_584, w_066_586, w_066_594, w_066_595, w_066_625, w_066_627;
  wire w_067_003, w_067_005, w_067_007, w_067_010, w_067_013, w_067_020, w_067_021, w_067_024, w_067_027, w_067_037, w_067_039, w_067_046, w_067_049, w_067_052, w_067_053, w_067_060, w_067_062, w_067_069, w_067_076, w_067_083, w_067_094, w_067_099, w_067_101, w_067_104, w_067_111, w_067_113, w_067_119, w_067_122, w_067_125, w_067_126, w_067_133, w_067_134, w_067_137, w_067_140, w_067_141, w_067_146, w_067_150, w_067_154, w_067_156, w_067_162, w_067_163, w_067_165, w_067_166, w_067_169, w_067_171, w_067_175, w_067_196, w_067_199, w_067_201, w_067_204, w_067_206, w_067_211, w_067_213, w_067_224, w_067_232, w_067_239, w_067_250, w_067_253, w_067_254, w_067_255, w_067_263, w_067_266, w_067_270, w_067_273, w_067_275, w_067_276, w_067_280, w_067_290, w_067_292, w_067_297, w_067_302, w_067_305, w_067_316, w_067_318, w_067_326, w_067_328, w_067_329, w_067_333, w_067_334, w_067_336, w_067_342, w_067_343, w_067_344, w_067_346, w_067_347, w_067_352, w_067_353, w_067_356, w_067_358, w_067_360, w_067_362, w_067_363, w_067_371, w_067_373, w_067_374, w_067_381, w_067_382, w_067_383, w_067_390, w_067_395;
  wire w_068_000, w_068_001, w_068_008, w_068_009, w_068_011, w_068_012, w_068_024, w_068_030, w_068_041, w_068_042, w_068_052, w_068_056, w_068_060, w_068_062, w_068_069, w_068_070, w_068_074, w_068_075, w_068_076, w_068_079, w_068_080, w_068_081, w_068_082, w_068_083, w_068_084, w_068_086, w_068_092, w_068_094, w_068_095, w_068_098, w_068_101, w_068_102, w_068_106, w_068_113, w_068_114, w_068_124, w_068_125, w_068_131, w_068_133, w_068_136, w_068_138, w_068_139, w_068_153, w_068_167, w_068_170, w_068_174, w_068_176, w_068_181, w_068_182, w_068_183, w_068_192, w_068_194, w_068_200, w_068_204, w_068_206, w_068_209, w_068_210, w_068_213, w_068_221, w_068_224, w_068_225, w_068_226, w_068_231, w_068_237, w_068_242, w_068_246, w_068_249, w_068_250, w_068_260, w_068_265, w_068_267, w_068_268, w_068_275, w_068_276, w_068_280, w_068_283, w_068_295, w_068_298, w_068_301, w_068_304, w_068_306, w_068_307, w_068_308, w_068_309, w_068_321, w_068_322, w_068_323, w_068_328, w_068_334, w_068_337, w_068_340, w_068_342, w_068_344, w_068_346, w_068_348, w_068_349, w_068_352, w_068_357, w_068_360, w_068_361;
  wire w_069_001, w_069_003, w_069_005, w_069_009, w_069_014, w_069_016, w_069_022, w_069_023, w_069_025, w_069_028, w_069_029, w_069_033, w_069_034, w_069_038, w_069_039, w_069_042, w_069_048, w_069_049, w_069_053, w_069_055, w_069_060, w_069_063, w_069_064, w_069_065, w_069_067, w_069_068, w_069_071, w_069_075, w_069_076, w_069_077, w_069_078, w_069_080, w_069_081, w_069_087, w_069_088, w_069_089, w_069_091, w_069_093, w_069_096, w_069_097, w_069_104, w_069_105, w_069_107, w_069_110, w_069_117, w_069_120, w_069_125, w_069_128, w_069_140, w_069_141, w_069_143, w_069_144, w_069_145, w_069_146, w_069_153, w_069_157, w_069_158, w_069_159, w_069_165, w_069_167, w_069_168, w_069_171, w_069_173, w_069_174, w_069_176, w_069_177, w_069_181, w_069_182, w_069_185, w_069_188, w_069_191, w_069_192, w_069_194, w_069_197, w_069_199, w_069_202, w_069_207, w_069_209, w_069_213, w_069_218, w_069_223, w_069_225, w_069_226, w_069_227, w_069_228, w_069_230, w_069_232, w_069_236, w_069_237, w_069_241, w_069_242, w_069_245, w_069_254, w_069_259, w_069_260, w_069_265;
  wire w_070_000, w_070_004, w_070_006, w_070_007, w_070_008, w_070_009, w_070_010, w_070_014, w_070_018, w_070_019, w_070_021, w_070_027, w_070_028, w_070_031, w_070_033, w_070_035, w_070_041, w_070_044, w_070_050, w_070_056, w_070_060, w_070_069, w_070_071, w_070_080, w_070_083, w_070_084, w_070_089, w_070_096, w_070_100, w_070_104, w_070_108, w_070_109, w_070_112, w_070_117, w_070_121, w_070_123, w_070_142, w_070_143, w_070_148, w_070_155, w_070_158, w_070_161, w_070_170, w_070_173, w_070_174, w_070_175, w_070_179, w_070_185, w_070_190, w_070_191, w_070_192, w_070_199, w_070_205, w_070_209, w_070_210, w_070_213, w_070_216, w_070_220, w_070_232, w_070_253, w_070_256, w_070_270, w_070_271, w_070_280, w_070_287, w_070_289, w_070_292, w_070_293, w_070_294, w_070_325, w_070_327, w_070_329, w_070_330, w_070_359, w_070_365, w_070_381, w_070_384, w_070_386, w_070_389, w_070_390, w_070_396, w_070_404, w_070_408, w_070_412, w_070_424, w_070_435, w_070_437, w_070_444, w_070_453, w_070_455, w_070_459, w_070_465, w_070_468, w_070_471, w_070_473, w_070_476, w_070_478, w_070_480, w_070_482, w_070_486, w_070_488, w_070_489, w_070_496, w_070_499, w_070_505, w_070_508, w_070_510, w_070_515, w_070_530, w_070_542, w_070_548, w_070_563, w_070_568, w_070_572, w_070_573, w_070_579;
  wire w_071_000, w_071_001, w_071_014, w_071_018, w_071_020, w_071_022, w_071_026, w_071_029, w_071_031, w_071_034, w_071_038, w_071_045, w_071_047, w_071_048, w_071_052, w_071_055, w_071_056, w_071_058, w_071_063, w_071_066, w_071_075, w_071_076, w_071_082, w_071_084, w_071_085, w_071_091, w_071_093, w_071_094, w_071_095, w_071_096, w_071_097, w_071_099, w_071_100, w_071_102, w_071_104, w_071_105, w_071_107, w_071_109, w_071_113, w_071_121, w_071_124, w_071_129, w_071_138, w_071_143, w_071_144, w_071_145, w_071_147, w_071_148, w_071_151, w_071_154, w_071_155, w_071_171, w_071_173, w_071_176, w_071_188, w_071_205, w_071_206, w_071_209, w_071_213, w_071_217, w_071_227, w_071_247, w_071_250, w_071_252, w_071_257, w_071_260, w_071_261, w_071_265, w_071_267, w_071_270, w_071_276, w_071_277, w_071_281, w_071_284, w_071_289, w_071_294, w_071_299, w_071_300, w_071_302, w_071_303, w_071_304, w_071_305, w_071_312, w_071_315, w_071_316, w_071_317, w_071_322;
  wire w_072_000, w_072_001, w_072_003, w_072_005, w_072_012, w_072_017, w_072_020, w_072_021, w_072_024, w_072_034, w_072_043, w_072_047, w_072_048, w_072_051, w_072_052, w_072_053, w_072_054, w_072_057, w_072_058, w_072_059, w_072_060, w_072_061, w_072_064, w_072_067, w_072_070, w_072_082, w_072_084, w_072_090, w_072_092, w_072_095, w_072_096, w_072_097, w_072_098, w_072_101, w_072_102, w_072_103, w_072_106, w_072_107, w_072_111, w_072_113, w_072_114, w_072_116, w_072_120, w_072_122, w_072_123, w_072_129, w_072_130, w_072_131, w_072_134, w_072_135, w_072_137, w_072_143, w_072_144, w_072_149, w_072_152, w_072_156, w_072_157, w_072_161, w_072_163, w_072_165, w_072_167, w_072_169, w_072_171, w_072_172, w_072_175, w_072_177, w_072_178, w_072_184, w_072_186, w_072_187, w_072_190, w_072_195, w_072_199, w_072_201, w_072_208, w_072_215, w_072_232, w_072_235, w_072_242, w_072_260, w_072_266, w_072_272, w_072_278, w_072_288, w_072_289, w_072_292, w_072_295;
  wire w_073_000, w_073_003, w_073_009, w_073_016, w_073_017, w_073_018, w_073_020, w_073_026, w_073_034, w_073_037, w_073_040, w_073_041, w_073_042, w_073_043, w_073_044, w_073_049, w_073_052, w_073_053, w_073_055, w_073_068, w_073_071, w_073_085, w_073_088, w_073_090, w_073_095, w_073_101, w_073_114, w_073_117, w_073_130, w_073_139, w_073_143, w_073_150, w_073_169, w_073_175, w_073_183, w_073_196, w_073_198, w_073_200, w_073_203, w_073_204, w_073_209, w_073_219, w_073_224, w_073_245, w_073_252, w_073_253, w_073_258, w_073_262, w_073_284, w_073_299, w_073_326, w_073_347, w_073_363, w_073_374, w_073_379, w_073_382, w_073_402, w_073_404, w_073_407, w_073_413, w_073_419, w_073_422, w_073_428, w_073_439, w_073_443, w_073_457, w_073_463, w_073_474, w_073_484, w_073_489, w_073_492, w_073_493, w_073_499, w_073_503, w_073_507, w_073_512, w_073_514, w_073_516, w_073_526, w_073_537, w_073_540, w_073_554, w_073_569, w_073_592, w_073_601, w_073_602, w_073_605, w_073_613, w_073_621, w_073_624, w_073_627, w_073_632, w_073_634, w_073_649, w_073_675, w_073_687, w_073_688, w_073_691, w_073_697, w_073_714, w_073_715, w_073_717, w_073_722, w_073_734, w_073_735, w_073_740;
  wire w_074_000, w_074_005, w_074_009, w_074_012, w_074_014, w_074_023, w_074_024, w_074_030, w_074_032, w_074_033, w_074_041, w_074_044, w_074_045, w_074_046, w_074_052, w_074_070, w_074_077, w_074_081, w_074_099, w_074_100, w_074_104, w_074_105, w_074_107, w_074_108, w_074_111, w_074_114, w_074_117, w_074_124, w_074_127, w_074_128, w_074_141, w_074_144, w_074_152, w_074_153, w_074_154, w_074_157, w_074_159, w_074_166, w_074_168, w_074_169, w_074_175, w_074_176, w_074_177, w_074_179, w_074_182, w_074_184, w_074_186, w_074_190, w_074_193, w_074_194, w_074_196, w_074_200, w_074_201, w_074_209, w_074_210, w_074_215, w_074_218, w_074_221, w_074_227, w_074_231, w_074_232, w_074_233, w_074_243, w_074_250, w_074_251, w_074_252, w_074_254, w_074_256, w_074_258, w_074_259, w_074_265, w_074_277, w_074_287, w_074_288, w_074_293, w_074_294, w_074_296, w_074_297, w_074_300, w_074_303, w_074_309, w_074_313, w_074_317, w_074_320, w_074_321, w_074_322, w_074_327, w_074_331, w_074_334, w_074_337, w_074_340, w_074_342, w_074_343, w_074_344, w_074_345, w_074_348, w_074_351, w_074_360, w_074_363, w_074_370, w_074_374, w_074_375;
  wire w_075_000, w_075_001, w_075_002, w_075_005, w_075_007, w_075_009, w_075_010, w_075_011, w_075_013, w_075_014, w_075_016, w_075_018, w_075_019, w_075_020, w_075_023, w_075_024, w_075_025, w_075_027, w_075_030, w_075_032, w_075_033, w_075_034, w_075_037, w_075_039, w_075_043, w_075_044, w_075_045, w_075_046, w_075_047, w_075_049, w_075_050, w_075_052, w_075_053, w_075_054, w_075_055, w_075_058, w_075_061, w_075_062, w_075_063, w_075_065, w_075_067, w_075_069, w_075_071, w_075_072, w_075_074, w_075_076, w_075_077, w_075_078, w_075_079, w_075_083, w_075_087, w_075_091, w_075_096, w_075_097, w_075_100, w_075_101, w_075_105, w_075_109, w_075_111, w_075_113, w_075_114, w_075_116, w_075_117, w_075_118, w_075_120, w_075_127, w_075_128, w_075_132, w_075_133, w_075_134, w_075_135, w_075_136, w_075_137, w_075_138, w_075_139, w_075_140, w_075_141, w_075_144, w_075_145, w_075_147, w_075_148, w_075_152, w_075_153, w_075_155, w_075_158, w_075_159, w_075_160, w_075_161;
  wire w_076_014, w_076_015, w_076_033, w_076_036, w_076_040, w_076_043, w_076_046, w_076_050, w_076_052, w_076_060, w_076_062, w_076_070, w_076_072, w_076_074, w_076_087, w_076_091, w_076_098, w_076_099, w_076_102, w_076_104, w_076_107, w_076_108, w_076_111, w_076_115, w_076_130, w_076_134, w_076_136, w_076_137, w_076_140, w_076_145, w_076_157, w_076_158, w_076_161, w_076_162, w_076_168, w_076_173, w_076_181, w_076_182, w_076_183, w_076_197, w_076_200, w_076_201, w_076_206, w_076_209, w_076_210, w_076_218, w_076_220, w_076_221, w_076_233, w_076_237, w_076_240, w_076_241, w_076_255, w_076_258, w_076_262, w_076_277, w_076_292, w_076_294, w_076_295, w_076_296, w_076_300, w_076_311, w_076_319, w_076_321, w_076_326, w_076_327, w_076_334, w_076_345, w_076_347, w_076_351, w_076_362, w_076_364, w_076_375, w_076_405, w_076_418, w_076_421, w_076_432, w_076_447, w_076_458, w_076_459, w_076_461, w_076_476, w_076_479, w_076_489, w_076_493, w_076_494, w_076_495, w_076_496, w_076_497, w_076_498, w_076_499, w_076_500, w_076_501, w_076_502;
  wire w_077_000, w_077_011, w_077_019, w_077_021, w_077_022, w_077_026, w_077_029, w_077_032, w_077_035, w_077_039, w_077_043, w_077_044, w_077_048, w_077_052, w_077_054, w_077_057, w_077_058, w_077_060, w_077_086, w_077_089, w_077_091, w_077_099, w_077_102, w_077_107, w_077_110, w_077_123, w_077_127, w_077_133, w_077_140, w_077_150, w_077_151, w_077_152, w_077_165, w_077_166, w_077_176, w_077_178, w_077_185, w_077_209, w_077_210, w_077_223, w_077_232, w_077_240, w_077_242, w_077_245, w_077_251, w_077_254, w_077_262, w_077_272, w_077_282, w_077_286, w_077_289, w_077_290, w_077_292, w_077_310, w_077_313, w_077_315, w_077_321, w_077_344, w_077_361, w_077_372, w_077_378, w_077_382, w_077_385, w_077_398, w_077_401, w_077_409, w_077_412, w_077_420, w_077_424, w_077_431, w_077_440, w_077_444, w_077_479, w_077_481, w_077_483, w_077_488, w_077_500, w_077_519, w_077_522, w_077_540, w_077_551, w_077_552, w_077_558, w_077_560, w_077_577, w_077_586, w_077_590, w_077_592, w_077_597, w_077_601, w_077_610, w_077_619, w_077_626, w_077_630, w_077_631, w_077_632, w_077_633, w_077_634;
  wire w_078_004, w_078_013, w_078_015, w_078_016, w_078_024, w_078_033, w_078_037, w_078_038, w_078_039, w_078_043, w_078_044, w_078_050, w_078_053, w_078_055, w_078_056, w_078_058, w_078_061, w_078_063, w_078_070, w_078_078, w_078_080, w_078_083, w_078_084, w_078_089, w_078_093, w_078_101, w_078_102, w_078_103, w_078_104, w_078_106, w_078_112, w_078_121, w_078_122, w_078_130, w_078_142, w_078_144, w_078_145, w_078_149, w_078_150, w_078_152, w_078_166, w_078_168, w_078_169, w_078_170, w_078_177, w_078_183, w_078_188, w_078_195, w_078_200, w_078_208, w_078_213, w_078_225, w_078_229, w_078_230, w_078_251, w_078_306, w_078_318, w_078_329, w_078_345, w_078_349, w_078_366, w_078_379, w_078_381, w_078_396, w_078_401, w_078_416, w_078_421, w_078_428, w_078_429, w_078_434, w_078_441, w_078_445, w_078_446, w_078_464, w_078_465, w_078_475, w_078_497, w_078_511, w_078_514, w_078_520, w_078_560, w_078_566, w_078_571, w_078_573, w_078_588, w_078_597;
  wire w_079_000, w_079_001, w_079_002, w_079_003, w_079_004, w_079_005, w_079_007, w_079_008, w_079_010, w_079_012, w_079_015, w_079_016, w_079_017, w_079_018, w_079_020, w_079_021, w_079_022, w_079_023, w_079_024, w_079_025, w_079_027, w_079_028, w_079_029, w_079_030, w_079_031, w_079_033, w_079_035, w_079_036, w_079_037, w_079_038, w_079_039, w_079_040, w_079_041, w_079_043, w_079_044, w_079_045, w_079_047, w_079_048, w_079_050, w_079_051, w_079_052, w_079_053, w_079_054, w_079_055, w_079_056, w_079_057, w_079_058, w_079_059, w_079_060, w_079_062;
  wire w_080_003, w_080_007, w_080_011, w_080_013, w_080_019, w_080_023, w_080_029, w_080_032, w_080_033, w_080_044, w_080_052, w_080_053, w_080_054, w_080_063, w_080_065, w_080_076, w_080_079, w_080_080, w_080_085, w_080_086, w_080_096, w_080_098, w_080_113, w_080_118, w_080_120, w_080_131, w_080_132, w_080_134, w_080_138, w_080_153, w_080_154, w_080_158, w_080_159, w_080_162, w_080_171, w_080_173, w_080_176, w_080_182, w_080_183, w_080_185, w_080_186, w_080_192, w_080_202, w_080_212, w_080_213, w_080_222, w_080_225, w_080_230, w_080_231, w_080_233, w_080_237, w_080_238, w_080_245, w_080_249, w_080_251, w_080_255, w_080_257, w_080_269, w_080_279, w_080_284, w_080_287, w_080_289, w_080_290, w_080_295, w_080_303, w_080_311, w_080_313, w_080_319, w_080_336, w_080_360, w_080_362, w_080_369, w_080_389, w_080_394, w_080_397, w_080_399, w_080_403, w_080_407, w_080_417, w_080_430, w_080_433, w_080_440, w_080_464, w_080_472, w_080_476, w_080_477, w_080_478, w_080_481;
  wire w_081_000, w_081_001, w_081_002, w_081_003, w_081_004, w_081_005, w_081_006, w_081_007, w_081_008, w_081_009, w_081_010, w_081_011, w_081_012, w_081_013, w_081_014, w_081_015, w_081_016, w_081_017, w_081_018, w_081_019, w_081_020, w_081_021, w_081_022;
  wire w_082_003, w_082_019, w_082_020, w_082_026, w_082_027, w_082_040, w_082_041, w_082_044, w_082_049, w_082_051, w_082_053, w_082_058, w_082_059, w_082_066, w_082_069, w_082_070, w_082_073, w_082_079, w_082_082, w_082_090, w_082_092, w_082_104, w_082_106, w_082_112, w_082_115, w_082_122, w_082_123, w_082_128, w_082_130, w_082_135, w_082_139, w_082_140, w_082_141, w_082_142, w_082_148, w_082_150, w_082_154, w_082_160, w_082_162, w_082_166, w_082_167, w_082_175, w_082_191, w_082_193, w_082_196, w_082_199, w_082_213, w_082_214, w_082_215, w_082_218, w_082_228, w_082_235, w_082_240, w_082_244, w_082_247, w_082_270, w_082_291, w_082_299, w_082_303, w_082_309, w_082_314, w_082_323, w_082_336, w_082_338, w_082_383, w_082_389, w_082_393, w_082_409, w_082_423, w_082_425, w_082_431, w_082_455, w_082_463, w_082_486, w_082_487, w_082_502, w_082_505, w_082_511, w_082_526, w_082_531, w_082_538, w_082_540, w_082_541, w_082_546, w_082_551, w_082_576, w_082_577;
  wire w_083_007, w_083_008, w_083_009, w_083_011, w_083_013, w_083_017, w_083_018, w_083_019, w_083_021, w_083_022, w_083_023, w_083_033, w_083_036, w_083_040, w_083_043, w_083_044, w_083_046, w_083_052, w_083_057, w_083_061, w_083_066, w_083_067, w_083_068, w_083_071, w_083_073, w_083_085, w_083_088, w_083_093, w_083_098, w_083_103, w_083_110, w_083_113, w_083_115, w_083_116, w_083_118, w_083_123, w_083_127, w_083_129, w_083_135, w_083_138, w_083_140, w_083_144, w_083_147, w_083_149, w_083_151, w_083_153, w_083_154, w_083_155, w_083_156, w_083_158, w_083_163, w_083_165, w_083_166, w_083_168, w_083_169, w_083_170, w_083_175, w_083_181, w_083_182, w_083_183, w_083_187, w_083_189, w_083_190, w_083_191, w_083_192, w_083_193;
  wire w_084_000, w_084_001, w_084_002, w_084_003, w_084_004, w_084_005, w_084_006, w_084_007, w_084_008, w_084_009, w_084_010, w_084_011, w_084_012, w_084_013, w_084_014, w_084_015, w_084_016, w_084_017, w_084_018, w_084_020, w_084_021, w_084_023, w_084_024, w_084_025, w_084_026, w_084_028, w_084_029, w_084_030, w_084_032, w_084_033, w_084_034, w_084_036, w_084_037, w_084_038, w_084_039, w_084_040, w_084_042, w_084_043, w_084_044, w_084_045, w_084_046, w_084_047, w_084_048;
  wire w_085_001, w_085_011, w_085_015, w_085_016, w_085_017, w_085_022, w_085_024, w_085_026, w_085_027, w_085_028, w_085_029, w_085_030, w_085_034, w_085_037, w_085_038, w_085_040, w_085_042, w_085_045, w_085_048, w_085_051, w_085_056, w_085_059, w_085_068, w_085_070, w_085_074, w_085_080, w_085_084, w_085_085, w_085_087, w_085_088, w_085_092, w_085_096, w_085_116, w_085_125, w_085_129, w_085_139, w_085_141, w_085_146, w_085_150, w_085_152, w_085_158, w_085_161, w_085_162, w_085_164, w_085_167, w_085_173, w_085_176, w_085_190, w_085_199, w_085_201, w_085_202, w_085_203, w_085_205, w_085_219, w_085_220, w_085_226, w_085_230, w_085_244, w_085_246, w_085_255, w_085_257, w_085_265, w_085_272, w_085_277, w_085_294, w_085_295, w_085_298, w_085_299, w_085_305, w_085_306, w_085_309, w_085_320, w_085_327, w_085_329, w_085_338, w_085_340, w_085_349, w_085_350, w_085_353, w_085_355, w_085_356, w_085_357, w_085_358, w_085_359, w_085_360, w_085_361, w_085_362, w_085_364;
  wire w_086_003, w_086_007, w_086_009, w_086_010, w_086_022, w_086_024, w_086_028, w_086_029, w_086_032, w_086_033, w_086_034, w_086_043, w_086_046, w_086_049, w_086_051, w_086_055, w_086_059, w_086_062, w_086_064, w_086_065, w_086_067, w_086_073, w_086_078, w_086_081, w_086_083, w_086_089, w_086_091, w_086_093, w_086_095, w_086_097, w_086_098, w_086_101, w_086_119, w_086_122, w_086_124, w_086_133, w_086_134, w_086_144, w_086_151, w_086_158, w_086_160, w_086_161, w_086_164, w_086_173, w_086_175, w_086_179, w_086_181, w_086_182, w_086_185, w_086_187, w_086_189, w_086_190, w_086_192, w_086_195, w_086_197, w_086_201, w_086_208, w_086_232, w_086_236, w_086_237, w_086_253, w_086_264, w_086_265, w_086_270, w_086_275, w_086_277, w_086_307, w_086_312, w_086_313, w_086_320, w_086_321, w_086_332, w_086_336, w_086_343;
  wire w_087_013, w_087_015, w_087_018, w_087_025, w_087_028, w_087_037, w_087_040, w_087_043, w_087_048, w_087_051, w_087_054, w_087_058, w_087_065, w_087_069, w_087_071, w_087_086, w_087_088, w_087_098, w_087_100, w_087_102, w_087_106, w_087_117, w_087_118, w_087_120, w_087_125, w_087_127, w_087_134, w_087_137, w_087_149, w_087_154, w_087_156, w_087_160, w_087_162, w_087_165, w_087_168, w_087_182, w_087_186, w_087_189, w_087_190, w_087_195, w_087_204, w_087_205, w_087_207, w_087_215, w_087_216, w_087_219, w_087_227, w_087_228, w_087_230, w_087_235, w_087_243, w_087_247, w_087_249, w_087_253, w_087_255, w_087_258, w_087_273, w_087_286, w_087_292, w_087_293, w_087_298, w_087_310, w_087_311, w_087_323, w_087_326, w_087_333, w_087_335, w_087_343, w_087_357, w_087_358, w_087_366, w_087_372, w_087_379, w_087_381, w_087_387, w_087_407, w_087_408, w_087_425, w_087_431;
  wire w_088_002, w_088_003, w_088_005, w_088_011, w_088_012, w_088_013, w_088_015, w_088_016, w_088_018, w_088_019, w_088_020, w_088_021, w_088_022, w_088_023, w_088_024, w_088_025, w_088_028, w_088_029, w_088_031, w_088_032, w_088_033, w_088_036, w_088_041, w_088_043, w_088_044, w_088_045, w_088_046, w_088_048, w_088_050, w_088_051, w_088_052, w_088_053, w_088_055, w_088_060, w_088_061, w_088_062, w_088_063, w_088_065, w_088_066, w_088_067, w_088_069, w_088_070, w_088_076, w_088_079, w_088_080, w_088_089, w_088_090, w_088_093, w_088_094, w_088_102, w_088_106, w_088_117, w_088_119, w_088_121, w_088_125, w_088_126, w_088_129, w_088_130, w_088_131, w_088_132, w_088_135, w_088_136, w_088_143;
  wire w_089_006, w_089_009, w_089_012, w_089_013, w_089_017, w_089_025, w_089_026, w_089_028, w_089_033, w_089_042, w_089_045, w_089_051, w_089_053, w_089_055, w_089_057, w_089_060, w_089_061, w_089_068, w_089_070, w_089_071, w_089_072, w_089_075, w_089_078, w_089_085, w_089_086, w_089_089, w_089_094, w_089_096, w_089_098, w_089_100, w_089_106, w_089_107, w_089_111, w_089_118, w_089_126, w_089_128, w_089_129, w_089_132, w_089_134, w_089_135, w_089_136, w_089_138, w_089_140, w_089_142, w_089_144, w_089_149, w_089_150, w_089_151, w_089_155, w_089_156, w_089_160, w_089_164, w_089_166, w_089_167, w_089_178, w_089_185, w_089_190, w_089_191, w_089_197, w_089_198, w_089_199, w_089_206, w_089_210, w_089_211, w_089_213, w_089_215, w_089_217, w_089_219, w_089_221, w_089_230, w_089_232, w_089_258, w_089_259, w_089_266, w_089_269, w_089_282, w_089_289, w_089_291, w_089_300;
  wire w_090_001, w_090_011, w_090_016, w_090_035, w_090_036, w_090_042, w_090_047, w_090_048, w_090_052, w_090_061, w_090_063, w_090_066, w_090_067, w_090_068, w_090_072, w_090_080, w_090_086, w_090_088, w_090_117, w_090_122, w_090_126, w_090_131, w_090_151, w_090_168, w_090_171, w_090_191, w_090_195, w_090_203, w_090_206, w_090_218, w_090_221, w_090_222, w_090_223, w_090_224, w_090_232, w_090_242, w_090_266, w_090_272, w_090_275, w_090_295, w_090_306, w_090_310, w_090_358, w_090_362, w_090_370, w_090_380, w_090_384, w_090_392, w_090_405, w_090_415, w_090_420, w_090_442, w_090_451, w_090_464, w_090_469, w_090_472, w_090_478, w_090_487, w_090_489, w_090_505, w_090_510, w_090_523, w_090_528, w_090_531, w_090_532, w_090_535, w_090_536, w_090_542, w_090_543, w_090_564;
  wire w_091_000, w_091_008, w_091_012, w_091_014, w_091_020, w_091_024, w_091_028, w_091_030, w_091_032, w_091_033, w_091_034, w_091_036, w_091_037, w_091_039, w_091_040, w_091_041, w_091_042, w_091_043, w_091_044, w_091_046, w_091_056, w_091_059, w_091_063, w_091_067, w_091_073, w_091_074, w_091_075, w_091_077, w_091_078, w_091_080, w_091_081, w_091_085, w_091_088, w_091_091, w_091_094, w_091_095, w_091_105, w_091_109, w_091_111, w_091_112, w_091_117, w_091_119, w_091_122, w_091_123, w_091_125, w_091_127, w_091_129, w_091_133, w_091_134, w_091_135, w_091_137, w_091_143, w_091_144, w_091_151, w_091_152, w_091_153, w_091_154, w_091_157, w_091_160, w_091_161, w_091_162, w_091_163, w_091_164, w_091_166, w_091_169, w_091_170, w_091_176;
  wire w_092_001, w_092_009, w_092_011, w_092_027, w_092_029, w_092_032, w_092_043, w_092_045, w_092_046, w_092_049, w_092_050, w_092_059, w_092_062, w_092_068, w_092_070, w_092_073, w_092_080, w_092_088, w_092_089, w_092_107, w_092_112, w_092_131, w_092_151, w_092_154, w_092_159, w_092_162, w_092_189, w_092_190, w_092_191, w_092_200, w_092_203, w_092_209, w_092_220, w_092_225, w_092_229, w_092_242, w_092_264, w_092_272, w_092_277, w_092_287, w_092_292, w_092_307, w_092_324, w_092_331, w_092_360, w_092_377, w_092_391, w_092_412, w_092_429, w_092_439, w_092_447, w_092_458, w_092_471, w_092_478, w_092_480, w_092_481, w_092_484, w_092_489, w_092_492, w_092_494, w_092_504, w_092_516, w_092_530, w_092_548, w_092_551, w_092_560, w_092_562, w_092_563, w_092_572, w_092_580, w_092_588, w_092_595, w_092_609, w_092_610, w_092_628, w_092_636, w_092_650, w_092_673, w_092_690, w_092_715, w_092_724, w_092_725, w_092_726, w_092_728, w_092_730, w_092_731, w_092_732, w_092_733, w_092_734, w_092_735, w_092_736, w_092_738;
  wire w_093_006, w_093_016, w_093_028, w_093_032, w_093_035, w_093_041, w_093_043, w_093_050, w_093_054, w_093_055, w_093_057, w_093_059, w_093_060, w_093_067, w_093_073, w_093_077, w_093_080, w_093_081, w_093_084, w_093_086, w_093_088, w_093_089, w_093_091, w_093_097, w_093_101, w_093_105, w_093_119, w_093_123, w_093_128, w_093_132, w_093_133, w_093_143, w_093_151, w_093_162, w_093_177, w_093_178, w_093_180, w_093_186, w_093_200, w_093_208, w_093_217, w_093_224, w_093_225, w_093_239, w_093_245, w_093_252, w_093_256, w_093_270, w_093_321, w_093_332, w_093_339, w_093_354, w_093_360, w_093_362, w_093_371, w_093_389, w_093_390, w_093_391, w_093_393, w_093_395, w_093_409, w_093_413, w_093_417, w_093_420, w_093_421, w_093_430, w_093_442, w_093_448, w_093_458, w_093_497, w_093_504, w_093_560, w_093_561, w_093_562, w_093_563, w_093_565;
  wire w_094_006, w_094_009, w_094_021, w_094_027, w_094_038, w_094_043, w_094_044, w_094_051, w_094_052, w_094_056, w_094_057, w_094_064, w_094_079, w_094_083, w_094_095, w_094_101, w_094_110, w_094_114, w_094_116, w_094_120, w_094_138, w_094_150, w_094_159, w_094_162, w_094_167, w_094_173, w_094_182, w_094_193, w_094_195, w_094_222, w_094_234, w_094_246, w_094_267, w_094_271, w_094_286, w_094_288, w_094_296, w_094_299, w_094_317, w_094_336, w_094_344, w_094_363, w_094_370, w_094_373, w_094_376, w_094_380, w_094_381, w_094_386, w_094_387, w_094_399, w_094_419, w_094_421, w_094_432, w_094_434, w_094_440, w_094_444, w_094_449, w_094_462, w_094_469, w_094_475, w_094_514, w_094_522, w_094_527, w_094_534, w_094_542, w_094_544, w_094_545, w_094_546, w_094_564, w_094_574, w_094_587, w_094_599, w_094_600, w_094_607, w_094_609, w_094_610, w_094_624, w_094_663, w_094_664, w_094_665, w_094_666, w_094_667, w_094_669;
  wire w_095_000, w_095_001, w_095_002, w_095_003, w_095_004, w_095_005, w_095_006, w_095_008, w_095_010, w_095_012, w_095_014, w_095_018, w_095_019, w_095_021, w_095_022, w_095_023, w_095_026, w_095_027, w_095_029, w_095_030, w_095_031, w_095_033, w_095_034, w_095_036, w_095_038, w_095_039, w_095_040, w_095_041, w_095_042, w_095_043, w_095_046, w_095_047, w_095_049, w_095_051, w_095_052, w_095_053, w_095_054, w_095_055, w_095_056, w_095_057;
  wire w_096_000, w_096_001, w_096_002, w_096_003, w_096_004, w_096_005;
  wire w_097_002, w_097_004, w_097_007, w_097_009, w_097_012, w_097_016, w_097_033, w_097_035, w_097_038, w_097_039, w_097_042, w_097_048, w_097_049, w_097_056, w_097_061, w_097_063, w_097_070, w_097_077, w_097_082, w_097_085, w_097_088, w_097_090, w_097_102, w_097_105, w_097_108, w_097_118, w_097_121, w_097_122, w_097_125, w_097_130, w_097_131, w_097_135, w_097_139, w_097_142, w_097_144, w_097_153, w_097_166, w_097_175, w_097_179, w_097_180, w_097_189, w_097_195, w_097_201, w_097_205, w_097_207, w_097_212, w_097_224, w_097_225, w_097_252, w_097_303, w_097_331, w_097_335, w_097_360, w_097_366, w_097_373, w_097_374, w_097_393, w_097_430, w_097_471, w_097_480, w_097_492, w_097_502, w_097_504, w_097_507, w_097_514, w_097_521, w_097_526, w_097_548, w_097_553, w_097_566, w_097_570;
  wire w_098_000, w_098_001, w_098_003, w_098_004, w_098_005, w_098_008, w_098_009, w_098_010, w_098_011, w_098_012, w_098_013, w_098_014, w_098_015, w_098_016, w_098_017, w_098_018, w_098_019, w_098_020, w_098_022, w_098_024, w_098_025, w_098_027, w_098_028, w_098_031, w_098_032, w_098_033, w_098_034, w_098_035, w_098_036, w_098_038, w_098_040, w_098_041, w_098_042, w_098_043, w_098_044, w_098_045, w_098_046, w_098_047, w_098_048, w_098_050, w_098_052, w_098_053, w_098_055, w_098_057, w_098_058, w_098_059, w_098_061, w_098_062, w_098_063, w_098_065, w_098_068, w_098_069, w_098_071, w_098_074;
  wire w_099_001, w_099_002, w_099_003, w_099_011, w_099_015, w_099_019, w_099_025, w_099_036, w_099_037, w_099_044, w_099_047, w_099_051, w_099_053, w_099_054, w_099_055, w_099_057, w_099_058, w_099_059, w_099_062, w_099_068, w_099_070, w_099_071, w_099_075, w_099_077, w_099_078, w_099_081, w_099_087, w_099_088, w_099_091, w_099_093, w_099_101, w_099_107, w_099_111, w_099_113, w_099_114, w_099_123, w_099_131, w_099_133, w_099_135, w_099_136, w_099_141, w_099_148, w_099_150, w_099_159, w_099_163, w_099_169, w_099_172, w_099_173, w_099_174, w_099_178, w_099_180, w_099_188, w_099_192, w_099_205, w_099_213, w_099_222, w_099_223, w_099_229, w_099_240, w_099_248, w_099_256, w_099_257, w_099_261, w_099_262, w_099_263, w_099_274, w_099_276, w_099_278, w_099_291, w_099_302, w_099_303, w_099_304, w_099_305, w_099_306, w_099_307, w_099_308, w_099_309, w_099_310, w_099_311, w_099_312, w_099_313, w_099_317, w_099_318, w_099_319, w_099_320, w_099_321, w_099_322, w_099_323, w_099_324, w_099_325, w_099_326, w_099_327, w_099_329;
  wire w_100_002, w_100_007, w_100_008, w_100_010, w_100_012, w_100_013, w_100_014, w_100_018, w_100_019, w_100_021, w_100_022, w_100_024, w_100_030, w_100_031, w_100_036, w_100_037, w_100_038, w_100_044, w_100_046, w_100_049, w_100_051, w_100_053, w_100_055, w_100_056, w_100_057, w_100_058, w_100_060, w_100_061, w_100_063, w_100_065, w_100_066, w_100_071, w_100_074, w_100_077, w_100_078, w_100_080, w_100_081, w_100_082, w_100_084, w_100_085, w_100_086, w_100_087, w_100_092, w_100_093, w_100_094, w_100_095, w_100_096, w_100_100, w_100_106, w_100_109, w_100_113, w_100_115, w_100_116, w_100_120, w_100_121, w_100_125, w_100_127, w_100_130;
  wire w_101_003, w_101_004, w_101_006, w_101_008, w_101_020, w_101_038, w_101_049, w_101_050, w_101_056, w_101_063, w_101_066, w_101_070, w_101_077, w_101_083, w_101_085, w_101_089, w_101_090, w_101_092, w_101_094, w_101_095, w_101_098, w_101_104, w_101_107, w_101_121, w_101_122, w_101_124, w_101_130, w_101_135, w_101_139, w_101_143, w_101_156, w_101_158, w_101_166, w_101_168, w_101_170, w_101_171, w_101_176, w_101_188, w_101_194, w_101_207, w_101_209, w_101_214, w_101_223, w_101_238, w_101_243, w_101_244, w_101_246, w_101_247, w_101_253, w_101_258, w_101_261, w_101_266, w_101_269, w_101_272, w_101_280, w_101_283, w_101_284, w_101_285, w_101_293, w_101_294, w_101_303, w_101_307, w_101_313, w_101_314, w_101_315, w_101_316, w_101_317, w_101_321, w_101_322, w_101_323, w_101_325;
  wire w_102_014, w_102_022, w_102_025, w_102_028, w_102_035, w_102_036, w_102_042, w_102_047, w_102_050, w_102_060, w_102_068, w_102_070, w_102_076, w_102_093, w_102_097, w_102_115, w_102_116, w_102_123, w_102_133, w_102_144, w_102_152, w_102_181, w_102_183, w_102_188, w_102_193, w_102_195, w_102_199, w_102_204, w_102_226, w_102_229, w_102_246, w_102_248, w_102_250, w_102_252, w_102_274, w_102_282, w_102_304, w_102_308, w_102_316, w_102_329, w_102_333, w_102_337, w_102_345, w_102_364, w_102_368, w_102_392, w_102_421, w_102_424, w_102_436, w_102_442, w_102_445, w_102_451, w_102_458, w_102_462, w_102_476, w_102_479, w_102_491, w_102_505, w_102_523, w_102_526, w_102_529, w_102_542, w_102_546, w_102_550, w_102_553, w_102_555, w_102_561, w_102_563, w_102_575, w_102_589, w_102_597, w_102_601, w_102_609, w_102_618, w_102_619, w_102_646, w_102_648, w_102_649, w_102_650, w_102_651, w_102_652, w_102_653, w_102_654, w_102_655, w_102_659, w_102_660, w_102_661, w_102_662, w_102_663, w_102_665, w_102_667, w_102_668, w_102_669, w_102_670, w_102_671, w_102_672, w_102_673, w_102_674, w_102_675, w_102_676, w_102_680, w_102_681, w_102_682, w_102_683, w_102_684, w_102_685, w_102_686, w_102_687, w_102_688, w_102_690;
  wire w_103_002, w_103_006, w_103_007, w_103_015, w_103_016, w_103_023, w_103_026, w_103_045, w_103_048, w_103_053, w_103_054, w_103_056, w_103_059, w_103_063, w_103_064, w_103_067, w_103_068, w_103_072, w_103_075, w_103_076, w_103_083, w_103_084, w_103_092, w_103_098, w_103_105, w_103_108, w_103_113, w_103_114, w_103_117, w_103_121, w_103_123, w_103_128, w_103_136, w_103_137, w_103_140, w_103_143, w_103_145, w_103_147, w_103_149, w_103_156, w_103_162, w_103_168, w_103_185, w_103_191, w_103_195, w_103_199, w_103_206, w_103_210, w_103_213, w_103_220, w_103_228, w_103_230, w_103_232, w_103_240, w_103_248, w_103_260, w_103_264, w_103_287, w_103_289, w_103_292, w_103_301, w_103_313;
  wire w_104_000, w_104_004, w_104_007, w_104_009, w_104_021, w_104_025, w_104_029, w_104_033, w_104_040, w_104_042, w_104_047, w_104_053, w_104_057, w_104_062, w_104_063, w_104_067, w_104_068, w_104_073, w_104_080, w_104_091, w_104_100, w_104_109, w_104_112, w_104_131, w_104_137, w_104_138, w_104_143, w_104_144, w_104_152, w_104_157, w_104_158, w_104_162, w_104_168, w_104_178, w_104_179, w_104_188, w_104_193, w_104_197, w_104_199, w_104_213, w_104_216, w_104_221, w_104_228, w_104_233, w_104_256, w_104_260, w_104_263, w_104_264, w_104_266, w_104_271, w_104_273, w_104_278, w_104_280, w_104_284, w_104_290, w_104_291, w_104_298, w_104_299, w_104_310, w_104_311, w_104_321, w_104_323, w_104_326, w_104_335, w_104_342, w_104_354, w_104_357, w_104_362, w_104_366, w_104_370;
  wire w_105_001, w_105_005, w_105_016, w_105_029, w_105_045, w_105_052, w_105_079, w_105_082, w_105_088, w_105_091, w_105_093, w_105_097, w_105_102, w_105_120, w_105_123, w_105_129, w_105_130, w_105_132, w_105_134, w_105_144, w_105_163, w_105_169, w_105_182, w_105_192, w_105_198, w_105_199, w_105_200, w_105_202, w_105_211, w_105_213, w_105_216, w_105_218, w_105_220, w_105_226, w_105_229, w_105_235, w_105_241, w_105_248, w_105_249, w_105_251, w_105_253, w_105_264, w_105_265, w_105_267, w_105_268, w_105_274, w_105_282, w_105_284, w_105_294, w_105_305, w_105_325, w_105_327, w_105_331, w_105_336, w_105_339, w_105_346, w_105_351, w_105_364, w_105_372, w_105_384, w_105_386, w_105_388;
  wire w_106_000, w_106_006, w_106_012, w_106_021, w_106_023, w_106_025, w_106_027, w_106_032, w_106_037, w_106_043, w_106_044, w_106_050, w_106_051, w_106_052, w_106_054, w_106_058, w_106_062, w_106_065, w_106_066, w_106_067, w_106_069, w_106_072, w_106_075, w_106_076, w_106_081, w_106_083, w_106_084, w_106_089, w_106_091, w_106_093, w_106_096, w_106_098, w_106_101, w_106_105, w_106_107, w_106_108, w_106_116, w_106_123, w_106_124, w_106_127, w_106_129, w_106_138, w_106_139, w_106_140, w_106_141, w_106_144, w_106_146, w_106_147, w_106_160, w_106_162, w_106_165, w_106_170, w_106_181, w_106_183, w_106_199, w_106_204, w_106_206;
  wire w_107_003, w_107_005, w_107_021, w_107_047, w_107_054, w_107_056, w_107_068, w_107_080, w_107_082, w_107_091, w_107_094, w_107_096, w_107_097, w_107_100, w_107_103, w_107_109, w_107_115, w_107_118, w_107_121, w_107_125, w_107_126, w_107_130, w_107_150, w_107_151, w_107_157, w_107_159, w_107_161, w_107_177, w_107_180, w_107_181, w_107_183, w_107_186, w_107_211, w_107_219, w_107_220, w_107_221, w_107_238, w_107_252, w_107_256, w_107_258, w_107_259, w_107_272, w_107_279, w_107_288, w_107_292, w_107_293, w_107_302, w_107_304, w_107_310, w_107_313, w_107_318, w_107_329, w_107_345, w_107_349, w_107_355, w_107_370, w_107_379, w_107_396, w_107_400, w_107_415, w_107_425;
  wire w_108_000, w_108_001, w_108_002, w_108_003, w_108_006, w_108_015, w_108_021, w_108_024, w_108_026, w_108_031, w_108_035, w_108_040, w_108_053, w_108_057, w_108_065, w_108_067, w_108_073, w_108_078, w_108_085, w_108_086, w_108_087, w_108_090, w_108_095, w_108_097, w_108_103, w_108_115, w_108_119, w_108_122, w_108_127, w_108_130, w_108_132, w_108_143, w_108_145, w_108_150, w_108_159, w_108_161, w_108_166, w_108_174, w_108_182, w_108_183, w_108_188, w_108_190, w_108_197, w_108_200, w_108_201, w_108_203, w_108_205, w_108_207;
  wire w_109_002, w_109_003, w_109_005, w_109_009, w_109_011, w_109_028, w_109_053, w_109_054, w_109_068, w_109_100, w_109_104, w_109_114, w_109_124, w_109_127, w_109_131, w_109_152, w_109_169, w_109_177, w_109_199, w_109_204, w_109_209, w_109_213, w_109_217, w_109_219, w_109_229, w_109_233, w_109_238, w_109_240, w_109_251, w_109_252, w_109_259, w_109_264, w_109_279, w_109_280, w_109_282, w_109_284, w_109_285, w_109_291, w_109_293, w_109_327, w_109_331, w_109_350, w_109_352, w_109_358, w_109_363, w_109_374, w_109_383, w_109_385, w_109_392, w_109_394, w_109_407, w_109_457, w_109_473, w_109_474, w_109_486;
  wire w_110_004, w_110_017, w_110_022, w_110_026, w_110_032, w_110_039, w_110_041, w_110_042, w_110_047, w_110_064, w_110_075, w_110_087, w_110_090, w_110_092, w_110_117, w_110_124, w_110_125, w_110_132, w_110_135, w_110_139, w_110_147, w_110_148, w_110_154, w_110_171, w_110_175, w_110_187, w_110_196, w_110_197, w_110_210, w_110_237, w_110_239, w_110_242, w_110_246, w_110_250, w_110_260, w_110_262, w_110_273, w_110_275, w_110_277, w_110_279, w_110_282, w_110_289, w_110_290, w_110_294, w_110_295, w_110_304, w_110_318, w_110_327, w_110_335, w_110_352, w_110_358, w_110_362, w_110_363, w_110_364, w_110_376, w_110_386, w_110_401, w_110_405, w_110_410, w_110_425, w_110_459, w_110_462, w_110_463, w_110_464, w_110_465, w_110_466, w_110_468, w_110_470, w_110_471, w_110_472, w_110_473, w_110_474, w_110_475, w_110_477;
  wire w_111_003, w_111_007, w_111_008, w_111_010, w_111_011, w_111_012, w_111_018, w_111_019, w_111_020, w_111_021, w_111_023, w_111_027, w_111_034, w_111_039, w_111_041, w_111_046, w_111_047, w_111_049, w_111_054, w_111_059, w_111_061, w_111_062, w_111_070, w_111_078, w_111_081, w_111_091, w_111_099, w_111_102, w_111_106;
  wire w_112_000, w_112_006, w_112_008, w_112_010, w_112_018, w_112_019, w_112_021, w_112_022, w_112_025, w_112_035, w_112_039, w_112_046, w_112_054, w_112_056, w_112_063, w_112_065, w_112_068, w_112_077, w_112_078, w_112_079, w_112_084, w_112_085, w_112_095, w_112_104, w_112_107, w_112_120, w_112_121, w_112_127, w_112_130, w_112_131, w_112_134, w_112_140, w_112_143, w_112_144, w_112_145, w_112_160, w_112_161, w_112_165, w_112_169, w_112_172, w_112_173, w_112_174, w_112_180, w_112_182, w_112_187, w_112_189, w_112_197;
  wire w_113_008, w_113_010, w_113_015, w_113_019, w_113_025, w_113_029, w_113_031, w_113_032, w_113_033, w_113_034, w_113_047, w_113_048, w_113_049, w_113_050, w_113_061, w_113_062, w_113_081, w_113_090, w_113_106, w_113_107, w_113_109, w_113_110, w_113_112, w_113_114, w_113_120, w_113_125, w_113_132, w_113_136, w_113_146, w_113_154, w_113_158, w_113_171, w_113_172, w_113_174, w_113_181, w_113_185, w_113_187, w_113_188, w_113_198, w_113_209, w_113_211, w_113_218, w_113_219, w_113_227, w_113_231, w_113_234, w_113_237, w_113_238, w_113_250, w_113_258, w_113_262, w_113_267, w_113_269, w_113_273, w_113_276, w_113_289, w_113_291, w_113_300, w_113_309, w_113_316, w_113_318, w_113_323, w_113_341, w_113_347, w_113_348;
  wire w_114_003, w_114_007, w_114_009, w_114_015, w_114_018, w_114_020, w_114_032, w_114_036, w_114_037, w_114_039, w_114_047, w_114_056, w_114_058, w_114_065, w_114_067, w_114_068, w_114_069, w_114_106, w_114_112, w_114_114, w_114_116, w_114_117, w_114_118, w_114_119, w_114_120, w_114_131, w_114_134, w_114_135, w_114_138, w_114_141, w_114_144, w_114_148, w_114_150, w_114_152, w_114_167, w_114_170, w_114_176, w_114_181, w_114_186, w_114_188, w_114_189, w_114_194, w_114_195, w_114_197, w_114_198, w_114_209, w_114_211, w_114_217, w_114_220, w_114_226;
  wire w_115_000, w_115_004, w_115_005, w_115_008, w_115_016, w_115_018, w_115_019, w_115_021, w_115_033, w_115_036, w_115_037, w_115_039, w_115_040, w_115_055, w_115_061, w_115_065, w_115_066, w_115_075, w_115_084, w_115_089, w_115_101, w_115_122, w_115_125, w_115_126, w_115_131, w_115_134, w_115_135, w_115_136, w_115_151, w_115_152, w_115_162, w_115_169, w_115_178, w_115_179, w_115_190, w_115_191, w_115_194, w_115_209, w_115_215, w_115_219, w_115_228, w_115_240, w_115_241, w_115_251;
  wire w_116_001, w_116_004, w_116_008, w_116_023, w_116_030, w_116_042, w_116_061, w_116_077, w_116_079, w_116_092, w_116_112, w_116_118, w_116_122, w_116_124, w_116_126, w_116_136, w_116_140, w_116_142, w_116_150, w_116_153, w_116_192, w_116_204, w_116_224, w_116_231, w_116_238, w_116_260, w_116_261, w_116_287, w_116_292, w_116_343, w_116_345, w_116_348, w_116_365, w_116_373, w_116_387, w_116_407, w_116_412, w_116_414, w_116_420, w_116_424, w_116_426, w_116_428, w_116_495, w_116_497, w_116_500, w_116_510, w_116_513, w_116_530, w_116_532, w_116_545, w_116_554, w_116_570, w_116_576, w_116_601, w_116_628, w_116_636, w_116_639, w_116_640, w_116_641, w_116_642, w_116_643, w_116_644, w_116_645, w_116_646, w_116_647, w_116_648, w_116_649;
  wire w_117_000, w_117_004, w_117_005, w_117_008, w_117_010, w_117_011, w_117_012, w_117_014, w_117_016, w_117_017, w_117_018, w_117_020, w_117_022, w_117_024, w_117_026, w_117_028, w_117_029, w_117_033, w_117_035, w_117_036, w_117_038, w_117_040, w_117_043, w_117_045, w_117_046, w_117_048, w_117_050, w_117_051, w_117_053, w_117_054, w_117_055, w_117_056, w_117_057, w_117_058, w_117_059, w_117_060, w_117_062, w_117_063, w_117_064, w_117_066, w_117_072, w_117_074, w_117_075, w_117_078, w_117_079, w_117_088;
  wire w_118_000, w_118_005, w_118_010, w_118_012, w_118_017, w_118_018, w_118_019, w_118_023, w_118_029, w_118_030, w_118_031, w_118_036, w_118_040, w_118_041, w_118_043, w_118_050, w_118_054, w_118_060, w_118_061, w_118_062, w_118_067, w_118_070, w_118_071, w_118_079, w_118_080, w_118_081, w_118_082, w_118_087, w_118_090, w_118_093, w_118_094, w_118_099, w_118_101, w_118_104, w_118_107, w_118_108, w_118_109, w_118_110, w_118_111, w_118_112, w_118_113, w_118_114, w_118_115, w_118_116, w_118_117, w_118_118, w_118_122, w_118_123, w_118_124, w_118_125, w_118_126, w_118_127, w_118_128, w_118_129, w_118_130, w_118_132, w_118_134;
  wire w_119_001, w_119_003, w_119_007, w_119_012, w_119_014, w_119_016, w_119_017, w_119_018, w_119_027, w_119_029, w_119_040, w_119_043, w_119_050, w_119_053, w_119_063, w_119_067, w_119_070, w_119_082, w_119_083, w_119_085, w_119_086, w_119_087, w_119_099, w_119_101, w_119_103, w_119_104, w_119_106, w_119_109, w_119_117, w_119_119, w_119_123, w_119_125, w_119_135, w_119_139, w_119_142, w_119_143, w_119_146, w_119_149, w_119_156, w_119_157, w_119_162, w_119_164, w_119_165, w_119_171, w_119_175, w_119_177, w_119_188, w_119_189;
  wire w_120_008, w_120_029, w_120_038, w_120_042, w_120_051, w_120_060, w_120_072, w_120_083, w_120_104, w_120_126, w_120_135, w_120_140, w_120_159, w_120_167, w_120_169, w_120_176, w_120_177, w_120_215, w_120_222, w_120_223, w_120_241, w_120_244, w_120_262, w_120_269, w_120_289, w_120_305, w_120_311, w_120_332, w_120_343, w_120_345, w_120_348, w_120_353, w_120_402, w_120_410, w_120_430, w_120_439, w_120_454, w_120_480, w_120_489, w_120_506, w_120_516, w_120_517, w_120_528, w_120_545, w_120_558, w_120_569, w_120_578, w_120_594, w_120_604, w_120_612, w_120_626, w_120_633, w_120_638, w_120_648, w_120_666, w_120_674, w_120_681, w_120_684, w_120_689, w_120_693, w_120_695, w_120_734;
  wire w_121_004, w_121_009, w_121_011, w_121_027, w_121_032, w_121_039, w_121_045, w_121_047, w_121_048, w_121_050, w_121_051, w_121_053, w_121_054, w_121_055, w_121_057, w_121_058, w_121_082, w_121_084, w_121_086, w_121_088, w_121_106, w_121_112, w_121_115, w_121_117, w_121_120, w_121_121, w_121_125, w_121_126, w_121_127, w_121_128, w_121_129, w_121_134, w_121_136, w_121_141, w_121_144, w_121_160, w_121_161, w_121_162, w_121_168, w_121_174, w_121_189, w_121_190, w_121_192, w_121_194, w_121_199, w_121_202, w_121_206, w_121_209, w_121_210, w_121_211;
  wire w_122_000, w_122_001, w_122_005, w_122_008, w_122_009, w_122_010, w_122_012, w_122_014, w_122_017, w_122_020, w_122_021, w_122_022, w_122_026, w_122_027, w_122_030, w_122_031, w_122_032, w_122_034, w_122_035, w_122_040, w_122_041, w_122_049, w_122_055, w_122_056, w_122_058, w_122_060, w_122_063, w_122_065, w_122_066, w_122_067, w_122_072, w_122_074, w_122_081, w_122_082, w_122_083, w_122_084, w_122_086, w_122_089, w_122_090, w_122_091, w_122_093, w_122_094, w_122_102, w_122_103, w_122_113, w_122_120, w_122_121, w_122_126;
  wire w_123_005, w_123_013, w_123_016, w_123_029, w_123_036, w_123_053, w_123_056, w_123_067, w_123_087, w_123_096, w_123_097, w_123_101, w_123_104, w_123_112, w_123_122, w_123_139, w_123_149, w_123_153, w_123_162, w_123_169, w_123_172, w_123_174, w_123_187, w_123_195, w_123_251, w_123_255, w_123_297, w_123_302, w_123_304, w_123_364, w_123_367, w_123_369, w_123_379, w_123_388, w_123_459, w_123_471, w_123_481, w_123_503, w_123_505, w_123_511, w_123_532, w_123_538, w_123_584, w_123_592;
  wire w_124_001, w_124_025, w_124_027, w_124_035, w_124_046, w_124_052, w_124_056, w_124_057, w_124_061, w_124_065, w_124_070, w_124_078, w_124_089, w_124_091, w_124_094, w_124_096, w_124_104, w_124_105, w_124_108, w_124_109, w_124_112, w_124_114, w_124_116, w_124_122, w_124_134, w_124_143, w_124_145, w_124_156, w_124_171, w_124_217, w_124_220, w_124_232, w_124_242, w_124_244, w_124_252, w_124_256, w_124_273, w_124_281, w_124_286, w_124_287, w_124_291, w_124_295, w_124_319, w_124_328, w_124_330;
  wire w_125_003, w_125_025, w_125_030, w_125_031, w_125_036, w_125_057, w_125_059, w_125_065, w_125_069, w_125_072, w_125_079, w_125_081, w_125_084, w_125_118, w_125_124, w_125_128, w_125_129, w_125_138, w_125_150, w_125_187, w_125_191, w_125_193, w_125_204, w_125_208, w_125_224, w_125_242, w_125_282, w_125_297, w_125_308, w_125_318, w_125_332, w_125_347, w_125_354, w_125_386, w_125_397, w_125_399, w_125_417, w_125_439, w_125_446, w_125_466, w_125_497, w_125_561, w_125_586;
  wire w_126_008, w_126_013, w_126_017, w_126_018, w_126_024, w_126_027, w_126_028, w_126_034, w_126_037, w_126_038, w_126_041, w_126_047, w_126_055, w_126_056, w_126_058, w_126_061, w_126_063, w_126_064, w_126_068, w_126_073, w_126_078, w_126_079, w_126_082, w_126_084, w_126_090, w_126_092, w_126_095, w_126_100, w_126_104, w_126_112, w_126_115, w_126_116, w_126_117, w_126_119, w_126_120, w_126_127, w_126_128, w_126_130, w_126_133, w_126_135, w_126_139, w_126_142, w_126_144, w_126_153, w_126_154, w_126_158, w_126_164, w_126_175, w_126_187, w_126_193;
  wire w_127_000, w_127_003, w_127_004, w_127_007, w_127_008, w_127_011, w_127_015, w_127_017, w_127_018, w_127_022, w_127_025, w_127_026, w_127_027, w_127_031, w_127_034, w_127_035, w_127_038, w_127_041, w_127_043, w_127_044, w_127_047, w_127_048, w_127_052, w_127_053, w_127_054, w_127_057, w_127_061, w_127_065, w_127_067, w_127_069, w_127_070, w_127_071, w_127_073, w_127_074;
  wire w_128_000, w_128_010, w_128_021, w_128_022, w_128_025, w_128_026, w_128_035, w_128_048, w_128_051, w_128_055, w_128_067, w_128_070, w_128_073, w_128_091, w_128_094, w_128_103, w_128_111, w_128_115, w_128_122, w_128_130, w_128_139, w_128_140, w_128_152, w_128_157, w_128_174, w_128_181, w_128_187, w_128_191, w_128_195, w_128_196, w_128_233, w_128_234, w_128_268, w_128_291, w_128_295, w_128_297, w_128_306, w_128_318, w_128_327, w_128_329, w_128_345, w_128_353, w_128_380, w_128_411, w_128_414, w_128_417, w_128_426, w_128_464, w_128_495, w_128_496, w_128_524, w_128_559, w_128_571, w_128_580, w_128_608, w_128_638, w_128_640;
  wire w_129_005, w_129_017, w_129_023, w_129_029, w_129_034, w_129_041, w_129_044, w_129_048, w_129_065, w_129_067, w_129_072, w_129_078, w_129_082, w_129_087, w_129_088, w_129_090, w_129_095, w_129_100, w_129_106, w_129_108, w_129_111, w_129_113, w_129_117, w_129_120, w_129_133, w_129_135, w_129_140, w_129_149, w_129_156, w_129_164, w_129_168, w_129_170, w_129_175, w_129_180, w_129_182, w_129_186, w_129_198, w_129_204, w_129_205, w_129_210, w_129_216, w_129_226, w_129_245, w_129_251, w_129_256, w_129_275, w_129_276, w_129_278, w_129_282, w_129_289, w_129_293, w_129_295, w_129_305, w_129_313, w_129_329, w_129_333, w_129_337, w_129_342, w_129_348, w_129_349, w_129_351, w_129_353, w_129_372, w_129_414;
  wire w_130_005, w_130_023, w_130_033, w_130_035, w_130_044, w_130_046, w_130_049, w_130_071, w_130_075, w_130_088, w_130_089, w_130_122, w_130_134, w_130_171, w_130_184, w_130_191, w_130_194, w_130_195, w_130_204, w_130_211, w_130_212, w_130_220, w_130_230, w_130_236, w_130_239, w_130_252, w_130_254, w_130_260, w_130_264, w_130_278, w_130_280, w_130_283, w_130_294, w_130_295, w_130_321, w_130_375, w_130_377, w_130_391, w_130_408, w_130_418, w_130_463, w_130_469, w_130_499, w_130_511, w_130_518, w_130_519, w_130_520, w_130_521, w_130_522, w_130_523, w_130_524, w_130_528, w_130_529, w_130_530, w_130_531, w_130_532, w_130_533, w_130_534, w_130_535, w_130_536, w_130_538;
  wire w_131_000, w_131_007, w_131_029, w_131_037, w_131_040, w_131_048, w_131_053, w_131_054, w_131_059, w_131_071, w_131_073, w_131_087, w_131_092, w_131_101, w_131_109, w_131_113, w_131_120, w_131_121, w_131_140, w_131_144, w_131_147, w_131_149, w_131_187, w_131_212, w_131_223, w_131_254, w_131_263, w_131_269, w_131_285, w_131_303, w_131_304, w_131_308, w_131_318, w_131_345, w_131_430, w_131_431, w_131_432, w_131_450, w_131_472, w_131_480, w_131_483, w_131_486, w_131_511, w_131_545, w_131_557, w_131_566;
  wire w_132_012, w_132_026, w_132_031, w_132_056, w_132_059, w_132_076, w_132_077, w_132_082, w_132_084, w_132_087, w_132_089, w_132_094, w_132_099, w_132_115, w_132_129, w_132_130, w_132_152, w_132_155, w_132_165, w_132_179, w_132_180, w_132_188, w_132_196, w_132_202, w_132_204, w_132_206, w_132_217, w_132_219, w_132_229, w_132_231, w_132_249, w_132_255, w_132_260, w_132_262, w_132_281, w_132_289, w_132_291, w_132_305, w_132_313, w_132_330, w_132_331, w_132_333, w_132_384, w_132_386, w_132_390, w_132_393, w_132_395, w_132_398, w_132_406, w_132_415, w_132_422, w_132_435, w_132_467, w_132_468, w_132_469, w_132_470, w_132_471, w_132_475, w_132_476, w_132_477, w_132_478, w_132_479, w_132_480, w_132_481, w_132_483, w_132_485, w_132_486, w_132_487, w_132_488, w_132_489, w_132_490, w_132_491, w_132_492, w_132_493, w_132_494, w_132_495, w_132_496;
  wire w_133_000, w_133_003, w_133_028, w_133_057, w_133_061, w_133_066, w_133_081, w_133_085, w_133_095, w_133_097, w_133_099, w_133_117, w_133_120, w_133_134, w_133_143, w_133_159, w_133_187, w_133_201, w_133_223, w_133_235, w_133_244, w_133_249, w_133_290, w_133_313, w_133_334, w_133_344, w_133_351, w_133_362, w_133_368, w_133_373, w_133_374, w_133_376, w_133_378;
  wire w_134_001, w_134_002, w_134_017, w_134_018, w_134_066, w_134_071, w_134_072, w_134_073, w_134_076, w_134_089, w_134_109, w_134_114, w_134_116, w_134_122, w_134_132, w_134_135, w_134_138, w_134_140, w_134_147, w_134_151, w_134_156, w_134_163, w_134_169, w_134_173, w_134_185, w_134_200, w_134_204, w_134_218, w_134_230, w_134_251, w_134_256, w_134_261, w_134_292, w_134_320, w_134_323, w_134_374, w_134_375, w_134_396, w_134_405, w_134_448, w_134_451, w_134_474, w_134_489, w_134_490, w_134_491, w_134_492, w_134_493, w_134_494, w_134_495, w_134_496, w_134_497, w_134_498, w_134_499, w_134_501;
  wire w_135_003, w_135_013, w_135_019, w_135_029, w_135_062, w_135_078, w_135_086, w_135_089, w_135_094, w_135_110, w_135_111, w_135_119, w_135_136, w_135_156, w_135_163, w_135_164, w_135_184, w_135_191, w_135_194, w_135_196, w_135_200, w_135_240, w_135_257, w_135_271, w_135_286, w_135_348, w_135_354, w_135_373, w_135_377, w_135_398, w_135_429, w_135_438, w_135_457, w_135_487, w_135_488, w_135_528, w_135_549, w_135_587, w_135_609, w_135_661;
  wire w_136_002, w_136_004, w_136_005, w_136_007, w_136_010, w_136_011, w_136_013, w_136_014, w_136_017, w_136_020, w_136_024, w_136_025, w_136_030, w_136_031, w_136_032, w_136_033, w_136_037, w_136_040, w_136_044, w_136_047, w_136_049, w_136_051, w_136_054, w_136_057, w_136_058, w_136_059, w_136_060, w_136_063;
  wire w_137_003, w_137_013, w_137_017, w_137_032, w_137_034, w_137_037, w_137_039, w_137_042, w_137_045, w_137_061, w_137_075, w_137_076, w_137_085, w_137_098, w_137_099, w_137_104, w_137_107, w_137_116, w_137_122, w_137_123, w_137_146, w_137_162, w_137_164, w_137_176, w_137_183, w_137_185, w_137_188, w_137_190, w_137_202, w_137_223, w_137_234, w_137_235, w_137_255, w_137_266, w_137_272, w_137_320, w_137_345, w_137_351, w_137_354, w_137_356, w_137_443, w_137_464, w_137_469, w_137_473;
  wire w_138_023, w_138_024, w_138_037, w_138_047, w_138_049, w_138_051, w_138_056, w_138_058, w_138_060, w_138_061, w_138_066, w_138_067, w_138_069, w_138_073, w_138_078, w_138_083, w_138_093, w_138_094, w_138_096, w_138_100, w_138_104, w_138_120, w_138_125, w_138_134, w_138_157, w_138_160, w_138_168, w_138_171, w_138_192, w_138_205, w_138_206, w_138_214, w_138_221, w_138_231, w_138_238, w_138_241, w_138_246, w_138_248, w_138_250, w_138_258, w_138_261, w_138_282, w_138_283, w_138_304, w_138_308, w_138_309, w_138_310, w_138_326;
  wire w_139_001, w_139_002, w_139_004, w_139_005, w_139_006, w_139_007, w_139_009, w_139_010, w_139_011, w_139_013, w_139_014, w_139_015, w_139_016, w_139_018, w_139_019, w_139_020, w_139_021, w_139_022, w_139_023, w_139_024, w_139_025, w_139_026, w_139_027;
  wire w_140_001, w_140_009, w_140_010, w_140_015, w_140_020, w_140_021, w_140_024, w_140_027, w_140_031, w_140_036, w_140_042, w_140_052, w_140_062, w_140_068, w_140_071, w_140_073, w_140_074, w_140_088, w_140_092, w_140_093, w_140_094, w_140_096, w_140_137, w_140_155, w_140_161, w_140_165, w_140_176, w_140_178, w_140_180, w_140_184, w_140_188, w_140_189, w_140_190, w_140_202, w_140_216, w_140_230, w_140_233, w_140_234, w_140_242, w_140_243, w_140_244, w_140_245, w_140_246, w_140_247, w_140_251, w_140_252, w_140_253, w_140_254, w_140_256;
  wire w_141_000, w_141_002, w_141_008, w_141_011, w_141_012, w_141_016, w_141_018, w_141_021, w_141_044, w_141_048, w_141_050, w_141_053, w_141_056, w_141_059, w_141_065, w_141_068, w_141_079, w_141_093, w_141_107, w_141_114, w_141_117, w_141_128, w_141_133, w_141_139, w_141_143, w_141_149, w_141_151, w_141_154, w_141_168, w_141_171, w_141_175, w_141_176;
  wire w_142_040, w_142_076, w_142_095, w_142_101, w_142_129, w_142_147, w_142_181, w_142_187, w_142_205, w_142_209, w_142_212, w_142_258, w_142_276, w_142_303, w_142_321, w_142_348, w_142_365, w_142_421, w_142_442, w_142_494, w_142_499, w_142_503, w_142_517, w_142_559, w_142_587, w_142_603, w_142_607, w_142_638, w_142_772, w_142_777, w_142_792;
  wire w_143_000, w_143_004, w_143_014, w_143_018, w_143_019, w_143_044, w_143_061, w_143_066, w_143_068, w_143_076, w_143_081, w_143_082, w_143_088, w_143_090, w_143_106, w_143_107, w_143_111, w_143_116, w_143_209, w_143_211, w_143_243, w_143_257, w_143_265, w_143_300, w_143_344, w_143_353, w_143_374, w_143_401, w_143_408, w_143_473, w_143_479, w_143_493, w_143_501, w_143_530, w_143_535, w_143_554, w_143_568, w_143_575, w_143_581, w_143_598, w_143_652;
  wire w_144_006, w_144_010, w_144_032, w_144_035, w_144_043, w_144_044, w_144_045, w_144_061, w_144_062, w_144_077, w_144_079, w_144_105, w_144_125, w_144_142, w_144_169, w_144_173, w_144_182, w_144_185, w_144_186, w_144_190, w_144_193, w_144_202, w_144_206, w_144_219, w_144_228, w_144_242, w_144_302, w_144_306, w_144_309, w_144_346, w_144_373, w_144_406, w_144_447, w_144_473, w_144_558, w_144_559, w_144_560, w_144_561, w_144_562, w_144_563, w_144_564, w_144_565;
  wire w_145_002, w_145_005, w_145_011, w_145_012, w_145_016, w_145_020, w_145_022, w_145_027, w_145_030, w_145_032, w_145_035, w_145_037, w_145_038, w_145_039, w_145_040, w_145_046, w_145_048, w_145_052, w_145_066, w_145_068, w_145_070, w_145_075, w_145_077, w_145_079;
  wire w_146_001, w_146_005, w_146_008, w_146_036, w_146_042, w_146_044, w_146_049, w_146_057, w_146_071, w_146_079, w_146_085, w_146_088, w_146_090, w_146_092, w_146_107, w_146_124, w_146_133, w_146_142, w_146_168, w_146_182, w_146_191, w_146_198, w_146_210, w_146_213, w_146_227, w_146_255, w_146_256, w_146_273, w_146_275, w_146_279, w_146_285, w_146_291, w_146_297, w_146_302, w_146_303, w_146_305, w_146_309, w_146_311, w_146_320, w_146_321, w_146_323, w_146_324;
  wire w_147_003, w_147_007, w_147_020, w_147_022, w_147_027, w_147_029, w_147_031, w_147_032, w_147_037, w_147_040, w_147_050, w_147_061, w_147_062, w_147_063, w_147_077, w_147_089, w_147_097, w_147_099, w_147_100, w_147_113, w_147_116, w_147_118, w_147_146, w_147_147, w_147_160, w_147_162, w_147_165, w_147_166, w_147_168, w_147_173, w_147_175, w_147_202, w_147_203, w_147_214, w_147_216, w_147_226;
  wire w_148_004, w_148_010, w_148_015, w_148_017, w_148_038, w_148_043, w_148_060, w_148_077, w_148_085, w_148_087, w_148_106, w_148_123, w_148_164, w_148_209, w_148_215, w_148_241, w_148_279, w_148_283, w_148_286, w_148_353, w_148_371, w_148_375, w_148_398, w_148_417, w_148_447, w_148_499, w_148_528, w_148_536, w_148_553, w_148_565, w_148_574, w_148_576, w_148_581, w_148_595, w_148_609, w_148_611, w_148_650, w_148_670, w_148_684, w_148_689, w_148_690, w_148_691, w_148_692, w_148_693, w_148_694, w_148_698, w_148_699, w_148_700, w_148_701, w_148_702, w_148_703, w_148_705, w_148_707, w_148_708, w_148_709, w_148_710, w_148_711, w_148_712, w_148_713, w_148_717, w_148_718, w_148_719, w_148_721;
  wire w_149_004, w_149_015, w_149_018, w_149_027, w_149_032, w_149_041, w_149_056, w_149_060, w_149_063, w_149_075, w_149_079, w_149_080, w_149_081, w_149_082, w_149_126, w_149_138, w_149_159, w_149_179, w_149_207, w_149_261, w_149_302, w_149_314, w_149_364, w_149_367, w_149_368, w_149_430, w_149_438, w_149_450, w_149_466, w_149_478, w_149_484, w_149_501, w_149_506, w_149_517, w_149_590, w_149_600, w_149_612, w_149_619, w_149_631, w_149_636;
  wire w_150_000, w_150_003, w_150_008, w_150_009, w_150_041, w_150_056, w_150_067, w_150_068, w_150_108, w_150_127, w_150_150, w_150_159, w_150_182, w_150_191, w_150_197, w_150_200, w_150_231, w_150_239, w_150_241, w_150_253, w_150_274, w_150_294, w_150_296, w_150_300, w_150_318, w_150_324, w_150_333, w_150_334, w_150_345, w_150_361, w_150_363, w_150_378, w_150_393, w_150_394, w_150_449;
  wire w_151_009, w_151_011, w_151_013, w_151_034, w_151_048, w_151_057, w_151_068, w_151_080, w_151_086, w_151_088, w_151_099, w_151_108, w_151_116, w_151_130, w_151_148, w_151_156, w_151_160, w_151_175, w_151_178, w_151_184, w_151_200, w_151_203, w_151_208, w_151_215, w_151_222, w_151_247, w_151_259, w_151_262, w_151_264, w_151_268, w_151_276, w_151_284, w_151_295, w_151_302, w_151_321, w_151_352, w_151_366, w_151_367, w_151_388, w_151_453;
  wire w_152_002, w_152_007, w_152_008, w_152_045, w_152_073, w_152_089, w_152_108, w_152_118, w_152_153, w_152_161, w_152_167, w_152_198, w_152_200, w_152_221, w_152_234, w_152_236, w_152_337, w_152_348, w_152_387, w_152_428, w_152_468, w_152_511, w_152_513, w_152_573, w_152_586, w_152_601, w_152_621, w_152_714, w_152_721, w_152_729;
  wire w_153_009, w_153_016, w_153_018, w_153_019, w_153_020, w_153_022, w_153_025, w_153_026, w_153_029, w_153_030, w_153_032, w_153_037, w_153_038, w_153_044, w_153_045, w_153_047, w_153_049, w_153_052, w_153_053, w_153_055, w_153_056, w_153_057, w_153_060, w_153_067, w_153_070, w_153_072, w_153_073, w_153_085, w_153_091;
  wire w_154_002, w_154_009, w_154_010, w_154_025, w_154_030, w_154_031, w_154_033, w_154_036, w_154_039, w_154_046, w_154_051, w_154_054, w_154_055, w_154_056, w_154_060, w_154_062, w_154_065, w_154_075, w_154_078, w_154_080, w_154_082, w_154_093, w_154_094, w_154_095, w_154_096, w_154_097, w_154_098, w_154_099, w_154_103, w_154_110, w_154_112, w_154_119, w_154_120, w_154_121, w_154_131;
  wire w_155_000, w_155_001, w_155_024, w_155_033, w_155_034, w_155_041, w_155_045, w_155_050, w_155_072, w_155_076, w_155_088, w_155_090, w_155_102, w_155_103, w_155_109, w_155_122, w_155_145, w_155_148, w_155_149, w_155_180, w_155_192, w_155_197, w_155_217, w_155_242, w_155_252, w_155_276, w_155_288, w_155_289, w_155_290, w_155_352, w_155_402, w_155_403, w_155_405, w_155_415, w_155_424, w_155_443, w_155_444, w_155_470, w_155_493, w_155_494, w_155_508, w_155_531;
  wire w_156_005, w_156_007, w_156_013, w_156_029, w_156_032, w_156_041, w_156_044, w_156_057, w_156_100, w_156_130, w_156_150, w_156_167, w_156_172, w_156_209, w_156_224, w_156_231, w_156_232, w_156_238, w_156_242, w_156_261, w_156_289, w_156_296, w_156_342, w_156_374, w_156_386, w_156_428, w_156_430, w_156_467, w_156_472, w_156_501, w_156_545;
  wire w_157_001, w_157_002, w_157_007, w_157_013, w_157_021, w_157_022, w_157_031, w_157_032, w_157_036, w_157_048, w_157_051, w_157_053, w_157_054, w_157_058, w_157_064, w_157_065, w_157_066, w_157_074, w_157_094, w_157_097, w_157_098, w_157_101, w_157_121, w_157_123, w_157_124, w_157_126, w_157_133, w_157_135, w_157_141, w_157_148, w_157_151, w_157_160, w_157_162, w_157_164;
  wire w_158_000, w_158_001, w_158_002, w_158_003, w_158_004;
  wire w_159_004, w_159_007, w_159_008, w_159_012, w_159_013, w_159_018, w_159_024, w_159_029, w_159_030, w_159_032, w_159_037, w_159_039, w_159_045, w_159_048, w_159_063, w_159_065, w_159_074, w_159_077, w_159_078, w_159_079, w_159_080, w_159_083, w_159_098, w_159_101, w_159_108;
  wire w_160_039, w_160_049, w_160_056, w_160_059, w_160_063, w_160_074, w_160_080, w_160_092, w_160_148, w_160_182, w_160_223, w_160_237, w_160_245, w_160_299, w_160_382, w_160_394, w_160_398, w_160_405, w_160_426, w_160_433, w_160_449, w_160_465, w_160_479, w_160_580, w_160_601, w_160_611, w_160_634, w_160_667, w_160_673, w_160_699, w_160_706, w_160_753, w_160_793;
  wire w_161_009, w_161_013, w_161_023, w_161_026, w_161_035, w_161_065, w_161_071, w_161_074, w_161_079, w_161_093, w_161_121, w_161_133, w_161_134, w_161_135, w_161_153, w_161_155, w_161_160, w_161_183, w_161_272, w_161_294, w_161_326, w_161_365, w_161_369, w_161_394, w_161_446, w_161_451, w_161_460, w_161_461, w_161_472, w_161_487, w_161_514, w_161_533, w_161_565, w_161_567, w_161_607;
  wire w_162_000, w_162_001, w_162_002, w_162_003, w_162_004, w_162_006, w_162_008, w_162_013, w_162_015, w_162_017, w_162_019, w_162_020, w_162_021, w_162_022, w_162_023, w_162_024, w_162_025;
  wire w_163_036, w_163_050, w_163_065, w_163_077, w_163_078, w_163_081, w_163_091, w_163_099, w_163_132, w_163_133, w_163_157, w_163_159, w_163_162, w_163_163, w_163_178, w_163_185, w_163_188, w_163_189, w_163_221, w_163_225, w_163_228, w_163_243, w_163_249, w_163_266, w_163_284, w_163_307, w_163_327, w_163_343, w_163_416, w_163_428, w_163_445, w_163_478, w_163_486, w_163_488, w_163_489, w_163_491, w_163_497, w_163_509, w_163_515, w_163_519, w_163_567, w_163_574, w_163_593;
  wire w_164_004, w_164_005, w_164_023, w_164_079, w_164_085, w_164_093, w_164_119, w_164_127, w_164_141, w_164_204, w_164_235, w_164_241, w_164_244, w_164_266, w_164_277, w_164_291, w_164_294, w_164_302, w_164_339, w_164_348, w_164_374, w_164_387, w_164_390, w_164_395, w_164_424, w_164_453, w_164_502, w_164_588, w_164_593;
  wire w_165_003, w_165_007, w_165_009, w_165_012, w_165_015, w_165_017, w_165_025, w_165_026, w_165_028, w_165_032, w_165_034, w_165_043, w_165_049, w_165_050, w_165_051, w_165_054, w_165_056, w_165_059, w_165_071, w_165_079, w_165_088, w_165_094, w_165_095, w_165_096, w_165_101, w_165_105, w_165_109, w_165_110, w_165_111, w_165_146, w_165_150, w_165_155;
  wire w_166_010, w_166_040, w_166_041, w_166_056, w_166_076, w_166_081, w_166_095, w_166_097, w_166_103, w_166_109, w_166_110, w_166_115, w_166_123, w_166_127, w_166_138, w_166_145, w_166_152, w_166_165, w_166_199, w_166_202, w_166_219, w_166_248, w_166_268, w_166_279, w_166_282, w_166_287, w_166_288, w_166_299, w_166_305, w_166_313, w_166_322;
  wire w_167_005, w_167_014, w_167_016, w_167_022, w_167_031, w_167_040, w_167_041, w_167_043, w_167_049, w_167_050, w_167_057, w_167_068, w_167_078, w_167_080, w_167_081, w_167_082, w_167_099, w_167_100, w_167_107, w_167_108, w_167_122, w_167_131, w_167_140, w_167_145, w_167_152, w_167_162, w_167_163, w_167_164, w_167_165, w_167_166, w_167_170, w_167_171, w_167_172, w_167_173, w_167_174, w_167_175, w_167_176, w_167_177, w_167_178, w_167_179, w_167_180, w_167_181, w_167_183;
  wire w_168_014, w_168_028, w_168_088, w_168_110, w_168_126, w_168_143, w_168_147, w_168_151, w_168_152, w_168_159, w_168_171, w_168_216, w_168_232, w_168_266, w_168_315, w_168_354, w_168_359, w_168_380, w_168_381, w_168_419, w_168_448, w_168_452, w_168_492, w_168_506, w_168_542;
  wire w_169_004, w_169_008, w_169_062, w_169_101, w_169_103, w_169_106, w_169_141, w_169_170, w_169_187, w_169_192, w_169_200, w_169_218, w_169_221, w_169_236, w_169_273, w_169_279, w_169_283, w_169_296, w_169_303, w_169_305, w_169_318, w_169_323, w_169_333, w_169_344, w_169_365, w_169_380, w_169_405, w_169_437;
  wire w_170_015, w_170_017, w_170_040, w_170_053, w_170_085, w_170_139, w_170_172, w_170_185, w_170_194, w_170_198, w_170_209, w_170_212, w_170_222, w_170_226, w_170_240, w_170_248, w_170_250, w_170_277, w_170_282, w_170_310, w_170_331, w_170_399, w_170_423;
  wire w_171_013, w_171_119, w_171_124, w_171_135, w_171_162, w_171_176, w_171_192, w_171_195, w_171_221, w_171_228, w_171_252, w_171_263, w_171_265, w_171_303, w_171_322, w_171_333, w_171_334, w_171_363, w_171_384, w_171_408, w_171_412, w_171_425, w_171_450, w_171_470, w_171_479, w_171_495, w_171_560, w_171_578, w_171_606, w_171_611, w_171_654, w_171_706, w_171_711, w_171_722, w_171_731;
  wire w_172_000, w_172_001, w_172_002, w_172_003, w_172_005, w_172_006, w_172_007, w_172_012, w_172_013, w_172_024, w_172_030, w_172_031, w_172_033, w_172_035, w_172_039, w_172_040, w_172_041, w_172_042, w_172_044, w_172_046, w_172_048, w_172_049, w_172_052, w_172_053;
  wire w_173_001, w_173_002, w_173_003, w_173_004, w_173_005, w_173_008, w_173_009, w_173_011, w_173_012, w_173_013, w_173_015, w_173_016, w_173_017, w_173_018, w_173_022, w_173_023, w_173_025, w_173_026, w_173_027, w_173_028, w_173_030, w_173_031;
  wire w_174_001, w_174_004, w_174_010, w_174_014, w_174_024, w_174_028, w_174_029, w_174_044, w_174_060, w_174_066, w_174_072, w_174_075, w_174_083, w_174_088, w_174_090, w_174_092, w_174_093, w_174_096, w_174_098, w_174_104, w_174_107, w_174_110;
  wire w_175_018, w_175_019, w_175_022, w_175_025, w_175_026, w_175_038, w_175_056, w_175_083, w_175_103, w_175_108, w_175_141, w_175_144, w_175_156, w_175_167, w_175_208, w_175_221, w_175_240, w_175_285, w_175_373, w_175_417, w_175_422, w_175_464, w_175_477, w_175_488, w_175_504, w_175_549, w_175_558, w_175_594, w_175_615;
  wire w_176_001, w_176_002, w_176_008, w_176_049, w_176_059, w_176_080, w_176_085, w_176_097, w_176_110, w_176_129, w_176_136, w_176_138, w_176_148, w_176_151, w_176_158, w_176_170;
  wire w_177_006, w_177_008, w_177_014, w_177_024, w_177_025, w_177_036, w_177_085, w_177_102, w_177_108, w_177_160, w_177_166, w_177_178, w_177_238, w_177_258, w_177_266, w_177_280, w_177_288, w_177_307, w_177_310, w_177_333, w_177_375, w_177_385, w_177_399, w_177_402, w_177_405;
  wire w_178_005, w_178_006, w_178_009, w_178_015, w_178_028, w_178_036, w_178_043, w_178_049, w_178_054, w_178_067, w_178_075, w_178_076, w_178_077, w_178_095, w_178_097, w_178_099, w_178_102, w_178_107, w_178_114, w_178_115, w_178_116, w_178_118, w_178_120, w_178_121, w_178_122, w_178_123, w_178_124, w_178_125, w_178_126, w_178_127, w_178_128, w_178_129, w_178_131;
  wire w_179_023, w_179_039, w_179_044, w_179_079, w_179_140, w_179_141, w_179_159, w_179_164, w_179_184, w_179_188, w_179_203, w_179_204, w_179_416, w_179_423, w_179_507, w_179_579, w_179_583, w_179_620, w_179_710, w_179_721, w_179_737, w_179_745, w_179_767, w_179_768;
  wire w_180_001, w_180_002, w_180_003, w_180_007, w_180_008, w_180_009, w_180_010, w_180_011, w_180_012, w_180_013, w_180_014, w_180_015, w_180_016, w_180_019, w_180_020, w_180_021, w_180_023, w_180_024, w_180_025, w_180_026;
  wire w_181_002, w_181_039, w_181_048, w_181_058, w_181_064, w_181_118, w_181_123, w_181_132, w_181_142, w_181_147, w_181_153, w_181_169, w_181_195, w_181_205, w_181_208, w_181_249, w_181_265;
  wire w_182_002, w_182_004, w_182_005, w_182_007, w_182_009, w_182_010, w_182_011, w_182_013, w_182_015, w_182_016, w_182_017, w_182_018, w_182_021, w_182_023, w_182_024, w_182_025, w_182_026;
  wire w_183_005, w_183_008, w_183_011, w_183_018, w_183_025, w_183_031, w_183_039, w_183_041, w_183_073, w_183_092, w_183_103, w_183_111, w_183_118, w_183_119, w_183_131, w_183_133, w_183_139, w_183_164, w_183_183, w_183_193, w_183_194, w_183_202, w_183_243, w_183_244, w_183_270;
  wire w_184_000, w_184_007, w_184_011, w_184_019, w_184_025, w_184_029, w_184_032, w_184_033, w_184_038, w_184_041, w_184_049, w_184_052, w_184_056, w_184_065, w_184_073, w_184_112, w_184_130, w_184_132;
  wire w_185_023, w_185_027, w_185_039, w_185_049, w_185_059, w_185_069, w_185_072, w_185_076, w_185_090, w_185_094, w_185_100, w_185_103, w_185_104, w_185_108, w_185_109, w_185_112, w_185_130, w_185_137, w_185_140, w_185_185, w_185_198, w_185_202, w_185_209, w_185_219, w_185_220, w_185_221, w_185_222, w_185_223, w_185_224, w_185_225, w_185_226, w_185_227, w_185_228, w_185_229, w_185_231;
  wire w_186_042, w_186_055, w_186_084, w_186_093, w_186_095, w_186_099, w_186_131, w_186_140, w_186_177, w_186_197, w_186_205, w_186_208, w_186_212, w_186_223, w_186_231, w_186_235, w_186_257, w_186_262, w_186_295, w_186_322, w_186_336, w_186_361, w_186_440, w_186_450, w_186_467, w_186_537;
  wire w_187_001, w_187_002, w_187_004, w_187_006, w_187_009, w_187_010, w_187_011, w_187_012, w_187_013, w_187_014, w_187_015, w_187_016, w_187_017, w_187_019, w_187_020, w_187_023, w_187_026, w_187_028, w_187_029, w_187_030, w_187_032, w_187_033, w_187_039, w_187_041;
  wire w_188_003, w_188_007, w_188_036, w_188_039, w_188_062, w_188_091, w_188_107, w_188_146, w_188_158, w_188_184, w_188_225, w_188_281, w_188_393, w_188_437, w_188_592, w_188_646;
  wire w_189_023, w_189_025, w_189_026, w_189_056, w_189_092, w_189_119, w_189_157, w_189_175, w_189_220, w_189_298, w_189_319, w_189_367, w_189_443, w_189_445, w_189_446, w_189_463, w_189_471, w_189_478, w_189_484, w_189_513, w_189_546, w_189_620, w_189_621, w_189_622, w_189_623;
  wire w_190_000, w_190_001, w_190_005, w_190_008, w_190_009, w_190_014, w_190_029, w_190_034, w_190_036, w_190_040, w_190_041, w_190_053, w_190_066, w_190_067, w_190_073, w_190_074, w_190_093, w_190_095, w_190_096, w_190_100, w_190_103, w_190_112, w_190_116;
  wire w_191_008, w_191_011, w_191_026, w_191_027, w_191_033, w_191_034, w_191_045, w_191_047, w_191_051, w_191_052, w_191_062, w_191_065, w_191_069, w_191_074, w_191_076, w_191_082, w_191_092, w_191_134, w_191_136, w_191_163, w_191_210, w_191_215, w_191_229, w_191_232, w_191_240, w_191_245, w_191_262, w_191_275, w_191_286, w_191_306, w_191_309, w_191_331, w_191_336, w_191_362;
  wire w_192_008, w_192_009, w_192_010, w_192_017, w_192_019, w_192_031, w_192_041, w_192_045, w_192_059, w_192_063, w_192_065, w_192_079, w_192_082, w_192_099, w_192_113, w_192_114, w_192_119, w_192_134, w_192_138, w_192_145, w_192_146, w_192_148, w_192_153, w_192_163, w_192_164, w_192_165, w_192_172, w_192_175, w_192_176, w_192_179, w_192_189, w_192_196, w_192_197, w_192_198, w_192_199, w_192_200, w_192_201, w_192_202, w_192_203, w_192_204, w_192_205, w_192_206, w_192_207;
  wire w_193_006, w_193_014, w_193_021, w_193_033, w_193_067, w_193_080, w_193_085, w_193_087, w_193_091, w_193_097, w_193_106, w_193_131, w_193_136, w_193_137, w_193_151, w_193_169, w_193_183, w_193_184, w_193_190, w_193_199, w_193_233, w_193_272, w_193_296, w_193_299, w_193_312, w_193_327, w_193_345, w_193_350;
  wire w_194_021, w_194_057, w_194_077, w_194_078, w_194_096, w_194_098, w_194_102, w_194_117, w_194_132, w_194_136, w_194_142, w_194_170, w_194_173, w_194_174, w_194_178, w_194_187, w_194_221, w_194_238, w_194_241, w_194_246, w_194_262, w_194_298, w_194_304, w_194_314, w_194_325;
  wire w_195_003, w_195_006, w_195_007, w_195_023, w_195_030, w_195_035, w_195_044, w_195_046, w_195_054, w_195_067, w_195_072, w_195_074, w_195_075, w_195_081, w_195_084, w_195_100, w_195_107, w_195_121, w_195_128, w_195_129, w_195_139, w_195_140, w_195_141, w_195_148, w_195_177, w_195_194, w_195_205, w_195_208, w_195_209, w_195_216, w_195_228, w_195_232, w_195_233, w_195_236, w_195_241;
  wire w_196_007, w_196_016, w_196_023, w_196_040, w_196_072, w_196_075, w_196_079, w_196_095, w_196_101, w_196_111, w_196_136, w_196_141, w_196_149, w_196_154, w_196_163, w_196_173, w_196_196, w_196_210, w_196_212, w_196_217, w_196_254;
  wire w_197_017, w_197_060, w_197_064, w_197_098, w_197_114, w_197_141, w_197_146, w_197_152, w_197_160, w_197_161, w_197_194, w_197_223, w_197_228, w_197_247, w_197_248, w_197_312, w_197_396, w_197_445;
  wire w_198_006, w_198_014, w_198_017, w_198_021, w_198_024, w_198_030, w_198_044, w_198_046, w_198_052, w_198_053, w_198_054, w_198_056, w_198_057, w_198_059, w_198_060, w_198_062, w_198_076, w_198_078;
  wire w_199_040, w_199_048, w_199_054, w_199_073, w_199_076, w_199_106, w_199_156, w_199_159, w_199_173, w_199_178, w_199_235, w_199_240, w_199_253, w_199_266, w_199_267, w_199_280, w_199_294, w_199_338, w_199_373;
  wire w_200_002, w_200_005, w_200_021, w_200_028, w_200_045, w_200_061, w_200_089, w_200_106, w_200_117, w_200_127, w_200_128, w_200_178, w_200_183, w_200_188, w_200_211, w_200_214, w_200_216, w_200_234, w_200_254, w_200_282, w_200_359, w_200_407, w_200_429, w_200_436, w_200_440, w_200_448, w_200_498;
  wire w_201_007, w_201_009, w_201_026, w_201_027, w_201_035, w_201_057, w_201_062, w_201_081, w_201_141, w_201_148, w_201_174, w_201_190, w_201_193, w_201_203, w_201_226, w_201_268, w_201_280, w_201_286, w_201_346, w_201_409, w_201_422, w_201_502;
  wire w_202_014, w_202_017, w_202_022, w_202_029, w_202_033, w_202_040, w_202_055, w_202_064, w_202_066, w_202_077, w_202_078, w_202_079, w_202_085, w_202_089, w_202_095, w_202_105, w_202_111, w_202_116, w_202_119, w_202_149, w_202_153, w_202_165, w_202_184, w_202_186, w_202_196, w_202_198, w_202_218, w_202_223, w_202_231, w_202_252, w_202_267, w_202_276, w_202_278, w_202_286, w_202_292, w_202_295;
  wire w_203_015, w_203_016, w_203_027, w_203_032, w_203_045, w_203_062, w_203_074, w_203_083, w_203_090, w_203_143, w_203_184, w_203_198, w_203_246, w_203_259, w_203_271, w_203_297, w_203_339, w_203_368, w_203_375, w_203_430, w_203_433, w_203_444, w_203_473, w_203_478;
  wire w_204_011, w_204_027, w_204_043, w_204_056, w_204_135, w_204_218, w_204_280, w_204_323, w_204_386, w_204_388, w_204_473, w_204_493, w_204_510, w_204_651;
  wire w_205_000, w_205_007, w_205_034, w_205_035, w_205_053, w_205_066, w_205_076, w_205_122, w_205_153, w_205_173, w_205_186, w_205_199, w_205_216, w_205_217, w_205_245, w_205_285, w_205_309, w_205_317, w_205_330, w_205_353, w_205_367, w_205_453, w_205_459, w_205_462, w_205_504, w_205_519, w_205_537;
  wire w_206_002, w_206_009, w_206_010, w_206_038, w_206_046, w_206_047, w_206_058, w_206_070, w_206_082, w_206_086, w_206_087, w_206_119, w_206_139, w_206_144, w_206_145, w_206_157, w_206_203;
  wire w_207_026, w_207_049, w_207_050, w_207_069, w_207_086, w_207_110, w_207_119, w_207_144, w_207_152, w_207_189, w_207_198, w_207_202, w_207_233, w_207_263, w_207_378, w_207_463, w_207_468, w_207_546;
  wire w_208_021, w_208_026, w_208_027, w_208_035, w_208_053, w_208_072, w_208_083, w_208_122, w_208_133, w_208_161, w_208_169, w_208_175, w_208_214, w_208_225, w_208_231, w_208_238, w_208_244, w_208_259, w_208_268, w_208_273, w_208_277, w_208_354, w_208_400, w_208_408;
  wire w_209_007, w_209_012, w_209_018, w_209_033, w_209_043, w_209_054, w_209_057, w_209_062, w_209_063, w_209_065, w_209_087, w_209_106, w_209_139, w_209_140, w_209_145, w_209_176, w_209_182, w_209_209, w_209_255, w_209_263, w_209_281, w_209_299, w_209_314, w_209_322, w_209_342, w_209_345;
  wire w_210_003, w_210_014, w_210_019, w_210_020, w_210_028, w_210_030, w_210_040, w_210_044, w_210_061, w_210_064, w_210_093, w_210_098, w_210_101, w_210_102, w_210_107, w_210_124, w_210_132, w_210_139, w_210_142;
  wire w_211_003, w_211_004, w_211_005, w_211_006, w_211_012, w_211_014, w_211_017, w_211_018, w_211_019, w_211_021, w_211_023, w_211_026, w_211_027, w_211_028, w_211_033, w_211_034, w_211_036, w_211_037, w_211_039, w_211_040, w_211_041, w_211_042, w_211_043, w_211_044, w_211_045, w_211_046, w_211_047, w_211_048, w_211_049, w_211_051;
  wire w_212_003, w_212_006, w_212_009, w_212_019, w_212_034, w_212_048, w_212_052, w_212_061, w_212_064, w_212_067, w_212_073, w_212_087, w_212_092, w_212_117, w_212_120, w_212_124, w_212_162, w_212_163, w_212_165, w_212_170, w_212_182, w_212_189, w_212_190, w_212_202, w_212_204, w_212_218, w_212_226;
  wire w_213_005, w_213_007, w_213_013, w_213_015, w_213_017, w_213_046, w_213_052, w_213_070, w_213_078, w_213_079, w_213_085, w_213_086, w_213_179, w_213_194, w_213_241, w_213_303, w_213_315, w_213_339, w_213_358, w_213_368, w_213_392, w_213_414, w_213_419, w_213_466, w_213_479, w_213_513, w_213_541, w_213_577, w_213_600, w_213_605, w_213_665;
  wire w_214_010, w_214_016, w_214_021, w_214_055, w_214_148, w_214_166, w_214_175, w_214_181, w_214_201, w_214_203, w_214_206, w_214_225, w_214_280, w_214_371, w_214_381, w_214_448, w_214_457, w_214_518, w_214_550, w_214_577, w_214_594, w_214_595, w_214_596, w_214_597, w_214_598, w_214_599, w_214_600, w_214_604, w_214_605, w_214_606, w_214_607, w_214_608, w_214_609, w_214_610, w_214_611, w_214_612, w_214_613, w_214_614, w_214_616;
  wire w_215_015, w_215_024, w_215_025, w_215_038, w_215_049, w_215_099, w_215_106, w_215_124, w_215_138, w_215_139, w_215_166, w_215_197, w_215_203, w_215_206, w_215_211, w_215_246, w_215_249, w_215_286, w_215_335, w_215_344, w_215_346, w_215_429, w_215_434, w_215_438, w_215_487, w_215_494, w_215_532, w_215_533;
  wire w_216_002, w_216_034, w_216_044, w_216_048, w_216_088, w_216_105, w_216_149, w_216_169, w_216_203, w_216_234, w_216_236, w_216_253, w_216_262, w_216_281, w_216_290, w_216_301, w_216_308, w_216_340, w_216_345, w_216_352, w_216_357, w_216_362, w_216_376, w_216_377, w_216_410;
  wire w_217_001, w_217_006, w_217_008, w_217_014, w_217_018, w_217_020, w_217_023, w_217_031, w_217_034, w_217_049, w_217_051, w_217_054, w_217_060, w_217_061, w_217_064, w_217_068, w_217_074, w_217_078, w_217_083;
  wire w_218_080, w_218_124, w_218_178, w_218_180, w_218_189, w_218_195, w_218_261, w_218_334, w_218_338, w_218_380, w_218_576, w_218_584, w_218_595, w_218_599, w_218_660, w_218_671, w_218_698, w_218_701, w_218_725, w_218_776, w_218_777, w_218_778, w_218_779, w_218_780, w_218_781, w_218_782, w_218_783, w_218_784, w_218_785, w_218_789, w_218_790, w_218_791, w_218_792, w_218_793, w_218_794, w_218_795, w_218_796, w_218_797, w_218_798, w_218_799, w_218_800, w_218_802;
  wire w_219_005, w_219_008, w_219_067, w_219_090, w_219_242, w_219_244, w_219_265, w_219_340, w_219_413, w_219_439, w_219_522, w_219_604, w_219_626, w_219_636, w_219_644, w_219_656, w_219_668, w_219_738;
  wire w_220_119, w_220_142, w_220_186, w_220_195, w_220_197, w_220_231, w_220_248, w_220_263, w_220_265, w_220_290, w_220_322, w_220_337, w_220_340, w_220_346, w_220_350, w_220_367, w_220_371, w_220_377, w_220_380;
  wire w_221_018, w_221_033, w_221_044, w_221_054, w_221_063, w_221_067, w_221_069, w_221_071, w_221_125, w_221_143, w_221_159, w_221_175, w_221_190, w_221_207, w_221_213, w_221_225;
  wire w_222_026, w_222_032, w_222_120, w_222_141, w_222_163, w_222_185, w_222_226, w_222_236, w_222_255, w_222_315, w_222_321, w_222_422, w_222_469, w_222_521, w_222_623, w_222_628;
  wire w_223_016, w_223_027, w_223_040, w_223_047, w_223_073, w_223_075, w_223_079, w_223_140, w_223_141, w_223_145, w_223_146, w_223_151, w_223_156, w_223_166, w_223_184, w_223_201, w_223_202, w_223_209, w_223_218, w_223_235, w_223_241, w_223_267, w_223_284;
  wire w_224_024, w_224_036, w_224_049, w_224_069, w_224_083, w_224_095, w_224_104, w_224_113, w_224_114, w_224_156, w_224_178, w_224_210, w_224_241, w_224_256, w_224_303, w_224_331, w_224_353, w_224_386, w_224_401, w_224_405, w_224_421, w_224_494, w_224_524;
  wire w_225_010, w_225_019, w_225_033, w_225_051, w_225_053, w_225_059, w_225_062, w_225_086, w_225_102, w_225_104, w_225_112, w_225_142, w_225_154, w_225_168, w_225_180, w_225_194, w_225_204, w_225_220, w_225_227, w_225_240;
  wire w_226_019, w_226_077, w_226_092, w_226_138, w_226_152, w_226_171, w_226_189, w_226_190, w_226_199, w_226_219, w_226_222, w_226_310, w_226_393, w_226_401, w_226_455, w_226_475, w_226_497, w_226_557, w_226_558, w_226_559;
  wire w_227_026, w_227_036, w_227_062, w_227_160, w_227_163, w_227_173, w_227_209, w_227_231, w_227_269, w_227_278, w_227_339, w_227_403, w_227_475, w_227_485, w_227_513, w_227_584, w_227_597, w_227_612, w_227_620, w_227_647, w_227_658;
  wire w_228_005, w_228_011, w_228_013, w_228_039, w_228_050, w_228_066, w_228_105, w_228_123, w_228_146, w_228_214, w_228_343, w_228_374, w_228_466, w_228_533, w_228_578, w_228_580, w_228_584, w_228_588, w_228_625, w_228_627;
  wire w_229_000, w_229_003, w_229_015, w_229_034, w_229_035, w_229_041, w_229_046, w_229_086, w_229_136, w_229_192, w_229_247, w_229_268, w_229_285, w_229_323, w_229_455;
  wire w_230_007, w_230_010, w_230_024, w_230_027, w_230_037, w_230_038, w_230_055, w_230_060, w_230_077, w_230_080, w_230_095, w_230_157, w_230_197, w_230_215, w_230_233, w_230_266, w_230_298, w_230_321, w_230_322, w_230_323, w_230_324, w_230_325, w_230_326, w_230_327, w_230_328, w_230_329, w_230_333, w_230_334, w_230_335, w_230_336, w_230_337, w_230_338, w_230_339, w_230_340, w_230_341, w_230_342, w_230_344;
  wire w_231_001, w_231_003, w_231_009, w_231_056, w_231_064, w_231_157, w_231_160, w_231_198, w_231_199, w_231_220, w_231_321, w_231_322, w_231_427, w_231_463, w_231_464, w_231_530, w_231_532, w_231_537, w_231_545, w_231_579;
  wire w_232_035, w_232_050, w_232_069, w_232_077, w_232_079, w_232_084, w_232_103, w_232_125, w_232_150, w_232_166, w_232_172, w_232_190, w_232_237, w_232_295, w_232_318, w_232_332, w_232_376, w_232_381, w_232_399, w_232_456, w_232_457, w_232_478, w_232_479, w_232_503, w_232_508, w_232_509, w_232_510, w_232_511, w_232_512, w_232_513, w_232_517, w_232_518, w_232_519, w_232_520, w_232_521, w_232_522, w_232_523, w_232_524, w_232_525, w_232_526, w_232_527, w_232_529;
  wire w_233_001, w_233_012, w_233_037, w_233_038, w_233_068, w_233_088, w_233_101, w_233_168, w_233_169, w_233_171, w_233_204, w_233_234, w_233_239, w_233_249, w_233_326, w_233_353, w_233_378, w_233_386;
  wire w_234_038, w_234_086, w_234_111, w_234_145, w_234_147, w_234_153, w_234_159, w_234_182, w_234_195, w_234_254, w_234_309, w_234_326, w_234_403, w_234_429;
  wire w_235_018, w_235_034, w_235_046, w_235_056, w_235_062, w_235_066, w_235_070, w_235_079, w_235_083, w_235_101, w_235_112, w_235_114, w_235_115, w_235_121, w_235_141, w_235_177, w_235_181, w_235_206;
  wire w_236_010, w_236_028, w_236_046, w_236_097, w_236_132, w_236_159, w_236_166, w_236_199;
  wire w_237_000, w_237_012, w_237_033, w_237_062, w_237_063, w_237_074, w_237_081, w_237_084, w_237_107, w_237_111, w_237_128, w_237_130, w_237_131, w_237_134;
  wire w_238_000, w_238_010, w_238_021, w_238_052, w_238_105, w_238_120, w_238_141, w_238_150, w_238_189, w_238_195, w_238_235, w_238_264, w_238_395, w_238_412, w_238_429, w_238_449;
  wire w_239_000;
  wire w_240_005, w_240_019, w_240_024, w_240_026, w_240_038, w_240_047, w_240_055, w_240_056, w_240_072, w_240_076, w_240_090, w_240_098, w_240_101, w_240_104, w_240_109, w_240_114, w_240_125, w_240_142, w_240_147, w_240_159, w_240_171, w_240_184;
  wire w_241_000, w_241_002, w_241_008, w_241_010, w_241_011, w_241_021, w_241_029, w_241_030, w_241_031, w_241_032, w_241_033, w_241_055, w_241_058, w_241_059, w_241_068, w_241_081, w_241_085;
  wire w_242_000, w_242_002, w_242_006, w_242_058, w_242_077, w_242_082, w_242_090, w_242_093, w_242_122, w_242_132, w_242_133, w_242_134, w_242_153, w_242_162, w_242_163;
  wire w_243_015, w_243_057, w_243_072, w_243_109, w_243_111, w_243_143, w_243_150, w_243_160, w_243_181, w_243_268, w_243_297;
  wire w_244_000, w_244_026, w_244_053, w_244_071, w_244_081, w_244_111, w_244_117, w_244_136, w_244_185, w_244_200, w_244_205, w_244_216, w_244_220, w_244_229, w_244_238, w_244_244, w_244_247, w_244_248, w_244_249, w_244_250, w_244_251, w_244_252, w_244_254;
  wire w_245_035, w_245_153, w_245_155, w_245_188, w_245_262, w_245_339, w_245_347, w_245_397, w_245_398, w_245_436, w_245_448, w_245_465, w_245_507, w_245_624, w_245_660, w_245_696, w_245_730, w_245_735;
  wire w_246_014, w_246_074, w_246_075, w_246_079, w_246_092, w_246_107, w_246_119, w_246_124, w_246_286, w_246_289, w_246_307, w_246_482, w_246_485, w_246_520, w_246_521, w_246_573, w_246_593, w_246_607, w_246_608;
  wire w_247_000, w_247_021, w_247_035, w_247_076, w_247_079, w_247_107, w_247_131, w_247_135, w_247_140, w_247_142, w_247_147, w_247_154, w_247_159, w_247_161, w_247_162, w_247_163, w_247_170, w_247_181, w_247_183, w_247_184;
  wire w_248_025, w_248_028, w_248_034, w_248_039, w_248_042, w_248_045, w_248_063, w_248_087, w_248_099, w_248_111, w_248_130, w_248_136, w_248_142;
  wire w_249_069, w_249_150, w_249_152, w_249_169, w_249_187, w_249_191, w_249_202, w_249_268, w_249_280, w_249_333, w_249_340;
  wire w_250_012, w_250_239, w_250_252, w_250_287, w_250_288, w_250_292, w_250_327, w_250_367, w_250_513, w_250_548, w_250_588, w_250_605, w_250_609;
  wire w_251_013, w_251_017, w_251_028, w_251_035, w_251_037, w_251_047, w_251_048, w_251_064, w_251_075, w_251_081, w_251_089, w_251_097, w_251_109, w_251_112, w_251_130, w_251_131, w_251_133;
  wire w_252_012, w_252_044, w_252_065, w_252_088, w_252_103, w_252_124, w_252_229, w_252_242, w_252_247, w_252_272, w_252_275, w_252_280, w_252_301, w_252_306, w_252_331, w_252_363, w_252_368, w_252_386, w_252_394, w_252_429, w_252_430, w_252_431, w_252_432, w_252_433, w_252_434, w_252_435, w_252_436, w_252_437;
  wire w_253_002, w_253_008, w_253_023, w_253_053, w_253_059, w_253_060, w_253_074, w_253_143, w_253_150, w_253_163, w_253_198, w_253_221, w_253_318, w_253_344, w_253_361, w_253_363, w_253_415;
  wire w_254_000, w_254_020, w_254_028, w_254_031, w_254_037, w_254_053, w_254_054, w_254_057, w_254_058, w_254_061, w_254_062, w_254_065, w_254_073, w_254_084, w_254_095, w_254_105, w_254_106, w_254_107, w_254_108, w_254_109, w_254_110, w_254_111, w_254_112, w_254_113;
  wire w_255_024, w_255_035, w_255_042, w_255_062, w_255_076, w_255_078, w_255_081, w_255_089, w_255_103, w_255_105;
  wire w_256_021, w_256_028, w_256_060, w_256_089, w_256_097, w_256_310, w_256_477, w_256_484, w_256_490, w_256_515, w_256_550, w_256_646, w_256_689;
  wire w_257_054, w_257_075, w_257_101, w_257_110, w_257_112, w_257_143, w_257_190, w_257_243, w_257_257, w_257_293, w_257_318;
  wire w_258_026, w_258_032, w_258_103, w_258_138, w_258_153, w_258_193, w_258_240, w_258_247, w_258_390, w_258_411, w_258_449, w_258_481;
  wire w_259_038, w_259_084, w_259_131, w_259_224, w_259_316, w_259_338, w_259_345, w_259_457, w_259_469, w_259_472, w_259_506, w_259_543, w_259_551;
  wire w_260_001, w_260_017, w_260_027, w_260_030, w_260_035, w_260_058, w_260_061, w_260_082, w_260_101, w_260_108, w_260_151, w_260_159, w_260_161, w_260_164, w_260_166, w_260_183, w_260_199, w_260_201, w_260_282, w_260_283, w_260_284, w_260_285, w_260_286, w_260_287, w_260_288, w_260_292, w_260_293, w_260_294, w_260_295, w_260_296, w_260_297, w_260_298, w_260_299, w_260_300, w_260_301, w_260_302, w_260_304;
  wire w_261_000, w_261_005, w_261_008, w_261_015, w_261_022, w_261_029, w_261_032, w_261_034, w_261_041, w_261_044, w_261_061, w_261_100;
  wire w_262_001, w_262_002, w_262_010, w_262_044, w_262_068, w_262_073, w_262_202, w_262_223, w_262_267, w_262_321, w_262_371, w_262_381, w_262_389;
  wire w_263_001, w_263_007, w_263_022, w_263_028, w_263_030, w_263_049, w_263_062, w_263_078, w_263_083, w_263_101, w_263_104, w_263_106, w_263_119, w_263_120, w_263_133;
  wire w_264_157, w_264_159, w_264_161, w_264_233, w_264_266, w_264_273, w_264_310, w_264_470, w_264_553, w_264_599, w_264_666, w_264_743;
  wire w_265_029, w_265_064, w_265_073, w_265_120, w_265_171, w_265_197, w_265_237, w_265_327, w_265_418, w_265_450, w_265_453, w_265_491, w_265_507, w_265_641, w_265_645, w_265_694;
  wire w_266_043, w_266_124, w_266_160, w_266_176, w_266_247, w_266_250, w_266_307, w_266_324, w_266_330, w_266_438, w_266_533, w_266_621, w_266_622, w_266_623, w_266_624, w_266_625, w_266_626, w_266_627, w_266_628, w_266_629, w_266_630, w_266_631, w_266_635, w_266_636, w_266_637, w_266_638, w_266_639, w_266_640, w_266_641, w_266_642, w_266_643, w_266_645;
  wire w_267_014, w_267_023, w_267_041, w_267_054, w_267_055, w_267_065, w_267_067, w_267_083, w_267_085, w_267_103, w_267_114, w_267_131, w_267_146, w_267_155, w_267_183, w_267_216, w_267_217, w_267_248, w_267_276, w_267_298;
  wire w_268_021, w_268_035, w_268_038, w_268_058, w_268_079, w_268_113, w_268_152, w_268_213, w_268_214, w_268_216, w_268_237, w_268_261, w_268_268;
  wire w_269_019, w_269_030, w_269_070, w_269_122, w_269_159, w_269_171, w_269_276, w_269_356, w_269_363, w_269_382, w_269_405, w_269_414, w_269_434, w_269_441, w_269_493, w_269_564, w_269_565;
  wire w_270_017, w_270_037, w_270_046, w_270_217, w_270_228, w_270_284, w_270_335;
  wire w_271_011, w_271_021, w_271_030, w_271_072, w_271_142, w_271_188, w_271_354, w_271_416, w_271_470, w_271_532, w_271_555, w_271_575, w_271_602, w_271_637, w_271_740;
  wire w_272_005, w_272_009, w_272_018, w_272_021, w_272_024, w_272_026, w_272_028, w_272_030, w_272_031, w_272_038, w_272_039, w_272_040, w_272_043;
  wire w_273_042, w_273_054, w_273_065, w_273_075, w_273_092, w_273_093, w_273_105, w_273_112, w_273_134, w_273_135, w_273_136, w_273_137, w_273_138, w_273_139, w_273_140, w_273_141, w_273_142;
  wire w_274_029, w_274_055, w_274_100, w_274_104, w_274_115, w_274_126, w_274_130, w_274_143, w_274_144, w_274_149, w_274_170, w_274_171, w_274_188, w_274_221, w_274_232, w_274_238;
  wire w_275_049, w_275_090, w_275_133, w_275_135, w_275_291, w_275_489, w_275_598, w_275_603, w_275_605, w_275_619, w_275_722;
  wire w_276_030, w_276_050, w_276_110, w_276_142, w_276_170, w_276_185, w_276_196, w_276_200, w_276_264, w_276_296, w_276_326, w_276_331, w_276_349, w_276_350, w_276_367;
  wire w_277_013, w_277_020, w_277_038, w_277_067, w_277_123, w_277_137, w_277_143, w_277_203, w_277_258, w_277_268, w_277_293, w_277_315, w_277_317, w_277_364, w_277_373, w_277_381;
  wire w_278_045, w_278_057, w_278_060, w_278_100, w_278_116, w_278_174;
  wire w_279_026, w_279_068, w_279_069, w_279_124, w_279_127, w_279_138, w_279_139, w_279_153, w_279_160, w_279_171, w_279_228, w_279_253, w_279_302;
  wire w_280_019, w_280_098, w_280_258, w_280_259, w_280_282, w_280_306, w_280_444, w_280_448, w_280_503, w_280_559, w_280_652, w_280_682, w_280_687;
  wire w_281_044, w_281_089, w_281_119, w_281_133, w_281_212, w_281_237, w_281_283, w_281_307, w_281_365, w_281_389, w_281_462, w_281_551, w_281_616, w_281_627, w_281_643, w_281_710, w_281_740;
  wire w_282_031, w_282_109, w_282_110, w_282_137, w_282_141, w_282_150, w_282_166, w_282_206, w_282_227, w_282_236, w_282_246, w_282_250, w_282_265, w_282_291, w_282_298, w_282_327, w_282_367, w_282_385, w_282_386, w_282_387, w_282_388, w_282_392, w_282_393, w_282_394, w_282_395, w_282_397;
  wire w_283_003, w_283_038, w_283_043, w_283_064, w_283_094, w_283_126, w_283_131, w_283_137, w_283_138, w_283_216, w_283_219, w_283_272, w_283_329, w_283_338, w_283_379;
  wire w_284_005, w_284_014, w_284_015, w_284_022, w_284_024, w_284_029, w_284_039, w_284_040, w_284_049, w_284_054, w_284_080, w_284_081, w_284_102, w_284_113, w_284_123, w_284_129, w_284_142, w_284_145;
  wire w_285_011, w_285_037, w_285_041, w_285_057, w_285_091, w_285_104, w_285_184, w_285_353, w_285_393, w_285_460, w_285_689, w_285_774;
  wire w_286_037, w_286_074, w_286_130, w_286_132, w_286_136, w_286_186, w_286_190, w_286_275, w_286_362, w_286_377, w_286_380, w_286_393;
  wire w_287_019, w_287_020, w_287_064, w_287_125, w_287_180, w_287_274, w_287_279, w_287_315, w_287_334, w_287_335, w_287_354, w_287_369, w_287_394;
  wire w_288_068, w_288_070, w_288_087, w_288_158, w_288_167, w_288_194, w_288_198, w_288_278, w_288_288, w_288_420, w_288_422, w_288_478, w_288_510, w_288_511, w_288_512, w_288_516, w_288_517, w_288_518, w_288_519, w_288_520, w_288_521, w_288_522, w_288_523, w_288_524, w_288_526;
  wire w_289_103, w_289_121, w_289_166, w_289_257, w_289_417, w_289_574;
  wire w_290_004, w_290_005, w_290_048, w_290_086, w_290_100, w_290_103, w_290_106, w_290_117, w_290_118, w_290_128, w_290_158, w_290_159, w_290_160, w_290_161, w_290_162, w_290_163, w_290_164, w_290_165, w_290_166, w_290_167;
  wire w_291_001, w_291_007, w_291_022, w_291_030, w_291_043, w_291_044, w_291_063, w_291_071, w_291_073, w_291_082, w_291_085, w_291_099, w_291_108, w_291_110, w_291_123, w_291_129;
  wire w_292_033, w_292_298, w_292_309, w_292_433, w_292_494, w_292_533, w_292_554;
  wire w_293_021, w_293_033, w_293_036, w_293_038, w_293_067, w_293_084, w_293_101, w_293_149, w_293_208, w_293_225, w_293_226, w_293_325, w_293_359, w_293_386;
  wire w_294_000, w_294_009, w_294_017, w_294_019, w_294_031, w_294_037, w_294_046, w_294_055, w_294_064, w_294_070, w_294_074, w_294_083, w_294_110, w_294_111, w_294_118, w_294_145, w_294_148;
  wire w_295_020, w_295_092, w_295_112, w_295_122, w_295_173, w_295_188, w_295_227, w_295_247, w_295_275, w_295_280, w_295_308, w_295_312, w_295_400;
  wire w_296_032, w_296_041, w_296_129, w_296_132, w_296_200, w_296_302, w_296_316, w_296_354;
  wire w_297_054, w_297_116;
  wire w_298_000, w_298_003, w_298_019, w_298_031, w_298_035, w_298_038, w_298_057, w_298_073, w_298_087, w_298_090, w_298_091, w_298_099, w_298_100;
  wire w_299_015, w_299_020, w_299_050, w_299_053, w_299_097, w_299_149, w_299_164, w_299_245, w_299_261, w_299_270, w_299_288, w_299_315, w_299_316, w_299_476, w_299_477, w_299_478, w_299_479, w_299_480, w_299_481, w_299_482, w_299_483, w_299_484, w_299_485, w_299_486, w_299_490, w_299_491, w_299_492, w_299_494;
  wire w_300_010, w_300_046, w_300_064, w_300_085, w_300_111, w_300_139, w_300_176, w_300_261, w_300_425, w_300_610;
  wire w_301_002, w_301_014, w_301_027, w_301_046, w_301_062, w_301_066, w_301_091, w_301_121, w_301_153, w_301_182, w_301_197, w_301_210, w_301_220;
  wire w_302_049, w_302_076, w_302_117, w_302_261, w_302_338, w_302_495, w_302_529, w_302_629;
  wire w_303_059, w_303_070, w_303_078, w_303_080, w_303_095, w_303_100, w_303_106, w_303_119, w_303_121, w_303_128;
  wire w_304_003, w_304_022, w_304_079, w_304_083, w_304_100, w_304_178, w_304_192, w_304_223, w_304_258, w_304_315, w_304_331, w_304_414, w_304_437, w_304_443, w_304_468, w_304_500;
  wire w_305_057, w_305_077, w_305_083, w_305_103, w_305_157, w_305_178, w_305_188, w_305_239, w_305_270, w_305_471, w_305_536;
  wire w_306_018, w_306_041, w_306_087, w_306_106, w_306_112, w_306_146, w_306_151, w_306_165, w_306_177, w_306_207, w_306_236, w_306_272, w_306_281;
  wire w_307_036, w_307_040, w_307_043, w_307_075, w_307_081, w_307_093, w_307_095, w_307_123, w_307_166, w_307_305, w_307_343, w_307_350, w_307_391, w_307_415;
  wire w_308_008, w_308_022, w_308_026, w_308_034, w_308_064, w_308_067, w_308_095, w_308_107, w_308_115, w_308_123, w_308_126, w_308_146, w_308_147, w_308_155;
  wire w_309_034, w_309_187, w_309_193, w_309_215, w_309_264, w_309_270, w_309_301, w_309_352, w_309_380, w_309_382, w_309_383, w_309_384, w_309_385, w_309_386, w_309_387, w_309_388, w_309_389, w_309_390, w_309_391;
  wire w_310_061, w_310_071, w_310_093, w_310_145, w_310_165, w_310_188, w_310_244, w_310_251, w_310_258, w_310_365, w_310_412, w_310_447, w_310_496, w_310_557, w_310_582;
  wire w_311_003, w_311_080, w_311_123, w_311_131, w_311_134, w_311_180, w_311_245, w_311_256, w_311_263, w_311_288, w_311_325, w_311_369, w_311_439;
  wire w_312_023, w_312_040, w_312_042, w_312_056, w_312_060, w_312_133, w_312_146, w_312_238, w_312_355, w_312_363, w_312_432;
  wire w_313_008, w_313_030, w_313_080, w_313_083, w_313_090, w_313_118, w_313_128, w_313_149, w_313_192, w_313_231, w_313_240, w_313_254, w_313_258, w_313_397, w_313_403;
  wire w_314_014, w_314_032, w_314_077, w_314_092, w_314_134, w_314_159, w_314_174, w_314_191, w_314_204, w_314_219, w_314_220, w_314_221, w_314_225, w_314_226, w_314_227, w_314_228, w_314_229, w_314_230, w_314_231, w_314_232, w_314_234;
  wire w_315_111, w_315_140, w_315_171, w_315_238, w_315_269, w_315_362, w_315_523, w_315_524, w_315_530, w_315_634, w_315_665, w_315_724;
  wire w_316_066, w_316_072, w_316_149, w_316_219, w_316_246, w_316_257, w_316_410, w_316_450, w_316_453;
  wire w_317_014, w_317_090, w_317_148, w_317_162, w_317_249, w_317_261, w_317_264, w_317_298;
  wire w_318_000, w_318_003, w_318_004, w_318_011, w_318_012, w_318_013, w_318_014, w_318_015;
  wire w_319_077, w_319_129, w_319_200, w_319_210, w_319_218, w_319_278, w_319_289, w_319_347;
  wire w_320_004, w_320_019, w_320_123, w_320_178, w_320_218, w_320_224, w_320_285, w_320_297, w_320_309, w_320_318, w_320_369, w_320_389, w_320_411;
  wire w_321_001, w_321_005, w_321_063, w_321_141, w_321_176, w_321_282, w_321_303, w_321_536;
  wire w_322_001, w_322_002, w_322_005, w_322_008, w_322_013, w_322_014, w_322_015, w_322_017, w_322_022;
  wire w_323_061, w_323_089, w_323_123, w_323_139, w_323_230, w_323_269, w_323_284;
  wire w_324_008, w_324_011, w_324_012, w_324_029, w_324_031, w_324_035, w_324_045, w_324_052;
  wire w_325_000, w_325_005, w_325_035, w_325_046, w_325_139, w_325_238, w_325_272, w_325_310;
  wire w_326_031, w_326_035, w_326_042, w_326_043, w_326_077, w_326_104, w_326_111, w_326_113, w_326_114, w_326_179;
  wire w_327_097, w_327_155, w_327_344, w_327_363, w_327_364, w_327_438, w_327_440, w_327_444;
  wire w_328_004, w_328_010, w_328_026, w_328_037, w_328_053, w_328_110, w_328_120, w_328_153;
  wire w_329_037, w_329_039, w_329_094, w_329_306, w_329_384;
  wire w_330_016, w_330_035, w_330_042, w_330_059, w_330_116, w_330_201, w_330_247, w_330_279;
  wire w_331_025, w_331_052, w_331_072, w_331_111, w_331_153, w_331_247, w_331_255, w_331_315, w_331_330, w_331_439, w_331_507, w_331_508, w_331_509, w_331_510, w_331_511, w_331_512, w_331_513, w_331_514, w_331_515, w_331_519, w_331_520, w_331_521, w_331_522, w_331_523, w_331_524, w_331_525, w_331_527;
  wire w_332_004, w_332_142, w_332_224, w_332_261, w_332_363, w_332_409, w_332_451, w_332_668, w_332_669, w_332_670, w_332_671, w_332_672, w_332_673, w_332_674, w_332_675;
  wire w_333_011, w_333_115, w_333_137, w_333_158, w_333_222, w_333_223, w_333_314;
  wire w_334_098, w_334_139, w_334_337, w_334_340, w_334_367, w_334_368, w_334_486, w_334_640;
  wire w_335_033, w_335_041, w_335_098, w_335_102, w_335_116, w_335_134, w_335_151, w_335_162;
  wire w_336_002, w_336_016, w_336_025, w_336_029, w_336_057, w_336_074, w_336_083, w_336_110, w_336_124, w_336_140, w_336_177, w_336_209, w_336_235;
  wire w_337_004, w_337_020, w_337_028, w_337_036, w_337_072, w_337_101, w_337_188, w_337_225, w_337_356, w_337_384, w_337_412;
  wire w_338_003, w_338_010, w_338_022, w_338_028, w_338_044, w_338_049, w_338_094, w_338_158, w_338_239, w_338_264, w_338_312;
  wire w_339_003, w_339_008, w_339_012, w_339_019, w_339_020, w_339_022, w_339_028, w_339_029, w_339_039, w_339_041;
  wire w_340_000, w_340_004, w_340_010, w_340_011, w_340_013, w_340_026, w_340_030, w_340_038, w_340_046, w_340_049, w_340_050, w_340_051, w_340_052, w_340_053, w_340_054, w_340_055, w_340_056, w_340_057, w_340_058;
  wire w_341_035, w_341_245, w_341_351, w_341_408, w_341_418, w_341_458, w_341_487, w_341_599, w_341_704, w_341_774;
  wire w_342_047, w_342_103, w_342_111, w_342_194, w_342_213, w_342_217, w_342_311, w_342_344, w_342_358, w_342_477;
  wire w_343_138, w_343_246, w_343_251, w_343_335, w_343_360, w_343_425, w_343_478, w_343_479, w_343_580, w_343_605, w_343_697;
  wire w_344_001, w_344_026, w_344_042, w_344_061, w_344_063, w_344_077, w_344_088, w_344_116, w_344_148, w_344_263, w_344_455;
  wire w_345_013, w_345_017, w_345_053, w_345_098, w_345_129, w_345_216, w_345_250;
  wire w_346_076, w_346_104, w_346_139, w_346_565;
  wire w_347_016, w_347_021, w_347_036, w_347_053, w_347_098, w_347_109, w_347_117, w_347_167, w_347_252, w_347_257, w_347_268, w_347_328, w_347_331;
  wire w_348_101, w_348_114, w_348_137, w_348_213, w_348_243;
  wire w_349_027, w_349_028, w_349_036, w_349_060, w_349_089, w_349_177, w_349_214, w_349_230, w_349_289, w_349_305;
  wire w_350_022, w_350_049, w_350_071, w_350_094, w_350_123;
  wire w_351_044, w_351_049, w_351_051, w_351_070, w_351_075, w_351_095, w_351_106, w_351_228, w_351_235, w_351_240, w_351_336;
  wire w_352_047, w_352_296, w_352_314, w_352_411;
  wire w_353_047, w_353_106, w_353_137, w_353_189, w_353_244, w_353_311, w_353_443, w_353_535, w_353_570;
  wire w_354_003, w_354_004, w_354_010, w_354_039, w_354_048, w_354_082, w_354_112, w_354_113, w_354_207;
  wire w_355_038, w_355_051, w_355_071, w_355_072, w_355_079, w_355_100, w_355_113, w_355_192, w_355_295, w_355_297, w_355_405;
  wire w_356_001, w_356_003, w_356_039, w_356_043, w_356_044, w_356_048, w_356_061, w_356_078, w_356_108;
  wire w_357_005, w_357_096, w_357_296, w_357_302, w_357_304, w_357_318, w_357_319, w_357_381, w_357_408, w_357_460, w_357_588, w_357_658;
  wire w_358_066, w_358_227, w_358_284, w_358_295;
  wire w_359_015, w_359_021, w_359_041, w_359_047, w_359_051, w_359_074, w_359_075, w_359_089, w_359_090, w_359_154, w_359_170, w_359_176, w_359_198, w_359_209, w_359_210, w_359_211, w_359_212, w_359_213, w_359_214, w_359_215, w_359_216, w_359_217, w_359_221, w_359_222, w_359_223, w_359_224, w_359_225, w_359_227;
  wire w_360_021, w_360_150, w_360_266, w_360_269, w_360_288, w_360_315, w_360_353, w_360_373, w_360_383, w_360_414, w_360_419, w_360_429, w_360_482, w_360_520, w_360_521, w_360_522, w_360_523, w_360_524;
  wire w_361_031, w_361_070, w_361_097, w_361_104, w_361_200, w_361_221, w_361_249, w_361_354, w_361_369;
  wire w_362_013, w_362_019, w_362_031, w_362_104, w_362_193, w_362_283, w_362_337, w_362_420;
  wire w_363_009, w_363_056, w_363_057, w_363_123, w_363_359, w_363_372;
  wire w_364_009, w_364_013, w_364_027;
  wire w_365_045, w_365_106, w_365_128, w_365_196, w_365_199, w_365_252, w_365_390;
  wire w_366_013, w_366_072, w_366_144, w_366_174, w_366_238, w_366_313, w_366_358;
  wire w_367_035, w_367_075, w_367_123, w_367_125, w_367_160, w_367_221, w_367_295, w_367_491, w_367_654, w_367_755;
  wire w_368_015, w_368_022, w_368_024, w_368_029, w_368_066, w_368_067, w_368_081, w_368_084, w_368_111;
  wire w_369_115, w_369_133, w_369_282, w_369_524, w_369_666, w_369_722, w_369_740, w_369_741, w_369_742, w_369_743, w_369_744, w_369_745, w_369_747, w_369_749, w_369_750, w_369_751, w_369_752, w_369_753, w_369_754, w_369_755, w_369_757, w_369_759, w_369_760, w_369_761, w_369_762, w_369_763, w_369_765, w_369_767, w_369_768, w_369_769, w_369_770, w_369_771, w_369_772, w_369_773, w_369_775;
  wire w_370_020, w_370_031, w_370_051, w_370_056, w_370_065, w_370_084, w_370_095, w_370_099;
  wire w_371_000;
  wire w_372_000, w_372_003, w_372_008, w_372_031, w_372_033, w_372_038;
  wire w_373_001, w_373_013, w_373_057, w_373_092, w_373_241, w_373_268, w_373_327;
  wire w_374_056, w_374_076, w_374_091, w_374_141;
  wire w_375_032, w_375_071, w_375_142, w_375_171, w_375_178, w_375_190, w_375_191, w_375_192, w_375_193, w_375_194, w_375_195, w_375_196, w_375_197, w_375_198, w_375_199, w_375_200, w_375_204, w_375_205, w_375_206, w_375_207, w_375_208, w_375_209, w_375_210, w_375_211, w_375_212, w_375_214;
  wire w_376_055, w_376_070, w_376_138, w_376_176, w_376_251, w_376_275, w_376_277, w_376_278, w_376_279, w_376_280, w_376_281, w_376_282, w_376_283, w_376_284, w_376_285, w_376_286, w_376_290, w_376_291, w_376_292, w_376_293, w_376_295;
  wire w_377_013, w_377_040, w_377_065, w_377_066, w_377_087;
  wire w_378_022, w_378_046, w_378_107, w_378_111, w_378_112, w_378_119;
  wire w_379_071, w_379_085, w_379_099, w_379_103, w_379_182, w_379_186;
  wire w_380_035, w_380_162, w_380_284, w_380_296, w_380_317, w_380_615, w_380_731;
  wire w_381_038, w_381_104, w_381_163, w_381_284, w_381_319, w_381_653, w_381_670;
  wire w_382_033, w_382_046, w_382_341, w_382_477, w_382_563, w_382_615;
  wire w_383_018, w_383_031, w_383_092, w_383_112, w_383_240, w_383_350, w_383_394, w_383_450, w_383_455, w_383_591, w_383_618, w_383_733, w_383_734, w_383_735, w_383_736, w_383_737, w_383_738, w_383_739, w_383_741, w_383_743, w_383_744, w_383_745, w_383_746, w_383_747, w_383_748, w_383_749, w_383_753, w_383_754, w_383_755, w_383_756, w_383_758, w_383_760, w_383_761, w_383_762, w_383_763, w_383_764, w_383_765, w_383_766, w_383_767, w_383_768, w_383_769, w_383_770, w_383_771, w_383_773, w_383_775, w_383_776, w_383_777, w_383_778, w_383_779, w_383_780, w_383_782;
  wire w_384_042, w_384_046, w_384_121, w_384_149, w_384_162;
  wire w_385_007, w_385_089, w_385_106, w_385_124, w_385_213, w_385_227, w_385_427, w_385_429;
  wire w_386_015, w_386_041, w_386_080, w_386_115, w_386_146, w_386_152, w_386_161, w_386_188, w_386_226, w_386_473;
  wire w_387_012, w_387_219, w_387_252;
  wire w_388_012, w_388_025, w_388_057, w_388_076, w_388_090, w_388_100, w_388_159;
  wire w_389_066, w_389_087, w_389_150, w_389_234, w_389_279, w_389_308, w_389_437;
  wire w_390_031, w_390_054, w_390_138, w_390_148, w_390_173, w_390_187, w_390_252;
  wire w_391_100, w_391_105, w_391_249, w_391_463, w_391_491, w_391_610, w_391_670, w_391_738;
  wire w_392_081, w_392_083, w_392_185, w_392_244, w_392_245, w_392_262, w_392_552, w_392_553, w_392_554, w_392_555, w_392_556, w_392_560, w_392_561, w_392_562, w_392_563, w_392_564, w_392_565, w_392_566, w_392_567, w_392_568, w_392_569, w_392_570, w_392_572;
  wire w_393_003, w_393_016, w_393_020, w_393_050, w_393_084, w_393_102, w_393_109, w_393_113, w_393_129, w_393_136, w_393_149, w_393_194, w_393_204, w_393_239, w_393_240, w_393_241, w_393_242, w_393_243, w_393_244, w_393_245, w_393_246, w_393_250, w_393_251, w_393_252, w_393_253, w_393_254, w_393_255, w_393_256, w_393_257, w_393_258, w_393_259, w_393_260, w_393_262;
  wire w_394_040, w_394_070, w_394_080, w_394_107;
  wire w_395_029, w_395_041, w_395_072, w_395_080, w_395_229, w_395_235, w_395_290, w_395_372;
  wire w_396_004, w_396_007, w_396_025, w_396_045, w_396_065;
  wire w_397_018, w_397_019, w_397_036, w_397_046, w_397_048, w_397_050, w_397_060, w_397_064, w_397_081, w_397_092, w_397_137, w_397_141;
  wire w_398_023, w_398_029, w_398_043, w_398_050, w_398_058, w_398_061, w_398_067, w_398_074;
  wire w_399_023, w_399_035, w_399_098, w_399_118, w_399_137, w_399_163, w_399_285, w_399_297;
  wire w_400_009, w_400_024, w_400_051, w_400_091;
  wire w_401_008, w_401_079, w_401_158, w_401_170, w_401_178, w_401_205, w_401_230, w_401_244, w_401_246;
  wire w_402_021, w_402_027, w_402_028, w_402_032, w_402_068, w_402_080, w_402_087, w_402_114, w_402_135;
  wire w_403_120, w_403_216, w_403_289, w_403_315, w_403_325, w_403_439;
  wire w_404_022, w_404_182, w_404_196, w_404_339, w_404_361, w_404_588, w_404_606, w_404_648;
  wire w_405_026, w_405_027, w_405_071, w_405_073, w_405_132, w_405_137, w_405_166, w_405_182;
  wire w_406_004, w_406_022, w_406_050, w_406_116, w_406_221, w_406_280, w_406_282;
  wire w_407_063, w_407_070, w_407_133, w_407_267, w_407_293, w_407_356, w_407_572, w_407_643;
  wire w_408_002, w_408_003, w_408_004, w_408_005;
  wire w_409_049, w_409_153, w_409_304, w_409_408, w_409_455;
  wire w_410_011, w_410_027, w_410_048, w_410_064, w_410_085, w_410_102, w_410_142;
  wire w_411_130, w_411_567, w_411_581;
  wire w_412_076, w_412_202, w_412_275, w_412_300, w_412_374, w_412_398;
  wire w_413_015, w_413_022, w_413_029, w_413_045, w_413_083;
  wire w_414_089, w_414_151, w_414_241, w_414_303, w_414_325;
  wire w_415_046, w_415_050, w_415_072, w_415_079, w_415_283;
  wire w_416_134, w_416_168, w_416_325, w_416_344, w_416_427;
  wire w_417_050, w_417_057, w_417_060, w_417_065, w_417_075, w_417_083, w_417_100, w_417_116, w_417_120, w_417_137;
  wire w_418_029, w_418_045, w_418_048, w_418_052, w_418_068, w_418_091, w_418_105;
  wire w_419_044, w_419_139, w_419_155, w_419_240, w_419_308, w_419_324, w_419_325, w_419_326, w_419_327, w_419_328, w_419_332, w_419_333, w_419_334, w_419_336;
  wire w_420_161, w_420_483, w_420_519, w_420_574, w_420_587, w_420_607, w_420_673;
  wire w_421_047, w_421_052, w_421_075, w_421_126, w_421_243;
  wire w_422_001, w_422_002, w_422_005, w_422_007, w_422_008, w_422_010, w_422_013;
  wire w_423_019, w_423_021, w_423_022, w_423_038, w_423_052, w_423_057, w_423_073, w_423_075, w_423_092;
  wire w_424_087, w_424_111, w_424_156, w_424_222, w_424_228;
  wire w_425_000, w_425_102, w_425_214, w_425_247, w_425_358, w_425_362, w_425_551, w_425_552, w_425_553, w_425_554, w_425_555, w_425_556, w_425_557, w_425_558, w_425_562, w_425_563, w_425_564, w_425_565, w_425_567;
  wire w_426_017, w_426_022, w_426_162;
  wire w_427_050, w_427_051, w_427_053, w_427_059;
  wire w_428_010, w_428_124, w_428_181;
  wire w_429_003, w_429_085, w_429_096, w_429_115, w_429_130, w_429_137, w_429_218, w_429_236, w_429_259;
  wire w_430_060, w_430_092, w_430_114, w_430_286, w_430_422, w_430_484, w_430_534;
  wire w_431_210;
  wire w_432_051, w_432_053, w_432_120, w_432_136, w_432_218, w_432_288, w_432_300, w_432_307, w_432_313;
  wire w_433_054, w_433_120, w_433_180, w_433_213, w_433_268, w_433_398, w_433_409, w_433_444;
  wire w_434_061, w_434_098, w_434_335, w_434_382, w_434_495;
  wire w_435_075, w_435_085, w_435_136, w_435_156;
  wire w_436_218, w_436_224, w_436_410, w_436_562, w_436_564;
  wire w_437_010, w_437_429;
  wire w_438_084, w_438_253, w_438_273;
  wire w_439_038, w_439_039, w_439_045, w_439_116, w_439_295, w_439_313;
  wire w_440_032, w_440_037, w_440_040, w_440_057, w_440_064, w_440_079;
  wire w_441_007, w_441_023, w_441_144, w_441_407, w_441_505;
  wire w_442_045, w_442_104, w_442_123, w_442_126, w_442_135, w_442_142, w_442_143, w_442_144, w_442_145, w_442_149, w_442_150, w_442_151, w_442_152, w_442_153, w_442_154, w_442_155, w_442_156, w_442_157, w_442_158, w_442_159, w_442_161;
  wire w_443_130, w_443_263, w_443_327;
  wire w_444_022, w_444_101, w_444_165, w_444_307, w_444_425, w_444_462, w_444_520, w_444_585, w_444_709;
  wire w_445_012, w_445_021, w_445_025, w_445_029, w_445_069, w_445_135, w_445_182, w_445_183, w_445_184, w_445_185, w_445_186, w_445_187, w_445_188, w_445_189, w_445_190, w_445_191, w_445_192, w_445_196, w_445_197, w_445_198, w_445_199, w_445_200, w_445_201, w_445_202, w_445_203, w_445_204, w_445_205, w_445_206, w_445_207, w_445_211, w_445_212, w_445_213, w_445_214, w_445_215;
  wire w_446_025, w_446_151, w_446_152, w_446_242, w_446_298, w_446_406, w_446_438, w_446_533, w_446_544, w_446_577;
  wire w_447_093, w_447_099, w_447_125, w_447_160, w_447_173, w_447_336, w_447_338;
  wire w_448_104, w_448_117, w_448_151, w_448_161, w_448_245, w_448_260, w_448_264, w_448_283;
  wire w_449_138, w_449_218, w_449_261;
  wire w_450_029, w_450_052, w_450_067, w_450_070, w_450_103, w_450_104, w_450_107, w_450_175;
  wire w_451_006, w_451_064, w_451_105, w_451_133, w_451_217, w_451_240;
  wire w_452_045, w_452_112, w_452_125, w_452_300, w_452_341;
  wire w_453_090, w_453_552;
  wire w_454_025, w_454_039, w_454_064, w_454_073, w_454_079, w_454_085, w_454_111, w_454_119, w_454_158, w_454_305, w_454_340;
  wire w_455_026, w_455_112, w_455_144, w_455_172, w_455_205, w_455_418;
  wire w_456_039, w_456_127, w_456_193;
  wire w_457_002, w_457_053, w_457_054, w_457_089, w_457_099, w_457_107, w_457_132, w_457_139, w_457_154, w_457_164;
  wire w_458_038, w_458_060, w_458_072;
  wire w_459_035, w_459_109, w_459_216;
  wire w_460_003, w_460_040, w_460_089, w_460_173, w_460_233, w_460_237;
  wire w_461_173, w_461_637;
  wire w_462_016, w_462_379, w_462_400, w_462_524, w_462_547;
  wire w_463_000, w_463_029, w_463_119, w_463_192;
  wire w_464_118, w_464_242, w_464_281, w_464_299, w_464_668, w_464_676;
  wire w_465_014, w_465_019, w_465_165, w_465_192, w_465_208, w_465_224, w_465_269, w_465_332;
  wire w_466_053, w_466_066, w_466_103, w_466_136, w_466_214, w_466_296;
  wire w_467_167, w_467_177, w_467_181, w_467_251, w_467_284, w_467_367;
  wire w_468_021, w_468_025, w_468_035, w_468_062, w_468_070, w_468_079, w_468_090, w_468_105, w_468_137, w_468_154;
  wire w_469_024, w_469_062, w_469_069, w_469_080;
  wire w_470_407, w_470_504;
  wire w_471_074, w_471_169, w_471_190;
  wire w_472_163;
  wire w_473_502;
  wire w_474_160, w_474_202, w_474_307;
  wire w_475_011, w_475_057, w_475_190, w_475_193, w_475_293, w_475_296, w_475_511;
  wire w_476_235, w_476_274, w_476_513;
  wire w_477_022, w_477_030, w_477_032, w_477_034, w_477_041, w_477_057, w_477_070;
  wire w_478_078, w_478_177, w_478_275, w_478_335, w_478_381;
  wire w_479_034, w_479_072, w_479_088, w_479_107, w_479_169, w_479_185, w_479_281, w_479_314, w_479_325;
  wire w_480_029, w_480_046, w_480_057, w_480_075, w_480_078, w_480_102, w_480_107;
  wire w_481_039, w_481_042, w_481_050, w_481_054, w_481_057, w_481_058, w_481_104, w_481_198, w_481_215, w_481_280;
  wire w_482_003, w_482_077, w_482_175, w_482_287, w_482_327, w_482_434;
  wire w_483_358, w_483_428, w_483_777;
  wire w_484_008, w_484_249, w_484_277, w_484_296, w_484_326, w_484_329, w_484_346, w_484_349, w_484_379;
  wire w_485_072, w_485_143;
  wire w_486_038, w_486_111;
  wire w_487_002, w_487_101, w_487_127, w_487_141, w_487_319, w_487_510;
  wire w_488_017, w_488_018, w_488_021, w_488_037, w_488_045, w_488_102;
  wire w_489_025, w_489_094, w_489_384, w_489_395;
  wire w_490_012, w_490_019, w_490_067, w_490_089, w_490_093;
  wire w_491_021, w_491_022, w_491_040, w_491_077;
  wire w_492_157, w_492_275, w_492_319, w_492_323;
  wire w_493_026, w_493_038, w_493_044, w_493_050, w_493_093, w_493_095, w_493_103, w_493_139;
  wire w_494_028, w_494_046, w_494_241;
  wire w_495_026, w_495_096, w_495_128, w_495_164, w_495_183, w_495_343, w_495_435;
  wire w_496_077, w_496_447, w_496_599, w_496_600, w_496_601, w_496_602, w_496_603, w_496_604;
  wire w_497_078, w_497_107;
  wire w_498_120, w_498_170, w_498_415, w_498_619;
  wire w_499_189, w_499_222, w_499_376, w_499_433, w_499_548, w_499_573, w_499_583;
  wire w_500_020, w_500_064, w_500_175, w_500_203, w_500_226, w_500_274, w_500_302, w_500_353;
  wire w_501_013, w_501_030;
  wire w_502_349, w_502_372, w_502_416, w_502_472, w_502_539, w_502_662, w_502_663, w_502_664, w_502_665, w_502_666, w_502_667, w_502_671, w_502_672, w_502_673, w_502_674, w_502_675, w_502_676, w_502_677, w_502_678, w_502_679, w_502_680, w_502_682, w_502_684, w_502_685, w_502_686, w_502_687, w_502_688, w_502_689, w_502_690, w_502_691, w_502_692, w_502_696, w_502_697, w_502_698, w_502_699, w_502_700, w_502_701, w_502_703;
  wire w_503_015, w_503_190, w_503_202, w_503_252, w_503_483, w_503_484, w_503_485, w_503_486, w_503_487, w_503_488, w_503_489, w_503_490, w_503_491, w_503_492;
  wire w_504_027, w_504_031, w_504_053;
  wire w_505_066, w_505_074, w_505_236;
  wire w_506_071, w_506_153, w_506_261, w_506_513, w_506_594, w_506_611, w_506_632, w_506_633, w_506_634, w_506_638, w_506_639, w_506_640, w_506_641, w_506_642, w_506_644;
  wire w_507_012, w_507_016, w_507_035, w_507_046;
  wire w_508_005, w_508_074, w_508_172, w_508_173, w_508_396;
  wire w_509_075, w_509_087, w_509_088, w_509_089, w_509_090, w_509_091, w_509_092, w_509_096, w_509_097, w_509_098, w_509_099, w_509_100, w_509_101, w_509_102, w_509_104;
  wire w_510_136, w_510_292, w_510_447, w_510_595, w_510_748;
  wire w_511_028, w_511_186, w_511_240, w_511_326, w_511_396;
  wire w_512_059, w_512_088, w_512_098, w_512_124, w_512_157, w_512_434, w_512_451;
  wire w_513_076, w_513_232, w_513_378, w_513_448, w_513_499, w_513_576;
  wire w_514_083, w_514_170, w_514_191, w_514_456;
  wire w_515_066, w_515_094, w_515_172, w_515_371;
  wire w_516_079, w_516_096, w_516_329, w_516_406;
  wire w_517_005, w_517_052, w_517_098, w_517_227;
  wire w_518_010, w_518_057, w_518_062;
  wire w_519_022, w_519_041;
  wire w_520_053, w_520_109, w_520_202, w_520_253, w_520_293, w_520_294, w_520_295, w_520_299, w_520_300, w_520_301, w_520_302, w_520_303, w_520_305;
  wire w_521_058, w_521_151, w_521_322, w_521_334;
  wire w_522_092, w_522_256, w_522_397, w_522_505, w_522_539;
  wire w_523_003, w_523_065, w_523_087, w_523_190, w_523_473;
  wire w_524_346, w_524_444, w_524_591, w_524_595, w_524_612;
  wire w_525_007, w_525_029, w_525_081, w_525_095;
  wire w_526_153;
  wire w_527_061, w_527_082, w_527_096, w_527_197, w_527_223, w_527_350, w_527_526;
  wire w_528_015, w_528_017, w_528_039, w_528_046;
  wire w_529_000, w_529_002, w_529_004;
  wire w_530_042, w_530_096, w_530_147, w_530_182, w_530_219;
  wire w_531_012, w_531_317, w_531_580;
  wire w_532_176, w_532_222, w_532_243, w_532_244, w_532_245, w_532_246, w_532_247, w_532_248, w_532_249, w_532_250, w_532_251, w_532_252, w_532_253, w_532_254, w_532_258, w_532_259, w_532_260, w_532_261, w_532_262, w_532_263, w_532_264, w_532_266;
  wire w_533_089, w_533_110, w_533_169, w_533_187, w_533_253, w_533_329, w_533_361, w_533_532, w_533_550;
  wire w_534_003, w_534_011, w_534_017, w_534_018, w_534_019, w_534_020, w_534_021, w_534_022, w_534_023, w_534_024;
  wire w_535_000, w_535_114, w_535_119, w_535_180, w_535_189, w_535_202, w_535_252, w_535_262, w_535_263, w_535_264, w_535_265, w_535_266, w_535_267, w_535_268, w_535_269, w_535_273, w_535_274, w_535_275, w_535_276, w_535_278, w_535_280, w_535_281, w_535_282, w_535_283, w_535_284, w_535_285, w_535_286, w_535_287, w_535_288, w_535_292, w_535_293, w_535_294, w_535_295, w_535_296, w_535_297, w_535_299;
  wire w_536_022, w_536_040;
  wire w_537_029, w_537_032, w_537_053, w_537_056, w_537_154, w_537_220, w_537_248, w_537_264;
  wire w_538_039, w_538_046, w_538_190, w_538_262;
  wire w_539_321, w_539_387, w_539_388, w_539_422, w_539_491, w_539_538, w_539_723;
  wire w_540_053, w_540_118;
  wire w_541_024, w_541_066;
  wire w_542_007, w_542_053, w_542_058, w_542_061, w_542_116, w_542_331;
  wire w_543_105, w_543_210, w_543_770, w_543_771, w_543_772, w_543_773, w_543_774, w_543_775, w_543_776, w_543_777, w_543_778, w_543_779, w_543_780, w_543_784, w_543_785, w_543_786, w_543_788;
  wire w_544_146, w_544_153;
  wire w_545_117, w_545_151, w_545_345, w_545_349;
  wire w_546_073, w_546_086, w_546_385, w_546_450, w_546_518, w_546_519, w_546_520, w_546_521, w_546_522, w_546_523, w_546_524;
  wire w_547_002, w_547_024, w_547_031, w_547_032, w_547_034, w_547_035, w_547_045;
  wire w_548_060, w_548_192, w_548_264;
  wire w_549_047, w_549_107, w_549_130;
  wire w_550_122, w_550_260;
  wire w_551_007, w_551_012, w_551_031, w_551_088, w_551_109;
  wire w_552_006, w_552_100, w_552_304;
  wire w_553_015, w_553_020, w_553_027, w_553_031;
  wire w_554_069;
  wire w_555_067, w_555_293;
  wire w_556_035, w_556_212, w_556_270, w_556_324, w_556_463;
  wire w_557_047, w_557_050, w_557_062, w_557_111, w_557_167, w_557_419, w_557_429, w_557_430, w_557_431, w_557_432;
  wire w_558_030, w_558_122, w_558_151;
  wire w_559_020, w_559_028, w_559_040;
  wire w_560_071, w_560_106, w_560_149, w_560_512, w_560_543;
  wire w_561_038, w_561_079, w_561_175, w_561_205, w_561_308, w_561_343;
  wire w_562_147, w_562_429, w_562_660;
  wire w_563_022, w_563_052, w_563_470;
  wire w_564_007, w_564_065, w_564_097, w_564_280, w_564_281, w_564_282, w_564_283, w_564_284, w_564_285, w_564_286, w_564_287, w_564_288, w_564_289, w_564_290, w_564_291;
  wire w_565_008, w_565_009, w_565_020;
  wire w_566_094, w_566_198;
  wire w_567_003, w_567_010, w_567_014, w_567_016, w_567_020, w_567_033, w_567_040, w_567_042;
  wire w_568_227, w_568_367, w_568_499;
  wire w_569_040, w_569_133;
  wire w_570_085, w_570_198, w_570_199, w_570_200, w_570_201, w_570_202, w_570_203, w_570_204, w_570_205, w_570_206, w_570_208, w_570_210, w_570_211, w_570_212, w_570_213, w_570_214, w_570_215, w_570_216, w_570_217, w_570_218, w_570_220;
  wire w_571_075, w_571_130, w_571_402;
  wire w_572_107, w_572_131, w_572_140;
  wire w_573_020, w_573_043, w_573_058, w_573_208, w_573_223, w_573_324;
  wire w_574_164, w_574_265, w_574_373;
  wire w_575_000, w_575_053, w_575_064, w_575_065, w_575_094, w_575_096, w_575_160, w_575_178, w_575_207;
  wire w_576_111, w_576_172, w_576_289, w_576_290, w_576_291, w_576_292, w_576_293, w_576_294, w_576_295, w_576_296, w_576_297, w_576_298;
  wire w_577_031, w_577_485, w_577_496;
  wire w_578_007, w_578_284, w_578_543, w_578_724;
  wire w_579_358, w_579_461, w_579_647;
  wire w_580_031, w_580_420;
  wire w_581_400;
  wire w_582_245, w_582_461, w_582_657, w_582_708;
  wire w_583_002, w_583_023, w_583_075, w_583_100, w_583_101, w_583_102, w_583_106, w_583_107, w_583_108, w_583_109, w_583_110, w_583_111, w_583_112, w_583_113, w_583_114, w_583_115, w_583_117;
  wire w_584_024, w_584_255, w_584_341, w_584_544, w_584_574, w_584_666, w_584_712;
  wire w_585_046, w_585_101, w_585_554, w_585_732, w_585_733, w_585_734, w_585_735, w_585_736, w_585_737, w_585_738, w_585_742, w_585_743, w_585_744, w_585_745, w_585_746, w_585_747, w_585_748, w_585_749, w_585_750, w_585_751, w_585_753, w_585_755, w_585_756, w_585_757, w_585_758, w_585_759, w_585_760, w_585_761, w_585_762, w_585_763, w_585_764, w_585_765, w_585_766;
  wire w_586_040, w_586_073, w_586_090, w_586_096, w_586_125, w_586_230, w_586_231, w_586_232, w_586_233, w_586_234, w_586_235, w_586_236;
  wire w_587_009, w_587_090, w_587_141, w_587_230, w_587_313;
  wire w_588_111, w_588_153, w_588_164;
  wire w_589_007, w_589_022, w_589_092, w_589_154, w_589_331;
  wire w_590_003, w_590_026, w_590_161;
  wire w_591_057, w_591_101, w_591_190, w_591_222, w_591_223, w_591_224, w_591_225, w_591_226, w_591_227, w_591_231, w_591_232, w_591_233, w_591_234, w_591_235, w_591_236, w_591_237, w_591_239;
  wire w_592_177, w_592_233, w_592_491;
  wire w_593_079, w_593_161;
  wire w_594_104, w_594_121;
  wire w_595_029, w_595_130, w_595_157, w_595_246;
  wire w_596_010, w_596_068, w_596_137, w_596_405;
  wire w_597_258;
  wire w_598_010, w_598_017, w_598_028;
  wire w_599_018, w_599_025, w_599_032;
  wire w_600_084, w_600_130, w_600_264, w_600_697;
  wire w_601_071, w_601_073, w_601_077, w_601_123, w_601_384, w_601_583;
  wire w_602_005, w_602_296;
  wire w_603_090, w_603_123, w_603_163, w_603_184, w_603_185, w_603_186, w_603_190, w_603_191, w_603_192, w_603_193, w_603_194, w_603_195, w_603_197;
  wire w_604_108, w_604_237;
  wire w_605_212, w_605_658;
  wire w_607_016;
  wire w_608_014, w_608_218, w_608_359, w_608_384;
  wire w_609_050, w_609_187, w_609_233;
  wire w_610_041, w_610_051, w_610_104;
  wire w_611_282, w_611_485;
  wire w_612_076, w_612_103;
  wire w_613_009, w_613_024, w_613_030, w_613_089;
  wire w_614_253, w_614_334;
  wire w_615_023, w_615_033, w_615_034, w_615_052, w_615_067, w_615_078, w_615_079;
  wire w_616_232, w_616_388;
  wire w_617_086, w_617_233;
  wire w_618_009, w_618_048, w_618_060;
  wire w_619_167, w_619_251, w_619_510;
  wire w_620_002, w_620_106, w_620_438, w_620_440;
  wire w_621_230, w_621_444;
  wire w_622_033, w_622_037, w_622_064, w_622_074;
  wire w_623_081, w_623_364;
  wire w_624_018, w_624_070;
  wire w_625_100, w_625_277;
  wire w_626_011, w_626_319, w_626_338, w_626_797, w_626_798, w_626_799, w_626_800, w_626_801, w_626_802, w_626_803, w_626_804, w_626_808, w_626_809, w_626_810, w_626_811, w_626_812, w_626_813, w_626_814, w_626_815, w_626_816, w_626_817, w_626_818, w_626_820, w_626_822, w_626_823, w_626_824, w_626_825, w_626_826, w_626_827, w_626_828, w_626_829, w_626_830, w_626_831, w_626_832, w_626_833;
  wire w_628_056, w_628_074, w_628_151;
  wire w_629_146, w_629_161, w_629_191, w_629_624;
  wire w_630_049, w_630_052;
  wire w_631_130, w_631_326;
  wire w_633_039, w_633_744;
  wire w_634_179, w_634_264, w_634_295;
  wire w_635_039, w_635_156, w_635_170, w_635_484;
  wire w_636_078, w_636_112, w_636_159;
  wire w_637_003, w_637_010, w_637_242;
  wire w_638_261, w_638_350, w_638_380, w_638_423, w_638_470;
  wire w_639_000, w_639_018;
  wire w_640_029, w_640_267, w_640_443, w_640_456, w_640_532, w_640_598, w_640_653;
  wire w_641_058, w_641_063, w_641_072;
  wire w_642_569;
  wire w_643_008, w_643_030, w_643_303;
  wire w_644_011;
  wire w_645_314;
  wire w_646_003, w_646_007, w_646_009, w_646_013;
  wire w_647_193, w_647_200, w_647_366, w_647_367, w_647_393, w_647_446, w_647_488;
  wire w_648_040, w_648_041, w_648_079;
  wire w_649_021, w_649_026, w_649_030, w_649_031, w_649_032, w_649_033, w_649_034, w_649_035, w_649_039, w_649_040, w_649_041, w_649_042, w_649_043, w_649_044, w_649_045, w_649_046, w_649_047, w_649_049;
  wire w_650_341, w_650_578, w_650_741;
  wire w_651_019, w_651_337, w_651_464;
  wire w_652_014, w_652_020, w_652_030, w_652_041, w_652_042, w_652_061;
  wire w_653_035, w_653_063, w_653_094, w_653_188, w_653_262;
  wire w_654_153, w_654_308, w_654_336, w_654_411, w_654_412, w_654_413, w_654_414, w_654_415, w_654_416, w_654_417;
  wire w_655_478;
  wire w_656_067, w_656_087, w_656_298, w_656_348, w_656_596, w_656_597, w_656_598, w_656_599, w_656_600, w_656_601, w_656_602, w_656_603, w_656_604, w_656_605, w_656_606, w_656_607;
  wire w_658_054, w_658_094, w_658_262;
  wire w_659_239;
  wire w_660_000, w_660_001;
  wire w_661_018, w_661_049;
  wire w_662_321;
  wire w_663_023, w_663_060, w_663_070, w_663_094;
  wire w_664_018, w_664_103, w_664_123, w_664_155;
  wire w_665_027, w_665_424;
  wire w_666_406, w_666_445;
  wire w_667_051, w_667_625;
  wire w_668_171;
  wire w_669_108, w_669_152, w_669_254, w_669_261, w_669_298, w_669_307;
  wire w_670_022, w_670_024, w_670_045;
  wire w_671_371;
  wire w_673_161, w_673_278, w_673_419;
  wire w_674_172, w_674_360;
  wire w_675_109, w_675_146, w_675_252, w_675_318;
  wire w_676_185, w_676_222, w_676_258;
  wire w_677_020, w_677_131;
  wire w_678_049, w_678_201, w_678_225, w_678_454;
  wire w_679_286, w_679_443, w_679_618;
  wire w_680_105, w_680_186;
  wire w_681_081, w_681_252, w_681_320;
  wire w_682_371, w_682_399, w_682_472, w_682_543, w_682_716, w_682_717, w_682_718, w_682_722, w_682_723, w_682_724, w_682_725, w_682_726, w_682_727, w_682_728, w_682_729, w_682_730, w_682_732;
  wire w_683_089, w_683_112, w_683_230, w_683_259;
  wire w_685_294, w_685_299;
  wire w_686_011, w_686_026, w_686_102, w_686_107;
  wire w_687_198;
  wire w_688_036, w_688_387, w_688_501, w_688_749, w_688_750, w_688_751, w_688_752, w_688_753, w_688_754, w_688_755, w_688_756, w_688_757, w_688_761, w_688_762, w_688_763, w_688_764, w_688_765, w_688_766, w_688_767, w_688_768, w_688_770;
  wire w_689_090, w_689_226, w_689_227, w_689_233, w_689_234, w_689_235, w_689_236, w_689_237, w_689_238, w_689_239, w_689_240, w_689_241;
  wire w_690_025, w_690_052, w_690_053, w_690_054, w_690_055, w_690_056;
  wire w_691_005, w_691_139;
  wire w_692_155, w_692_168;
  wire w_693_031, w_693_163, w_693_193, w_693_292, w_693_319, w_693_324;
  wire w_694_002, w_694_018, w_694_021, w_694_029;
  wire w_695_052, w_695_313, w_695_314, w_695_315, w_695_316, w_695_320, w_695_321, w_695_322, w_695_323, w_695_325;
  wire w_696_115;
  wire w_697_033, w_697_187, w_697_213;
  wire w_699_036, w_699_231, w_699_724;
  wire w_701_033, w_701_054, w_701_157;
  wire w_702_148;
  wire w_703_135, w_703_220, w_703_306;
  wire w_704_043, w_704_140, w_704_722, w_704_723, w_704_724, w_704_725, w_704_726, w_704_727, w_704_728, w_704_729, w_704_730, w_704_731, w_704_732;
  wire w_705_454, w_705_455, w_705_456, w_705_457, w_705_458, w_705_459, w_705_460, w_705_461, w_705_462, w_705_463;
  wire w_706_205, w_706_227;
  wire w_707_117, w_707_118;
  wire w_708_064, w_708_269;
  wire w_709_559;
  wire w_710_119;
  wire w_711_004, w_711_018, w_711_030, w_711_048, w_711_051, w_711_052, w_711_053, w_711_054, w_711_058, w_711_059, w_711_060, w_711_061, w_711_062, w_711_063, w_711_064, w_711_065, w_711_067;
  wire w_712_033, w_712_065;
  wire w_714_000, w_714_009, w_714_021, w_714_046;
  wire w_716_018, w_716_029;
  wire w_717_116;
  wire w_718_123, w_718_200, w_718_258, w_718_277, w_718_646;
  wire w_719_004, w_719_150, w_719_250, w_719_393;
  wire w_721_517;
  wire w_722_415;
  wire w_723_559, w_723_597;
  wire w_724_311, w_724_391, w_724_451;
  wire w_725_058, w_725_102, w_725_342;
  wire w_726_165, w_726_379, w_726_437;
  wire w_727_106;
  wire w_728_136, w_728_394, w_728_548, w_728_789, w_728_790, w_728_791, w_728_792, w_728_793, w_728_794, w_728_795, w_728_796, w_728_797;
  wire w_729_360;
  wire w_730_122, w_730_150, w_730_159, w_730_160, w_730_161, w_730_162, w_730_163, w_730_164, w_730_165, w_730_166, w_730_167, w_730_168, w_730_169;
  wire w_731_077, w_731_087, w_731_103, w_731_119, w_731_122, w_731_147, w_731_181, w_731_186, w_731_200, w_731_201, w_731_202, w_731_203, w_731_207, w_731_208, w_731_209, w_731_210, w_731_211, w_731_212, w_731_213, w_731_214, w_731_216;
  wire w_732_016;
  wire w_733_045, w_733_100, w_733_108;
  wire w_734_086, w_734_104;
  wire w_735_051;
  wire w_736_059, w_736_091, w_736_389;
  wire w_737_012, w_737_115, w_737_621, w_737_622, w_737_623, w_737_624, w_737_625, w_737_626, w_737_630, w_737_631, w_737_632, w_737_633, w_737_634, w_737_636;
  wire w_739_093, w_739_105;
  wire w_740_115, w_740_318;
  wire w_741_144;
  wire w_742_030;
  wire w_743_021, w_743_031, w_743_118, w_743_119, w_743_120, w_743_121, w_743_122, w_743_123, w_743_124, w_743_125, w_743_126, w_743_127, w_743_128, w_743_129, w_743_133, w_743_134, w_743_135, w_743_136, w_743_138;
  wire w_744_058, w_744_072;
  wire w_746_141, w_746_634, w_746_635, w_746_636, w_746_637, w_746_638, w_746_639, w_746_640, w_746_641, w_746_642;
  wire w_747_019;
  wire w_748_126, w_748_161, w_748_267;
  wire w_749_059, w_749_131, w_749_176;
  wire w_750_434, w_750_448;
  wire w_751_282, w_751_314, w_751_322;
  wire w_752_418;
  wire w_753_377, w_753_543;
  wire w_754_136, w_754_167;
  wire w_755_016;
  wire w_756_003, w_756_070, w_756_072, w_756_472, w_756_473, w_756_474, w_756_475, w_756_476;
  wire w_757_133;
  wire w_758_227;
  wire w_759_047, w_759_108, w_759_124, w_759_642, w_759_649;
  wire w_761_018, w_761_022;
  wire w_762_061, w_762_123, w_762_253;
  wire w_764_054, w_764_241, w_764_380, w_764_381, w_764_382, w_764_383, w_764_384, w_764_385, w_764_386, w_764_387, w_764_388;
  wire w_765_198;
  wire w_766_300, w_766_316, w_766_317, w_766_318, w_766_319, w_766_320, w_766_321, w_766_322, w_766_323, w_766_324, w_766_325, w_766_326, w_766_327, w_766_331, w_766_332, w_766_333, w_766_334, w_766_335, w_766_336, w_766_337, w_766_338, w_766_339, w_766_340, w_766_341, w_766_342, w_766_344;
  wire w_767_284;
  wire w_768_276, w_768_277, w_768_278, w_768_279, w_768_280, w_768_281, w_768_282, w_768_283, w_768_284, w_768_285, w_768_286, w_768_287, w_768_291, w_768_292, w_768_293, w_768_294, w_768_296;
  wire w_770_055, w_770_072;
  wire w_772_073, w_772_265, w_772_266, w_772_267, w_772_268, w_772_269, w_772_270, w_772_271, w_772_272, w_772_273, w_772_274, w_772_278, w_772_279, w_772_280, w_772_281, w_772_283;
  wire w_773_230, w_773_231, w_773_232, w_773_233, w_773_234, w_773_235, w_773_236;
  wire w_774_008;
  wire w_775_193;
  wire w_776_012, w_776_102;
  wire w_777_101;
  wire w_778_006;
  wire w_779_209, w_779_213;
  wire w_780_023;
  wire w_781_000;
  wire w_782_041, w_782_320;
  wire w_783_159, w_783_184, w_783_235;
  wire w_784_109, w_784_272, w_784_375, w_784_523, w_784_524, w_784_525, w_784_529, w_784_530, w_784_531, w_784_532, w_784_534, w_784_536, w_784_537, w_784_538, w_784_539, w_784_540, w_784_541, w_784_542, w_784_543, w_784_544, w_784_545, w_784_546, w_784_547;
  wire w_785_011;
  wire w_786_008, w_786_009;
  wire w_787_032;
  wire w_788_008, w_788_021, w_788_095, w_788_134, w_788_145;
  wire w_789_050, w_789_143, w_789_340;
  wire w_790_120, w_790_123, w_790_297, w_790_401;
  wire w_791_006;
  wire w_792_343;
  wire w_793_014, w_793_040, w_793_053;
  wire w_794_102;
  wire w_795_180;
  wire w_797_003;
  wire w_799_000;
  wire w_800_000, w_800_001, w_800_002, w_800_003, w_800_004, w_800_005, w_800_006, w_800_007, w_800_008, w_800_009, w_800_010, w_800_011, w_800_012, w_800_013, w_800_014, w_800_015, w_800_016, w_800_017, w_800_018, w_800_019, w_800_020, w_800_021, w_800_022, w_800_023, w_800_024, w_800_025, w_800_026, w_800_027, w_800_028, w_800_029, w_800_030, w_800_031, w_800_032, w_800_033, w_800_034, w_800_035, w_800_036, w_800_037, w_800_038, w_800_039, w_800_040, w_800_041, w_800_042, w_800_043, w_800_044, w_800_045, w_800_046, w_800_047, w_800_048, w_800_049, w_800_050, w_800_051, w_800_052, w_800_053, w_800_054, w_800_055, w_800_056, w_800_057, w_800_058, w_800_059, w_800_060, w_800_061, w_800_062, w_800_063, w_800_064, w_800_065, w_800_066, w_800_067, w_800_068, w_800_069, w_800_070, w_800_071, w_800_072, w_800_073, w_800_074, w_800_075, w_800_076, w_800_077, w_800_078, w_800_079, w_800_080, w_800_081, w_800_082, w_800_083, w_800_084, w_800_085, w_800_086, w_800_087, w_800_088, w_800_089, w_800_090, w_800_091, w_800_092, w_800_093, w_800_094, w_800_095, w_800_096, w_800_097, w_800_098, w_800_099, w_800_100, w_800_101, w_800_102, w_800_103, w_800_104, w_800_105, w_800_106, w_800_107, w_800_108, w_800_109, w_800_110, w_800_111, w_800_112, w_800_113, w_800_114, w_800_115, w_800_116, w_800_117, w_800_118, w_800_119, w_800_120, w_800_121, w_800_122, w_800_123, w_800_124, w_800_125, w_800_126, w_800_127, w_800_128, w_800_129, w_800_130, w_800_131, w_800_132, w_800_133, w_800_134, w_800_135, w_800_136, w_800_137, w_800_138, w_800_139, w_800_140, w_800_141, w_800_142, w_800_143, w_800_144, w_800_145, w_800_146, w_800_147, w_800_148, w_800_149, w_800_150, w_800_151, w_800_152, w_800_153, w_800_154, w_800_155, w_800_156, w_800_157, w_800_158, w_800_159, w_800_160, w_800_161, w_800_162, w_800_163, w_800_164, w_800_165, w_800_166, w_800_167, w_800_168, w_800_169, w_800_170, w_800_171, w_800_172, w_800_173, w_800_174, w_800_175, w_800_176, w_800_177, w_800_178, w_800_179, w_800_180, w_800_181, w_800_182, w_800_183, w_800_184, w_800_185, w_800_186, w_800_187, w_800_188, w_800_189, w_800_190, w_800_191, w_800_192, w_800_193, w_800_194, w_800_195, w_800_196, w_800_197, w_800_198, w_800_199, w_800_200, w_800_201, w_800_202, w_800_203, w_800_204, w_800_205, w_800_206, w_800_207, w_800_208, w_800_209, w_800_210, w_800_211, w_800_212, w_800_213, w_800_214, w_800_215, w_800_216, w_800_217, w_800_218, w_800_219, w_800_220, w_800_221, w_800_222, w_800_223, w_800_224, w_800_225, w_800_226, w_800_227, w_800_228, w_800_229, w_800_230, w_800_231, w_800_232, w_800_233, w_800_234, w_800_235, w_800_236, w_800_237, w_800_238, w_800_239, w_800_240, w_800_241, w_800_242, w_800_243, w_800_244, w_800_245, w_800_246, w_800_247, w_800_248, w_800_249, w_800_250, w_800_251, w_800_252, w_800_253, w_800_254, w_800_255, w_800_256, w_800_257, w_800_258, w_800_259, w_800_260, w_800_261, w_800_262, w_800_263, w_800_264, w_800_265, w_800_266, w_800_267, w_800_268, w_800_269, w_800_270, w_800_271, w_800_272, w_800_273, w_800_274, w_800_275, w_800_276, w_800_277, w_800_278, w_800_279, w_800_280, w_800_281, w_800_282, w_800_283, w_800_284, w_800_285, w_800_286, w_800_287, w_800_288, w_800_289, w_800_290, w_800_291, w_800_292, w_800_293, w_800_294, w_800_295, w_800_296, w_800_297, w_800_298, w_800_299, w_800_300, w_800_301, w_800_302, w_800_303, w_800_304, w_800_305, w_800_306, w_800_307, w_800_308, w_800_309, w_800_310, w_800_311, w_800_312, w_800_313, w_800_314, w_800_315, w_800_316, w_800_317, w_800_318, w_800_319, w_800_320, w_800_321, w_800_322, w_800_323, w_800_324, w_800_325, w_800_326, w_800_327, w_800_328, w_800_329, w_800_330, w_800_331, w_800_332, w_800_333, w_800_334, w_800_335, w_800_336, w_800_337, w_800_338, w_800_339, w_800_340, w_800_341, w_800_342, w_800_343, w_800_344, w_800_345, w_800_346, w_800_347, w_800_348, w_800_349, w_800_350, w_800_351, w_800_352, w_800_353, w_800_354, w_800_355, w_800_356, w_800_357, w_800_358, w_800_359, w_800_360, w_800_361, w_800_362, w_800_363, w_800_364, w_800_365, w_800_366, w_800_367, w_800_368, w_800_369, w_800_370, w_800_371, w_800_372, w_800_373, w_800_374, w_800_375, w_800_376, w_800_377, w_800_378, w_800_379, w_800_380, w_800_381, w_800_382, w_800_383, w_800_384, w_800_385, w_800_386, w_800_387, w_800_388, w_800_389, w_800_390, w_800_391, w_800_392, w_800_393, w_800_394, w_800_395, w_800_396, w_800_397, w_800_398, w_800_399, w_800_400, w_800_401, w_800_402, w_800_403, w_800_404, w_800_405, w_800_406, w_800_407, w_800_408, w_800_409, w_800_410, w_800_411, w_800_412, w_800_413, w_800_414, w_800_415, w_800_416, w_800_417, w_800_418, w_800_419, w_800_420, w_800_421, w_800_422, w_800_423, w_800_424, w_800_425, w_800_426, w_800_427, w_800_428, w_800_429, w_800_430, w_800_431, w_800_432, w_800_433, w_800_434, w_800_435, w_800_436, w_800_437, w_800_438, w_800_439, w_800_440, w_800_441, w_800_442, w_800_443, w_800_444, w_800_445, w_800_446, w_800_447, w_800_448, w_800_449, w_800_450, w_800_451, w_800_452, w_800_453, w_800_454, w_800_455, w_800_456, w_800_457, w_800_458, w_800_459, w_800_460, w_800_461, w_800_462, w_800_463, w_800_464, w_800_465, w_800_466, w_800_467, w_800_468, w_800_469, w_800_470, w_800_471, w_800_472, w_800_473, w_800_474, w_800_475, w_800_476, w_800_477, w_800_478, w_800_479, w_800_480, w_800_481, w_800_482, w_800_483, w_800_484, w_800_485, w_800_486, w_800_487, w_800_488, w_800_489, w_800_490, w_800_491, w_800_492, w_800_493, w_800_494, w_800_495, w_800_496, w_800_497, w_800_498, w_800_499, w_800_500, w_800_501, w_800_502, w_800_503, w_800_504, w_800_505, w_800_506, w_800_507, w_800_508, w_800_509, w_800_510, w_800_511, w_800_512, w_800_513, w_800_514, w_800_515, w_800_516, w_800_517, w_800_518, w_800_519, w_800_520, w_800_521, w_800_522, w_800_523, w_800_524, w_800_525, w_800_526, w_800_527, w_800_528, w_800_529, w_800_530, w_800_531, w_800_532, w_800_533, w_800_534, w_800_535, w_800_536, w_800_537, w_800_538, w_800_539, w_800_540, w_800_541, w_800_542, w_800_543, w_800_544, w_800_545, w_800_546, w_800_547, w_800_548, w_800_549, w_800_550, w_800_551, w_800_552, w_800_553, w_800_554, w_800_555, w_800_556, w_800_557, w_800_558, w_800_559, w_800_560, w_800_561, w_800_562, w_800_563, w_800_564, w_800_565, w_800_566, w_800_567, w_800_568, w_800_569, w_800_570, w_800_571, w_800_572, w_800_573, w_800_574, w_800_575, w_800_576, w_800_577, w_800_578, w_800_579, w_800_580, w_800_581, w_800_582, w_800_583, w_800_584, w_800_585, w_800_586, w_800_587, w_800_588, w_800_589, w_800_590, w_800_591, w_800_592, w_800_593, w_800_594, w_800_595, w_800_596, w_800_597, w_800_598, w_800_599, w_800_600, w_800_601, w_800_602, w_800_603, w_800_604, w_800_605, w_800_606, w_800_607, w_800_608, w_800_609, w_800_610, w_800_611, w_800_612, w_800_613, w_800_614, w_800_615, w_800_616, w_800_617, w_800_618, w_800_619, w_800_620, w_800_621, w_800_622, w_800_623, w_800_624, w_800_625, w_800_626, w_800_627, w_800_628, w_800_629, w_800_630, w_800_631, w_800_632, w_800_633, w_800_634, w_800_635, w_800_636, w_800_637, w_800_638, w_800_639, w_800_640, w_800_641, w_800_642, w_800_643, w_800_644, w_800_645, w_800_646, w_800_647, w_800_648, w_800_649, w_800_650, w_800_651, w_800_652, w_800_653, w_800_654, w_800_655, w_800_656, w_800_657, w_800_658, w_800_659, w_800_660, w_800_661, w_800_662, w_800_663, w_800_664, w_800_665, w_800_666, w_800_667, w_800_668, w_800_669, w_800_670, w_800_671, w_800_672, w_800_673, w_800_674, w_800_675, w_800_676, w_800_677, w_800_678, w_800_679, w_800_680, w_800_681, w_800_682, w_800_683, w_800_684, w_800_685, w_800_686, w_800_687, w_800_688, w_800_689, w_800_690, w_800_691, w_800_692, w_800_693, w_800_694, w_800_695, w_800_696, w_800_697, w_800_698, w_800_699, w_800_700, w_800_701, w_800_702, w_800_703, w_800_704, w_800_705, w_800_706, w_800_707, w_800_708, w_800_709, w_800_710, w_800_711, w_800_712, w_800_713, w_800_714, w_800_715, w_800_716, w_800_717;
  not1 I001_000(w_001_000, w_000_000);
  nand2 I001_001(w_001_001, w_000_001, w_000_002);
  not1 I001_002(w_001_002, w_000_003);
  or2  I001_003(w_001_003, w_000_004, w_000_005);
  nand2 I001_004(w_001_004, w_000_006, w_000_007);
  nand2 I001_005(w_001_005, w_000_008, w_000_009);
  not1 I001_006(w_001_006, w_000_010);
  and2 I001_007(w_001_007, w_000_011, w_000_012);
  nand2 I001_008(w_001_008, w_000_013, w_000_014);
  not1 I001_009(w_001_009, w_000_015);
  nand2 I001_010(w_001_010, w_000_016, w_000_017);
  or2  I001_011(w_001_011, w_000_018, w_000_019);
  not1 I001_012(w_001_012, w_000_020);
  nand2 I001_013(w_001_013, w_000_021, w_000_022);
  nand2 I001_014(w_001_014, w_000_023, w_000_024);
  or2  I001_015(w_001_015, w_000_025, w_000_026);
  and2 I001_016(w_001_016, w_000_027, w_000_028);
  and2 I001_017(w_001_017, w_000_029, w_000_030);
  or2  I001_018(w_001_018, w_000_031, w_000_032);
  and2 I001_019(w_001_019, w_000_033, w_000_034);
  not1 I001_020(w_001_020, w_000_035);
  and2 I001_021(w_001_021, w_000_036, w_000_037);
  or2  I001_022(w_001_022, w_000_038, w_000_039);
  and2 I001_023(w_001_023, w_000_040, w_000_041);
  or2  I001_024(w_001_024, w_000_042, w_000_043);
  and2 I001_025(w_001_025, w_000_044, w_000_045);
  or2  I001_026(w_001_026, w_000_046, w_000_047);
  not1 I001_027(w_001_027, w_000_048);
  nand2 I001_028(w_001_028, w_000_049, w_000_050);
  and2 I001_029(w_001_029, w_000_051, w_000_052);
  and2 I001_030(w_001_030, w_000_053, w_000_054);
  nand2 I001_031(w_001_031, w_000_055, w_000_056);
  and2 I001_032(w_001_032, w_000_057, w_000_058);
  and2 I001_033(w_001_033, w_000_059, w_000_060);
  not1 I001_034(w_001_034, w_000_061);
  not1 I001_035(w_001_035, w_000_062);
  nand2 I001_036(w_001_036, w_000_063, w_000_064);
  nand2 I002_000(w_002_000, w_001_016, w_000_065);
  and2 I002_001(w_002_001, w_000_066, w_001_021);
  not1 I002_002(w_002_002, w_001_006);
  or2  I002_003(w_002_003, w_000_067, w_000_068);
  nand2 I002_004(w_002_004, w_001_016, w_001_007);
  nand2 I002_005(w_002_005, w_001_009, w_001_034);
  or2  I002_006(w_002_006, w_001_001, w_001_032);
  nand2 I002_007(w_002_007, w_001_032, w_000_069);
  and2 I002_008(w_002_008, w_001_000, w_001_004);
  and2 I002_009(w_002_009, w_000_070, w_000_071);
  and2 I002_010(w_002_010, w_001_033, w_001_002);
  nand2 I002_011(w_002_011, w_001_022, w_000_072);
  or2  I002_012(w_002_012, w_000_073, w_000_074);
  and2 I002_013(w_002_013, w_000_075, w_001_027);
  nand2 I002_014(w_002_014, w_001_035, w_001_000);
  and2 I002_015(w_002_015, w_000_076, w_001_028);
  nand2 I002_016(w_002_016, w_001_008, w_001_021);
  nand2 I002_017(w_002_017, w_001_030, w_001_008);
  not1 I002_018(w_002_018, w_000_077);
  nand2 I002_019(w_002_019, w_000_078, w_000_004);
  nand2 I002_020(w_002_020, w_001_028, w_000_079);
  and2 I002_021(w_002_021, w_000_018, w_000_080);
  or2  I002_022(w_002_022, w_001_021, w_000_081);
  nand2 I002_023(w_002_023, w_000_082, w_000_083);
  and2 I002_024(w_002_024, w_001_007, w_000_084);
  nand2 I002_025(w_002_025, w_000_085, w_001_001);
  not1 I002_026(w_002_026, w_000_086);
  nand2 I002_027(w_002_027, w_001_004, w_000_087);
  not1 I002_028(w_002_028, w_000_088);
  nand2 I002_029(w_002_029, w_000_089, w_000_090);
  nand2 I002_030(w_002_030, w_000_091, w_001_024);
  not1 I002_031(w_002_031, w_000_092);
  and2 I002_032(w_002_032, w_000_093, w_000_094);
  or2  I002_033(w_002_033, w_000_095, w_000_096);
  and2 I002_034(w_002_034, w_001_018, w_000_097);
  and2 I002_035(w_002_035, w_000_098, w_001_010);
  and2 I002_036(w_002_036, w_001_025, w_001_015);
  not1 I002_037(w_002_037, w_001_035);
  and2 I002_038(w_002_038, w_001_029, w_001_025);
  and2 I002_039(w_002_039, w_001_025, w_001_024);
  not1 I002_040(w_002_040, w_001_015);
  not1 I002_041(w_002_041, w_000_099);
  not1 I002_042(w_002_042, w_000_100);
  not1 I002_043(w_002_043, w_000_101);
  or2  I002_044(w_002_044, w_000_102, w_000_103);
  and2 I002_045(w_002_045, w_000_104, w_001_002);
  and2 I002_046(w_002_046, w_000_105, w_001_014);
  or2  I002_047(w_002_047, w_001_024, w_001_011);
  nand2 I002_048(w_002_048, w_001_010, w_000_106);
  nand2 I002_049(w_002_049, w_000_107, w_001_036);
  nand2 I002_050(w_002_050, w_000_108, w_000_109);
  and2 I002_051(w_002_051, w_000_069, w_000_110);
  not1 I002_052(w_002_052, w_000_092);
  and2 I002_053(w_002_053, w_000_111, w_001_030);
  not1 I002_054(w_002_054, w_001_018);
  not1 I002_055(w_002_055, w_000_112);
  not1 I002_056(w_002_056, w_000_113);
  not1 I002_057(w_002_057, w_001_026);
  nand2 I002_058(w_002_058, w_000_114, w_001_017);
  and2 I002_059(w_002_059, w_001_036, w_001_028);
  not1 I002_060(w_002_060, w_001_001);
  not1 I002_061(w_002_061, w_001_025);
  or2  I002_062(w_002_062, w_001_014, w_001_030);
  or2  I002_063(w_002_063, w_001_021, w_000_115);
  and2 I002_064(w_002_064, w_000_116, w_000_117);
  or2  I002_065(w_002_065, w_000_118, w_000_119);
  and2 I002_066(w_002_066, w_000_120, w_000_036);
  and2 I002_067(w_002_067, w_001_019, w_001_015);
  or2  I002_068(w_002_068, w_000_090, w_000_121);
  not1 I002_069(w_002_069, w_000_122);
  and2 I002_070(w_002_070, w_000_123, w_001_020);
  not1 I002_071(w_002_071, w_001_004);
  nand2 I002_072(w_002_072, w_001_024, w_000_124);
  or2  I002_073(w_002_073, w_000_125, w_001_018);
  or2  I002_074(w_002_074, w_001_014, w_000_126);
  or2  I002_075(w_002_075, w_000_127, w_000_027);
  not1 I002_076(w_002_076, w_000_128);
  not1 I002_077(w_002_077, w_000_097);
  nand2 I002_078(w_002_078, w_001_017, w_000_028);
  nand2 I002_079(w_002_079, w_000_129, w_001_020);
  nand2 I002_080(w_002_080, w_001_024, w_000_130);
  and2 I002_081(w_002_081, w_001_016, w_000_131);
  or2  I002_082(w_002_082, w_000_132, w_001_032);
  nand2 I002_083(w_002_083, w_001_019, w_000_133);
  or2  I002_084(w_002_084, w_001_019, w_000_134);
  nand2 I002_085(w_002_085, w_001_011, w_001_013);
  not1 I002_086(w_002_086, w_000_135);
  or2  I002_087(w_002_087, w_000_136, w_001_005);
  and2 I002_088(w_002_088, w_001_023, w_001_007);
  or2  I002_090(w_002_090, w_000_139, w_000_140);
  or2  I002_091(w_002_091, w_000_141, w_001_018);
  and2 I002_092(w_002_092, w_000_142, w_000_143);
  not1 I002_093(w_002_093, w_000_144);
  not1 I002_094(w_002_094, w_001_035);
  nand2 I002_096(w_002_096, w_000_145, w_001_013);
  nand2 I002_097(w_002_097, w_000_146, w_000_147);
  and2 I002_098(w_002_098, w_000_012, w_001_010);
  or2  I002_099(w_002_099, w_001_015, w_001_034);
  and2 I002_100(w_002_100, w_001_032, w_000_148);
  not1 I002_101(w_002_101, w_000_084);
  and2 I002_102(w_002_102, w_001_014, w_000_149);
  or2  I002_103(w_002_103, w_001_000, w_001_013);
  or2  I002_104(w_002_104, w_000_150, w_001_030);
  nand2 I002_105(w_002_105, w_001_004, w_001_033);
  nand2 I002_106(w_002_106, w_001_034, w_001_011);
  not1 I002_107(w_002_107, w_001_003);
  not1 I002_108(w_002_108, w_001_002);
  or2  I002_109(w_002_109, w_001_025, w_000_151);
  or2  I002_110(w_002_110, w_001_036, w_001_030);
  nand2 I002_112(w_002_112, w_000_152, w_000_153);
  nand2 I002_113(w_002_113, w_001_012, w_001_009);
  not1 I002_114(w_002_114, w_001_014);
  nand2 I002_115(w_002_115, w_001_029, w_000_154);
  not1 I002_116(w_002_116, w_001_022);
  and2 I002_118(w_002_118, w_000_156, w_000_018);
  or2  I002_119(w_002_119, w_000_157, w_000_158);
  or2  I002_120(w_002_120, w_001_003, w_000_159);
  nand2 I002_121(w_002_121, w_001_004, w_001_033);
  and2 I002_123(w_002_123, w_000_161, w_001_012);
  and2 I002_124(w_002_124, w_001_020, w_000_091);
  nand2 I002_125(w_002_125, w_001_014, w_001_013);
  not1 I002_127(w_002_127, w_001_030);
  or2  I002_128(w_002_128, w_000_162, w_001_020);
  or2  I002_129(w_002_129, w_001_008, w_000_163);
  nand2 I002_130(w_002_130, w_001_029, w_001_022);
  nand2 I002_133(w_002_133, w_001_003, w_001_025);
  or2  I002_134(w_002_134, w_001_014, w_000_166);
  and2 I002_135(w_002_135, w_001_026, w_000_167);
  or2  I002_137(w_002_137, w_001_011, w_001_014);
  nand2 I002_139(w_002_139, w_001_014, w_001_017);
  or2  I002_141(w_002_141, w_000_171, w_001_027);
  and2 I002_142(w_002_142, w_001_015, w_000_011);
  nand2 I002_144(w_002_144, w_001_004, w_000_172);
  nand2 I002_145(w_002_145, w_000_040, w_001_028);
  not1 I002_146(w_002_146, w_000_173);
  nand2 I002_147(w_002_147, w_000_174, w_001_003);
  nand2 I002_148(w_002_148, w_000_175, w_000_176);
  nand2 I002_149(w_002_149, w_000_177, w_000_043);
  not1 I002_150(w_002_150, w_000_178);
  not1 I002_151(w_002_151, w_001_033);
  not1 I002_152(w_002_152, w_001_019);
  not1 I002_154(w_002_154, w_001_029);
  or2  I002_155(w_002_155, w_001_014, w_001_021);
  or2  I002_157(w_002_157, w_001_026, w_000_181);
  or2  I002_158(w_002_158, w_000_182, w_000_134);
  not1 I002_159(w_002_159, w_001_006);
  nand2 I002_161(w_002_161, w_001_026, w_000_183);
  and2 I002_162(w_002_162, w_000_184, w_001_030);
  not1 I002_163(w_002_163, w_001_031);
  nand2 I002_165(w_002_165, w_001_023, w_001_009);
  and2 I002_166(w_002_166, w_000_081, w_001_013);
  nand2 I002_167(w_002_167, w_000_185, w_000_186);
  or2  I002_168(w_002_168, w_001_028, w_001_000);
  nand2 I002_170(w_002_170, w_001_022, w_001_012);
  not1 I002_171(w_002_171, w_000_151);
  or2  I002_172(w_002_172, w_000_189, w_001_032);
  nand2 I002_173(w_002_173, w_001_027, w_001_022);
  not1 I002_174(w_002_174, w_001_024);
  and2 I002_175(w_002_175, w_000_177, w_001_002);
  and2 I002_176(w_002_176, w_000_190, w_000_191);
  or2  I002_178(w_002_178, w_000_193, w_001_033);
  and2 I002_179(w_002_179, w_000_194, w_000_195);
  and2 I002_180(w_002_180, w_001_022, w_000_196);
  and2 I002_181(w_002_181, w_000_197, w_001_017);
  not1 I002_182(w_002_182, w_001_014);
  nand2 I002_183(w_002_183, w_000_198, w_001_022);
  or2  I002_184(w_002_184, w_001_008, w_000_199);
  nand2 I002_186(w_002_186, w_000_200, w_001_029);
  and2 I002_188(w_002_188, w_000_202, w_001_031);
  and2 I002_189(w_002_189, w_001_004, w_001_006);
  or2  I002_190(w_002_190, w_001_028, w_000_152);
  or2  I002_191(w_002_191, w_001_032, w_000_098);
  and2 I002_192(w_002_192, w_001_036, w_001_029);
  and2 I002_193(w_002_193, w_000_203, w_000_204);
  not1 I002_194(w_002_194, w_001_000);
  and2 I002_195(w_002_195, w_000_045, w_000_205);
  or2  I002_196(w_002_196, w_001_005, w_001_034);
  or2  I002_198(w_002_198, w_001_030, w_001_036);
  and2 I002_200(w_002_200, w_000_206, w_000_207);
  or2  I002_201(w_002_201, w_000_208, w_001_032);
  nand2 I002_202(w_002_202, w_000_209, w_001_017);
  nand2 I002_204(w_002_204, w_000_187, w_000_190);
  or2  I002_205(w_002_205, w_000_210, w_001_015);
  or2  I002_206(w_002_206, w_001_013, w_001_033);
  and2 I002_207(w_002_207, w_000_106, w_000_211);
  nand2 I002_209(w_002_209, w_001_023, w_000_212);
  or2  I002_210(w_002_210, w_000_170, w_000_213);
  and2 I002_211(w_002_211, w_001_007, w_001_011);
  not1 I002_212(w_002_212, w_000_183);
  nand2 I002_213(w_002_213, w_001_032, w_000_214);
  or2  I002_214(w_002_214, w_000_215, w_001_024);
  or2  I002_215(w_002_215, w_000_216, w_000_217);
  or2  I002_216(w_002_216, w_001_026, w_000_218);
  nand2 I002_217(w_002_217, w_001_008, w_000_156);
  and2 I002_218(w_002_218, w_001_016, w_000_219);
  not1 I002_219(w_002_219, w_001_029);
  or2  I002_220(w_002_220, w_001_021, w_000_220);
  not1 I002_221(w_002_221, w_000_221);
  nand2 I002_222(w_002_222, w_000_222, w_000_223);
  nand2 I002_223(w_002_223, w_001_022, w_001_001);
  nand2 I002_224(w_002_224, w_000_224, w_001_030);
  nand2 I002_225(w_002_225, w_000_225, w_001_031);
  not1 I002_226(w_002_226, w_001_019);
  and2 I002_227(w_002_227, w_000_129, w_000_068);
  nand2 I002_228(w_002_228, w_000_226, w_001_007);
  and2 I002_229(w_002_229, w_001_007, w_001_006);
  or2  I002_230(w_002_230, w_001_003, w_001_000);
  or2  I002_231(w_002_231, w_000_227, w_001_005);
  or2  I002_233(w_002_233, w_001_015, w_001_023);
  or2  I002_234(w_002_234, w_001_017, w_000_162);
  not1 I002_236(w_002_236, w_001_012);
  and2 I002_237(w_002_237, w_000_229, w_000_230);
  or2  I002_238(w_002_238, w_001_007, w_000_231);
  not1 I002_239(w_002_239, w_001_036);
  not1 I002_240(w_002_240, w_000_221);
  not1 I002_243(w_002_243, w_001_003);
  or2  I002_244(w_002_244, w_000_234, w_000_033);
  nand2 I002_246(w_002_246, w_001_028, w_000_235);
  not1 I002_247(w_002_247, w_000_236);
  not1 I002_249(w_002_249, w_001_010);
  not1 I002_250(w_002_250, w_001_003);
  nand2 I002_251(w_002_251, w_001_009, w_000_237);
  and2 I002_252(w_002_252, w_001_000, w_001_026);
  or2  I002_253(w_002_253, w_000_238, w_001_012);
  nand2 I002_256(w_002_256, w_000_037, w_000_239);
  not1 I002_257(w_002_257, w_001_020);
  and2 I002_258(w_002_258, w_001_009, w_001_018);
  and2 I002_259(w_002_259, w_000_021, w_000_240);
  nand2 I002_260(w_002_260, w_001_006, w_000_241);
  nand2 I002_261(w_002_261, w_000_045, w_000_242);
  nand2 I002_262(w_002_262, w_001_004, w_000_243);
  not1 I002_263(w_002_263, w_000_244);
  and2 I002_264(w_002_264, w_000_245, w_000_246);
  and2 I002_265(w_002_265, w_001_020, w_000_247);
  not1 I002_266(w_002_266, w_000_248);
  or2  I002_267(w_002_267, w_001_025, w_001_009);
  nand2 I002_268(w_002_268, w_001_013, w_001_016);
  and2 I002_269(w_002_269, w_001_034, w_001_000);
  nand2 I002_270(w_002_270, w_001_014, w_001_001);
  and2 I002_271(w_002_271, w_000_171, w_000_249);
  nand2 I002_272(w_002_272, w_000_250, w_001_016);
  not1 I002_273(w_002_273, w_000_251);
  not1 I002_274(w_002_274, w_000_252);
  or2  I002_275(w_002_275, w_001_016, w_001_022);
  not1 I002_276(w_002_276, w_000_253);
  or2  I002_277(w_002_277, w_000_239, w_001_004);
  not1 I002_278(w_002_278, w_000_254);
  not1 I002_279(w_002_279, w_001_024);
  and2 I002_280(w_002_280, w_001_012, w_001_013);
  or2  I002_282(w_002_282, w_000_026, w_000_255);
  or2  I002_283(w_002_283, w_000_256, w_001_006);
  nand2 I002_285(w_002_285, w_001_017, w_001_009);
  and2 I002_286(w_002_286, w_001_034, w_000_257);
  not1 I002_287(w_002_287, w_001_013);
  or2  I002_288(w_002_288, w_001_001, w_000_250);
  and2 I002_289(w_002_289, w_000_258, w_001_013);
  or2  I002_290(w_002_290, w_001_021, w_000_107);
  or2  I002_291(w_002_291, w_001_015, w_000_259);
  and2 I002_292(w_002_292, w_001_009, w_000_260);
  or2  I002_293(w_002_293, w_000_261, w_001_023);
  nand2 I002_295(w_002_295, w_001_016, w_001_019);
  nand2 I002_296(w_002_296, w_000_264, w_000_265);
  or2  I002_297(w_002_297, w_001_021, w_001_007);
  and2 I002_298(w_002_298, w_001_028, w_001_035);
  or2  I002_299(w_002_299, w_000_266, w_000_267);
  nand2 I002_300(w_002_300, w_001_027, w_000_187);
  nand2 I002_301(w_002_301, w_001_031, w_000_194);
  and2 I002_302(w_002_302, w_000_268, w_000_218);
  and2 I002_303(w_002_303, w_001_017, w_001_025);
  or2  I002_304(w_002_304, w_001_031, w_000_098);
  or2  I002_305(w_002_305, w_000_178, w_001_011);
  or2  I002_306(w_002_306, w_000_269, w_000_270);
  not1 I002_307(w_002_307, w_000_271);
  or2  I002_308(w_002_308, w_000_272, w_001_014);
  nand2 I002_309(w_002_309, w_001_011, w_001_017);
  or2  I002_310(w_002_310, w_000_261, w_000_273);
  nand2 I002_311(w_002_311, w_001_007, w_000_274);
  nand2 I002_312(w_002_312, w_001_034, w_000_275);
  not1 I002_313(w_002_313, w_001_023);
  or2  I002_315(w_002_315, w_001_005, w_000_276);
  or2  I002_316(w_002_316, w_001_032, w_000_277);
  not1 I002_317(w_002_317, w_000_216);
  or2  I002_318(w_002_318, w_001_034, w_001_033);
  nand2 I002_319(w_002_319, w_001_026, w_000_278);
  nand2 I002_320(w_002_320, w_001_004, w_000_262);
  not1 I002_321(w_002_321, w_001_030);
  and2 I002_322(w_002_322, w_000_197, w_000_279);
  not1 I002_323(w_002_323, w_000_280);
  and2 I002_324(w_002_324, w_000_118, w_001_002);
  not1 I002_326(w_002_326, w_001_027);
  not1 I002_327(w_002_327, w_000_283);
  nand2 I002_328(w_002_328, w_000_284, w_001_019);
  nand2 I002_329(w_002_329, w_000_285, w_000_182);
  or2  I002_330(w_002_330, w_001_035, w_001_025);
  or2  I002_331(w_002_331, w_001_032, w_000_286);
  not1 I002_334(w_002_334, w_000_270);
  and2 I002_335(w_002_335, w_001_007, w_001_026);
  not1 I002_337(w_002_337, w_001_026);
  nand2 I002_338(w_002_338, w_000_289, w_001_006);
  nand2 I002_340(w_002_340, w_001_005, w_001_003);
  or2  I002_341(w_002_341, w_001_021, w_000_290);
  or2  I002_342(w_002_342, w_001_018, w_001_024);
  not1 I002_343(w_002_343, w_000_291);
  not1 I002_344(w_002_344, w_001_006);
  nand2 I002_345(w_002_345, w_000_292, w_001_010);
  or2  I002_346(w_002_346, w_000_293, w_001_000);
  and2 I002_347(w_002_347, w_000_294, w_001_026);
  or2  I002_349(w_002_349, w_000_296, w_000_297);
  or2  I002_350(w_002_350, w_000_298, w_000_299);
  or2  I002_351(w_002_351, w_001_016, w_000_300);
  or2  I002_352(w_002_352, w_001_002, w_000_301);
  and2 I002_353(w_002_353, w_001_026, w_001_033);
  or2  I002_354(w_002_354, w_000_302, w_000_252);
  nand2 I002_357(w_002_357, w_000_303, w_001_030);
  nand2 I002_358(w_002_358, w_000_304, w_001_021);
  and2 I002_359(w_002_359, w_001_024, w_001_001);
  not1 I002_360(w_002_360, w_000_305);
  nand2 I002_361(w_002_361, w_001_008, w_000_262);
  and2 I002_362(w_002_362, w_001_021, w_000_306);
  and2 I002_363(w_002_363, w_001_018, w_001_006);
  or2  I002_365(w_002_365, w_001_033, w_000_307);
  not1 I002_366(w_002_366, w_000_012);
  or2  I002_367(w_002_367, w_001_029, w_000_308);
  not1 I002_368(w_002_368, w_001_000);
  not1 I002_369(w_002_369, w_001_009);
  not1 I002_370(w_002_370, w_001_021);
  and2 I002_372(w_002_372, w_001_024, w_000_309);
  nand2 I002_373(w_002_373, w_001_011, w_000_310);
  and2 I002_374(w_002_374, w_000_311, w_000_104);
  nand2 I002_375(w_002_375, w_001_010, w_001_013);
  or2  I002_376(w_002_376, w_000_236, w_000_312);
  not1 I002_377(w_002_377, w_000_173);
  or2  I002_378(w_002_378, w_001_030, w_001_028);
  or2  I002_379(w_002_379, w_001_008, w_000_313);
  and2 I002_380(w_002_380, w_001_036, w_000_314);
  not1 I002_383(w_002_383, w_001_010);
  or2  I002_384(w_002_384, w_001_034, w_001_016);
  not1 I002_385(w_002_385, w_000_318);
  nand2 I002_386(w_002_386, w_001_000, w_000_319);
  nand2 I002_389(w_002_389, w_000_321, w_001_022);
  and2 I002_390(w_002_390, w_000_322, w_001_033);
  nand2 I002_391(w_002_391, w_000_323, w_001_019);
  and2 I002_392(w_002_392, w_000_324, w_000_325);
  nand2 I002_393(w_002_393, w_001_013, w_000_326);
  not1 I002_396(w_002_396, w_000_034);
  or2  I002_397(w_002_397, w_000_328, w_000_108);
  and2 I002_398(w_002_398, w_000_329, w_000_330);
  and2 I002_400(w_002_400, w_000_331, w_000_330);
  and2 I002_401(w_002_401, w_001_029, w_000_156);
  or2  I002_402(w_002_402, w_000_332, w_000_333);
  not1 I002_403(w_002_403, w_001_014);
  not1 I002_405(w_002_405, w_001_007);
  not1 I002_406(w_002_406, w_000_123);
  or2  I002_407(w_002_407, w_000_215, w_001_025);
  or2  I002_408(w_002_408, w_001_021, w_000_335);
  and2 I002_409(w_002_409, w_000_292, w_000_336);
  or2  I002_411(w_002_411, w_000_260, w_000_337);
  nand2 I002_412(w_002_412, w_001_020, w_001_011);
  nand2 I002_413(w_002_413, w_000_338, w_000_339);
  or2  I002_414(w_002_414, w_001_015, w_000_065);
  or2  I002_415(w_002_415, w_000_176, w_001_013);
  not1 I002_416(w_002_416, w_001_025);
  nand2 I002_417(w_002_417, w_000_199, w_001_005);
  and2 I002_418(w_002_418, w_001_000, w_001_001);
  not1 I002_419(w_002_419, w_000_340);
  or2  I002_420(w_002_420, w_000_341, w_001_034);
  or2  I002_421(w_002_421, w_000_119, w_001_020);
  not1 I002_423(w_002_423, w_000_342);
  not1 I002_424(w_002_424, w_000_030);
  nand2 I002_425(w_002_425, w_001_005, w_000_047);
  or2  I002_426(w_002_426, w_000_343, w_001_018);
  nand2 I002_427(w_002_427, w_001_013, w_001_032);
  and2 I002_428(w_002_428, w_001_004, w_000_061);
  and2 I002_429(w_002_429, w_000_344, w_000_269);
  nand2 I002_433(w_002_433, w_000_348, w_001_003);
  or2  I002_434(w_002_434, w_000_349, w_001_014);
  and2 I002_435(w_002_435, w_001_021, w_000_350);
  not1 I002_436(w_002_436, w_000_184);
  and2 I002_438(w_002_438, w_000_351, w_001_031);
  and2 I002_439(w_002_439, w_000_139, w_000_035);
  nand2 I002_440(w_002_440, w_000_352, w_000_353);
  not1 I002_441(w_002_441, w_000_278);
  and2 I002_442(w_002_442, w_001_018, w_001_033);
  not1 I002_443(w_002_443, w_001_008);
  or2  I002_444(w_002_444, w_001_035, w_000_354);
  not1 I002_445(w_002_445, w_000_165);
  nand2 I002_446(w_002_446, w_000_355, w_000_249);
  nand2 I002_447(w_002_447, w_001_006, w_000_001);
  not1 I002_448(w_002_448, w_000_356);
  not1 I002_449(w_002_449, w_000_357);
  not1 I002_450(w_002_450, w_000_358);
  not1 I002_451(w_002_451, w_000_359);
  or2  I002_452(w_002_452, w_001_030, w_001_029);
  or2  I002_453(w_002_453, w_001_034, w_000_360);
  and2 I002_455(w_002_455, w_001_005, w_001_025);
  not1 I002_457(w_002_457, w_001_019);
  or2  I002_458(w_002_458, w_001_018, w_000_362);
  not1 I002_459(w_002_459, w_001_025);
  and2 I002_460(w_002_460, w_000_363, w_000_364);
  or2  I002_461(w_002_461, w_000_365, w_000_366);
  nand2 I002_462(w_002_462, w_000_367, w_000_368);
  or2  I002_464(w_002_464, w_001_009, w_000_370);
  or2  I002_465(w_002_465, w_000_371, w_001_034);
  and2 I002_466(w_002_466, w_001_031, w_000_282);
  nand2 I002_467(w_002_467, w_001_011, w_001_009);
  or2  I002_468(w_002_468, w_000_166, w_001_019);
  and2 I002_469(w_002_469, w_000_008, w_000_372);
  or2  I002_470(w_002_470, w_001_027, w_001_009);
  nand2 I002_471(w_002_471, w_000_373, w_001_032);
  and2 I002_472(w_002_472, w_001_025, w_000_075);
  or2  I002_473(w_002_473, w_000_200, w_001_007);
  not1 I002_474(w_002_474, w_000_349);
  and2 I002_475(w_002_475, w_001_031, w_000_243);
  and2 I002_477(w_002_477, w_000_096, w_001_033);
  not1 I002_478(w_002_478, w_000_228);
  not1 I002_479(w_002_479, w_001_031);
  not1 I002_480(w_002_480, w_000_374);
  not1 I002_481(w_002_481, w_001_019);
  or2  I002_482(w_002_482, w_001_034, w_001_014);
  or2  I002_485(w_002_485, w_000_377, w_000_378);
  not1 I002_486(w_002_486, w_001_010);
  and2 I002_487(w_002_487, w_000_021, w_001_015);
  not1 I002_488(w_002_488, w_000_078);
  or2  I002_489(w_002_489, w_001_018, w_001_009);
  nand2 I002_490(w_002_490, w_000_175, w_000_379);
  and2 I002_491(w_002_491, w_000_380, w_000_302);
  not1 I002_493(w_002_493, w_001_012);
  nand2 I002_494(w_002_494, w_001_035, w_001_025);
  and2 I002_495(w_002_495, w_000_381, w_000_382);
  not1 I002_496(w_002_496, w_000_181);
  and2 I002_497(w_002_497, w_001_033, w_000_062);
  nand2 I002_498(w_002_498, w_001_015, w_001_031);
  or2  I002_499(w_002_499, w_000_383, w_000_372);
  nand2 I002_500(w_002_500, w_001_011, w_001_020);
  not1 I002_501(w_002_501, w_000_384);
  not1 I002_502(w_002_502, w_001_030);
  not1 I002_503(w_002_503, w_000_228);
  not1 I002_504(w_002_504, w_001_029);
  or2  I002_505(w_002_505, w_000_065, w_001_011);
  not1 I002_507(w_002_507, w_001_004);
  or2  I002_509(w_002_509, w_000_300, w_000_320);
  or2  I002_510(w_002_510, w_000_150, w_001_019);
  or2  I002_511(w_002_511, w_000_386, w_000_324);
  not1 I002_512(w_002_512, w_000_109);
  not1 I002_513(w_002_513, w_000_354);
  or2  I002_514(w_002_514, w_001_016, w_000_260);
  nand2 I002_515(w_002_515, w_001_003, w_001_007);
  nand2 I002_516(w_002_516, w_001_030, w_001_000);
  nand2 I002_517(w_002_517, w_001_017, w_000_186);
  or2  I002_518(w_002_518, w_001_009, w_001_024);
  or2  I002_519(w_002_519, w_001_023, w_001_009);
  nand2 I002_520(w_002_520, w_000_387, w_001_022);
  and2 I002_522(w_002_522, w_000_232, w_001_022);
  or2  I002_523(w_002_523, w_000_225, w_001_031);
  nand2 I002_524(w_002_524, w_000_286, w_000_388);
  or2  I002_526(w_002_526, w_001_034, w_001_025);
  and2 I002_528(w_002_528, w_001_014, w_000_035);
  not1 I002_529(w_002_529, w_001_020);
  and2 I002_530(w_002_530, w_000_391, w_001_003);
  and2 I002_531(w_002_531, w_000_063, w_001_017);
  and2 I002_532(w_002_532, w_000_392, w_001_034);
  not1 I002_533(w_002_533, w_000_393);
  and2 I002_534(w_002_534, w_001_000, w_000_394);
  not1 I002_535(w_002_535, w_001_004);
  not1 I002_536(w_002_536, w_000_038);
  not1 I002_537(w_002_537, w_000_395);
  and2 I002_538(w_002_538, w_001_007, w_001_002);
  or2  I002_540(w_002_540, w_001_010, w_000_396);
  and2 I002_541(w_002_541, w_000_302, w_001_032);
  and2 I002_542(w_002_542, w_001_020, w_001_003);
  and2 I002_543(w_002_543, w_001_023, w_000_339);
  not1 I002_545(w_002_545, w_000_119);
  nand2 I002_547(w_002_547, w_001_030, w_001_022);
  or2  I002_548(w_002_548, w_001_013, w_001_036);
  nand2 I002_549(w_002_549, w_000_331, w_000_399);
  and2 I002_550(w_002_550, w_000_400, w_000_401);
  and2 I002_551(w_002_551, w_000_402, w_000_403);
  and2 I002_552(w_002_552, w_000_404, w_000_405);
  and2 I002_553(w_002_553, w_001_030, w_001_012);
  or2  I002_554(w_002_554, w_001_026, w_000_170);
  or2  I002_557(w_002_557, w_000_368, w_000_108);
  or2  I002_558(w_002_558, w_000_408, w_001_026);
  and2 I002_560(w_002_560, w_001_005, w_000_326);
  not1 I002_561(w_002_561, w_000_376);
  or2  I002_562(w_002_562, w_001_019, w_000_259);
  not1 I002_563(w_002_563, w_001_029);
  and2 I002_564(w_002_564, w_001_027, w_000_409);
  and2 I002_565(w_002_565, w_000_410, w_000_411);
  not1 I002_566(w_002_566, w_001_007);
  and2 I002_567(w_002_567, w_000_412, w_000_413);
  and2 I002_568(w_002_568, w_000_414, w_001_024);
  not1 I002_569(w_002_569, w_000_376);
  or2  I002_570(w_002_570, w_001_010, w_000_338);
  not1 I002_571(w_002_571, w_001_029);
  and2 I002_572(w_002_572, w_001_028, w_000_320);
  not1 I002_574(w_002_574, w_000_415);
  and2 I002_575(w_002_575, w_000_416, w_001_031);
  or2  I002_576(w_002_576, w_000_417, w_001_006);
  and2 I002_577(w_002_577, w_001_011, w_001_008);
  or2  I002_578(w_002_578, w_000_148, w_001_026);
  and2 I002_579(w_002_579, w_000_418, w_001_034);
  or2  I002_580(w_002_580, w_001_007, w_001_021);
  not1 I002_581(w_002_581, w_001_005);
  or2  I002_582(w_002_582, w_000_419, w_000_070);
  or2  I002_583(w_002_583, w_001_017, w_000_420);
  not1 I002_584(w_002_584, w_000_159);
  not1 I002_585(w_002_585, w_001_000);
  not1 I002_586(w_002_586, w_001_013);
  nand2 I002_587(w_002_587, w_000_030, w_001_021);
  or2  I002_588(w_002_588, w_000_096, w_001_011);
  not1 I002_589(w_002_589, w_001_003);
  and2 I002_590(w_002_590, w_000_403, w_000_421);
  or2  I002_591(w_002_591, w_000_339, w_000_152);
  or2  I002_592(w_002_592, w_001_026, w_000_304);
  or2  I002_593(w_002_593, w_000_313, w_000_422);
  and2 I002_594(w_002_594, w_001_019, w_001_027);
  or2  I002_595(w_002_595, w_000_348, w_001_006);
  not1 I002_596(w_002_596, w_001_026);
  or2  I002_597(w_002_597, w_001_008, w_000_423);
  not1 I002_598(w_002_598, w_000_032);
  and2 I002_599(w_002_599, w_001_018, w_000_061);
  and2 I002_600(w_002_600, w_000_424, w_000_425);
  nand2 I002_601(w_002_601, w_000_157, w_000_248);
  not1 I002_602(w_002_602, w_001_000);
  or2  I002_603(w_002_603, w_001_014, w_001_002);
  nand2 I002_604(w_002_604, w_000_426, w_000_427);
  not1 I002_605(w_002_605, w_000_139);
  not1 I002_606(w_002_606, w_000_342);
  or2  I002_607(w_002_607, w_001_028, w_001_023);
  not1 I002_608(w_002_608, w_000_428);
  not1 I002_609(w_002_609, w_000_160);
  not1 I002_610(w_002_610, w_000_023);
  and2 I002_612(w_002_612, w_001_001, w_000_093);
  or2  I002_613(w_002_613, w_000_430, w_001_027);
  nand2 I002_614(w_002_614, w_000_431, w_001_011);
  not1 I002_615(w_002_615, w_001_031);
  not1 I002_616(w_002_616, w_001_019);
  not1 I002_617(w_002_617, w_000_432);
  not1 I002_618(w_002_618, w_000_433);
  or2  I002_619(w_002_619, w_001_022, w_001_025);
  not1 I002_620(w_002_620, w_000_434);
  and2 I002_621(w_002_621, w_001_021, w_000_435);
  and2 I002_622(w_002_622, w_001_028, w_000_232);
  nand2 I002_623(w_002_623, w_000_436, w_000_037);
  and2 I002_624(w_002_624, w_001_001, w_000_437);
  or2  I002_625(w_002_625, w_001_018, w_000_438);
  nand2 I002_626(w_002_626, w_001_033, w_001_024);
  nand2 I002_627(w_002_627, w_001_000, w_000_057);
  not1 I002_628(w_002_628, w_000_439);
  nand2 I002_629(w_002_629, w_001_026, w_000_061);
  or2  I002_631(w_002_631, w_000_271, w_000_441);
  nand2 I002_632(w_002_632, w_000_287, w_000_279);
  or2  I002_633(w_002_633, w_001_007, w_000_442);
  and2 I002_634(w_002_634, w_000_443, w_001_022);
  nand2 I002_635(w_002_635, w_000_444, w_001_010);
  or2  I002_636(w_002_636, w_001_018, w_000_445);
  not1 I002_638(w_002_638, w_000_103);
  or2  I002_639(w_002_639, w_000_446, w_001_004);
  nand2 I002_640(w_002_640, w_000_136, w_001_001);
  or2  I002_642(w_002_642, w_000_448, w_000_170);
  and2 I002_643(w_002_643, w_001_022, w_000_282);
  not1 I002_644(w_002_644, w_000_449);
  and2 I002_645(w_002_645, w_000_353, w_001_010);
  nand2 I002_646(w_002_646, w_000_450, w_001_007);
  nand2 I002_647(w_002_647, w_000_338, w_000_144);
  and2 I002_648(w_002_648, w_000_283, w_001_000);
  nand2 I002_650(w_002_650, w_001_004, w_001_010);
  not1 I002_651(w_002_651, w_001_001);
  not1 I002_652(w_002_652, w_001_017);
  nand2 I002_653(w_002_653, w_000_050, w_001_026);
  or2  I002_654(w_002_654, w_001_035, w_001_030);
  nand2 I002_655(w_002_655, w_000_451, w_001_027);
  and2 I002_656(w_002_656, w_001_018, w_000_452);
  or2  I002_657(w_002_657, w_001_021, w_000_090);
  and2 I002_658(w_002_658, w_000_388, w_000_453);
  not1 I002_659(w_002_659, w_001_029);
  and2 I002_660(w_002_660, w_000_140, w_001_023);
  nand2 I002_661(w_002_661, w_001_031, w_001_007);
  and2 I002_662(w_002_662, w_000_454, w_001_005);
  nand2 I002_664(w_002_664, w_000_372, w_000_440);
  and2 I002_665(w_002_665, w_000_380, w_000_431);
  nand2 I002_666(w_002_666, w_001_013, w_001_027);
  nand2 I002_667(w_002_667, w_001_009, w_000_455);
  or2  I002_668(w_002_668, w_001_009, w_000_128);
  nand2 I002_669(w_002_669, w_001_004, w_000_456);
  not1 I002_671(w_002_671, w_001_000);
  not1 I002_672(w_002_672, w_001_007);
  and2 I002_673(w_002_673, w_001_030, w_001_015);
  nand2 I002_674(w_002_674, w_000_457, w_000_458);
  not1 I002_676(w_002_676, w_001_013);
  or2  I002_677(w_002_677, w_001_004, w_001_029);
  and2 I002_678(w_002_678, w_001_030, w_000_327);
  nand2 I002_679(w_002_679, w_001_001, w_001_027);
  nand2 I002_681(w_002_681, w_000_446, w_001_010);
  not1 I002_682(w_002_682, w_000_108);
  and2 I002_683(w_002_683, w_001_010, w_001_012);
  and2 I002_684(w_002_684, w_000_129, w_001_003);
  not1 I002_685(w_002_685, w_001_017);
  or2  I002_686(w_002_686, w_000_460, w_000_461);
  nand2 I002_688(w_002_688, w_000_072, w_000_175);
  or2  I002_690(w_002_690, w_001_029, w_000_181);
  not1 I002_691(w_002_691, w_001_019);
  and2 I002_692(w_002_692, w_000_420, w_001_030);
  nand2 I002_693(w_002_693, w_001_032, w_001_012);
  nand2 I002_694(w_002_694, w_001_008, w_000_462);
  or2  I002_695(w_002_695, w_000_463, w_000_298);
  nand2 I002_696(w_002_696, w_000_464, w_001_032);
  not1 I002_697(w_002_697, w_001_010);
  and2 I002_698(w_002_698, w_000_465, w_000_372);
  nand2 I002_699(w_002_699, w_001_009, w_001_035);
  or2  I002_701(w_002_701, w_000_250, w_001_007);
  nand2 I002_702(w_002_702, w_001_010, w_000_467);
  or2  I002_703(w_002_703, w_000_006, w_000_241);
  nand2 I002_705(w_002_705, w_000_251, w_000_469);
  or2  I002_706(w_002_706, w_001_000, w_001_012);
  and2 I002_707(w_002_707, w_000_386, w_000_470);
  and2 I002_708(w_002_708, w_001_007, w_001_016);
  nand2 I002_709(w_002_709, w_000_471, w_001_011);
  not1 I002_710(w_002_710, w_001_014);
  not1 I002_711(w_002_711, w_001_023);
  or2  I003_000(w_003_000, w_000_235, w_002_605);
  or2  I003_001(w_003_001, w_002_548, w_001_014);
  or2  I003_002(w_003_002, w_001_002, w_001_014);
  or2  I003_003(w_003_003, w_000_464, w_000_022);
  nand2 I003_004(w_003_004, w_002_560, w_000_126);
  or2  I003_005(w_003_005, w_001_018, w_000_472);
  or2  I003_006(w_003_006, w_001_004, w_001_021);
  not1 I003_007(w_003_007, w_001_015);
  not1 I003_008(w_003_008, w_002_058);
  nand2 I003_009(w_003_009, w_001_028, w_000_473);
  not1 I003_010(w_003_010, w_000_474);
  or2  I003_011(w_003_011, w_000_475, w_001_029);
  and2 I003_012(w_003_012, w_000_476, w_002_496);
  not1 I003_013(w_003_013, w_000_281);
  not1 I003_014(w_003_014, w_000_302);
  or2  I003_015(w_003_015, w_000_424, w_000_472);
  nand2 I003_016(w_003_016, w_002_647, w_001_003);
  nand2 I003_017(w_003_017, w_001_031, w_000_040);
  or2  I003_018(w_003_018, w_001_016, w_002_621);
  and2 I003_019(w_003_019, w_002_669, w_000_477);
  nand2 I003_020(w_003_020, w_001_016, w_001_019);
  or2  I003_021(w_003_021, w_000_172, w_002_229);
  and2 I003_022(w_003_022, w_001_014, w_000_478);
  or2  I003_023(w_003_023, w_000_026, w_001_027);
  not1 I003_024(w_003_024, w_001_023);
  and2 I003_025(w_003_025, w_001_025, w_000_224);
  and2 I003_026(w_003_026, w_001_020, w_002_040);
  nand2 I003_027(w_003_027, w_001_018, w_001_015);
  nand2 I003_028(w_003_028, w_000_204, w_002_550);
  nand2 I003_029(w_003_029, w_002_078, w_001_017);
  and2 I003_030(w_003_030, w_001_003, w_000_232);
  nand2 I003_031(w_003_031, w_001_021, w_000_479);
  not1 I003_032(w_003_032, w_001_018);
  not1 I003_033(w_003_033, w_001_017);
  not1 I003_034(w_003_034, w_002_369);
  not1 I003_035(w_003_035, w_002_112);
  and2 I003_036(w_003_036, w_000_447, w_000_255);
  or2  I003_037(w_003_037, w_001_030, w_002_052);
  or2  I003_038(w_003_038, w_000_415, w_001_025);
  not1 I003_039(w_003_039, w_000_420);
  not1 I003_040(w_003_040, w_000_470);
  and2 I003_041(w_003_041, w_001_026, w_000_239);
  or2  I003_042(w_003_042, w_000_480, w_002_504);
  or2  I003_043(w_003_043, w_000_151, w_002_108);
  and2 I003_044(w_003_044, w_000_023, w_000_172);
  or2  I003_045(w_003_045, w_000_139, w_002_346);
  not1 I003_046(w_003_046, w_000_319);
  and2 I003_047(w_003_047, w_002_077, w_000_481);
  or2  I003_048(w_003_048, w_000_482, w_002_447);
  not1 I003_049(w_003_049, w_001_022);
  and2 I003_050(w_003_050, w_002_207, w_000_096);
  nand2 I003_051(w_003_051, w_002_471, w_000_483);
  and2 I003_052(w_003_052, w_001_019, w_000_143);
  and2 I003_053(w_003_053, w_001_018, w_001_023);
  nand2 I003_054(w_003_054, w_000_396, w_001_000);
  or2  I003_055(w_003_055, w_000_296, w_001_007);
  nand2 I003_056(w_003_056, w_002_217, w_002_167);
  or2  I003_057(w_003_057, w_001_009, w_000_074);
  or2  I003_058(w_003_058, w_000_484, w_000_100);
  not1 I003_059(w_003_059, w_000_066);
  and2 I003_060(w_003_060, w_002_200, w_002_438);
  or2  I003_061(w_003_061, w_001_031, w_002_074);
  not1 I003_062(w_003_062, w_001_031);
  not1 I003_063(w_003_063, w_000_485);
  and2 I003_064(w_003_064, w_000_486, w_002_552);
  and2 I003_065(w_003_065, w_002_530, w_001_027);
  not1 I003_066(w_003_066, w_000_430);
  not1 I003_067(w_003_067, w_001_029);
  nand2 I003_068(w_003_068, w_001_001, w_001_036);
  or2  I003_069(w_003_069, w_002_020, w_001_020);
  not1 I003_070(w_003_070, w_000_024);
  or2  I003_071(w_003_071, w_002_269, w_000_487);
  nand2 I003_072(w_003_072, w_002_320, w_000_309);
  not1 I003_073(w_003_073, w_000_488);
  and2 I003_074(w_003_074, w_001_001, w_002_020);
  or2  I003_075(w_003_075, w_001_027, w_002_086);
  nand2 I003_076(w_003_076, w_002_370, w_001_013);
  and2 I003_077(w_003_077, w_002_034, w_000_021);
  nand2 I003_078(w_003_078, w_000_153, w_000_396);
  not1 I003_079(w_003_079, w_001_002);
  and2 I003_080(w_003_080, w_002_045, w_000_489);
  nand2 I003_081(w_003_081, w_000_458, w_002_612);
  and2 I003_082(w_003_082, w_002_162, w_001_020);
  and2 I003_083(w_003_083, w_000_490, w_001_004);
  not1 I003_084(w_003_084, w_002_016);
  nand2 I004_000(w_004_000, w_001_035, w_003_034);
  not1 I004_001(w_004_001, w_000_491);
  not1 I004_002(w_004_002, w_001_025);
  and2 I004_003(w_004_003, w_000_431, w_002_105);
  and2 I004_004(w_004_004, w_003_003, w_002_439);
  nand2 I004_005(w_004_005, w_003_084, w_003_020);
  or2  I004_006(w_004_006, w_001_000, w_001_001);
  or2  I004_007(w_004_007, w_003_013, w_000_086);
  and2 I004_008(w_004_008, w_001_006, w_002_538);
  or2  I004_009(w_004_009, w_002_523, w_001_034);
  and2 I004_010(w_004_010, w_001_020, w_000_492);
  not1 I004_011(w_004_011, w_003_060);
  or2  I004_012(w_004_012, w_002_590, w_002_547);
  or2  I004_013(w_004_013, w_000_137, w_002_607);
  nand2 I004_014(w_004_014, w_003_013, w_003_081);
  nand2 I004_015(w_004_015, w_001_019, w_001_017);
  or2  I004_016(w_004_016, w_002_079, w_001_010);
  nand2 I004_017(w_004_017, w_002_030, w_001_017);
  nand2 I004_019(w_004_019, w_000_349, w_001_009);
  and2 I004_020(w_004_020, w_000_493, w_001_012);
  not1 I004_021(w_004_021, w_001_017);
  and2 I004_022(w_004_022, w_002_011, w_002_008);
  not1 I004_023(w_004_023, w_003_033);
  or2  I004_024(w_004_024, w_001_030, w_003_071);
  not1 I004_025(w_004_025, w_001_016);
  not1 I004_026(w_004_026, w_002_030);
  not1 I004_027(w_004_027, w_003_077);
  or2  I004_028(w_004_028, w_003_023, w_003_022);
  not1 I004_029(w_004_029, w_001_034);
  not1 I004_030(w_004_030, w_002_052);
  or2  I004_031(w_004_031, w_000_494, w_000_495);
  nand2 I004_032(w_004_032, w_001_007, w_000_496);
  and2 I004_033(w_004_033, w_003_001, w_003_011);
  and2 I004_034(w_004_034, w_001_021, w_000_357);
  or2  I004_035(w_004_035, w_003_005, w_000_456);
  nand2 I004_036(w_004_036, w_002_282, w_001_018);
  not1 I004_037(w_004_037, w_003_032);
  not1 I004_038(w_004_038, w_003_066);
  or2  I004_039(w_004_039, w_000_216, w_002_297);
  and2 I004_040(w_004_040, w_001_004, w_003_074);
  nand2 I004_041(w_004_041, w_001_031, w_003_005);
  not1 I004_042(w_004_042, w_003_022);
  nand2 I004_043(w_004_043, w_003_078, w_001_026);
  nand2 I004_044(w_004_044, w_001_009, w_002_005);
  nand2 I004_045(w_004_045, w_001_020, w_000_497);
  or2  I004_046(w_004_046, w_002_170, w_001_017);
  or2  I004_047(w_004_047, w_001_027, w_001_035);
  nand2 I004_048(w_004_048, w_000_498, w_001_001);
  not1 I004_049(w_004_049, w_000_499);
  and2 I004_050(w_004_050, w_001_026, w_003_050);
  or2  I004_051(w_004_051, w_001_023, w_000_470);
  and2 I004_052(w_004_052, w_001_010, w_001_014);
  not1 I004_053(w_004_053, w_002_439);
  nand2 I004_054(w_004_054, w_003_048, w_000_193);
  nand2 I004_055(w_004_055, w_001_018, w_001_034);
  and2 I004_056(w_004_056, w_001_034, w_000_500);
  and2 I004_057(w_004_057, w_003_029, w_002_244);
  or2  I004_058(w_004_058, w_002_002, w_001_009);
  or2  I004_059(w_004_059, w_002_075, w_003_076);
  not1 I004_060(w_004_060, w_003_055);
  not1 I004_061(w_004_061, w_003_055);
  not1 I004_062(w_004_062, w_000_203);
  nand2 I004_063(w_004_063, w_001_019, w_000_501);
  nand2 I004_064(w_004_064, w_003_062, w_002_145);
  nand2 I004_065(w_004_065, w_002_386, w_001_032);
  nand2 I004_066(w_004_066, w_001_026, w_001_034);
  or2  I004_067(w_004_067, w_001_026, w_000_502);
  and2 I004_068(w_004_068, w_003_075, w_002_472);
  not1 I004_069(w_004_069, w_001_000);
  or2  I004_070(w_004_070, w_002_353, w_000_141);
  not1 I004_071(w_004_071, w_002_638);
  or2  I004_072(w_004_072, w_000_224, w_003_027);
  not1 I004_074(w_004_074, w_002_406);
  not1 I004_075(w_004_075, w_003_076);
  not1 I004_076(w_004_076, w_002_009);
  not1 I004_077(w_004_077, w_000_118);
  nand2 I004_078(w_004_078, w_001_003, w_000_189);
  not1 I004_079(w_004_079, w_003_022);
  nand2 I004_081(w_004_081, w_000_379, w_001_027);
  nand2 I004_082(w_004_082, w_003_015, w_001_025);
  not1 I004_083(w_004_083, w_000_212);
  or2  I004_084(w_004_084, w_001_020, w_001_035);
  or2  I004_085(w_004_085, w_003_072, w_001_007);
  not1 I004_086(w_004_086, w_000_505);
  not1 I004_087(w_004_087, w_001_011);
  nand2 I004_088(w_004_088, w_000_506, w_000_384);
  and2 I004_089(w_004_089, w_001_029, w_003_023);
  or2  I004_090(w_004_090, w_001_034, w_001_035);
  nand2 I004_091(w_004_091, w_002_587, w_001_029);
  and2 I004_092(w_004_092, w_000_507, w_002_088);
  nand2 I004_093(w_004_093, w_002_280, w_002_159);
  and2 I004_094(w_004_094, w_001_016, w_003_007);
  and2 I004_095(w_004_095, w_003_015, w_003_017);
  not1 I004_096(w_004_096, w_000_472);
  or2  I004_097(w_004_097, w_001_003, w_000_179);
  or2  I004_098(w_004_098, w_001_006, w_001_017);
  not1 I004_099(w_004_099, w_003_046);
  not1 I004_100(w_004_100, w_002_678);
  and2 I004_101(w_004_101, w_001_018, w_001_002);
  or2  I004_102(w_004_102, w_003_062, w_000_425);
  or2  I004_103(w_004_103, w_003_004, w_001_035);
  or2  I004_104(w_004_104, w_003_024, w_001_013);
  or2  I004_105(w_004_105, w_003_081, w_003_038);
  not1 I004_106(w_004_106, w_002_606);
  and2 I004_107(w_004_107, w_000_485, w_000_154);
  nand2 I004_108(w_004_108, w_001_008, w_001_000);
  or2  I004_109(w_004_109, w_001_019, w_002_304);
  not1 I004_110(w_004_110, w_003_040);
  nand2 I004_111(w_004_111, w_002_540, w_000_508);
  not1 I004_113(w_004_113, w_003_010);
  not1 I004_114(w_004_114, w_003_035);
  not1 I004_115(w_004_115, w_001_024);
  and2 I004_116(w_004_116, w_001_034, w_000_510);
  or2  I004_117(w_004_117, w_002_024, w_002_300);
  nand2 I004_118(w_004_118, w_001_002, w_002_481);
  and2 I004_119(w_004_119, w_003_021, w_003_084);
  nand2 I004_120(w_004_120, w_003_039, w_002_202);
  and2 I004_121(w_004_121, w_002_129, w_003_054);
  and2 I004_122(w_004_122, w_003_046, w_000_175);
  not1 I004_123(w_004_123, w_002_614);
  not1 I004_124(w_004_124, w_000_114);
  not1 I004_125(w_004_125, w_001_002);
  and2 I004_126(w_004_126, w_003_044, w_003_013);
  and2 I004_128(w_004_128, w_003_003, w_002_528);
  and2 I004_129(w_004_129, w_001_012, w_003_061);
  or2  I004_130(w_004_130, w_002_100, w_003_052);
  nand2 I004_131(w_004_131, w_003_059, w_001_029);
  or2  I004_132(w_004_132, w_001_024, w_003_050);
  not1 I004_133(w_004_133, w_000_511);
  nand2 I004_134(w_004_134, w_001_014, w_003_047);
  and2 I004_135(w_004_135, w_001_028, w_000_327);
  not1 I004_136(w_004_136, w_003_048);
  nand2 I004_137(w_004_137, w_001_014, w_003_017);
  and2 I004_138(w_004_138, w_002_393, w_001_023);
  not1 I004_139(w_004_139, w_002_487);
  or2  I004_140(w_004_140, w_002_633, w_001_000);
  or2  I004_141(w_004_141, w_003_047, w_000_399);
  and2 I004_142(w_004_142, w_002_612, w_000_365);
  not1 I004_143(w_004_143, w_003_050);
  not1 I004_144(w_004_144, w_000_512);
  or2  I004_145(w_004_145, w_002_272, w_003_039);
  or2  I004_146(w_004_146, w_003_051, w_000_513);
  not1 I004_147(w_004_147, w_002_056);
  and2 I004_148(w_004_148, w_003_064, w_003_016);
  or2  I004_149(w_004_149, w_002_515, w_003_013);
  nand2 I004_150(w_004_150, w_000_514, w_002_134);
  nand2 I004_151(w_004_151, w_003_032, w_000_515);
  not1 I004_152(w_004_152, w_000_249);
  nand2 I004_153(w_004_153, w_003_022, w_003_077);
  or2  I004_154(w_004_154, w_002_013, w_001_028);
  not1 I004_155(w_004_155, w_000_037);
  and2 I004_156(w_004_156, w_002_552, w_003_062);
  and2 I004_157(w_004_157, w_000_067, w_002_166);
  not1 I004_158(w_004_158, w_001_035);
  nand2 I004_159(w_004_159, w_003_054, w_003_064);
  not1 I004_160(w_004_160, w_002_066);
  or2  I004_161(w_004_161, w_003_006, w_003_008);
  and2 I004_162(w_004_162, w_001_029, w_000_516);
  nand2 I004_163(w_004_163, w_003_009, w_003_078);
  not1 I004_164(w_004_164, w_003_037);
  or2  I004_165(w_004_165, w_001_035, w_002_658);
  or2  I004_166(w_004_166, w_001_012, w_000_517);
  not1 I004_167(w_004_167, w_002_220);
  and2 I004_168(w_004_168, w_001_006, w_003_076);
  and2 I004_169(w_004_169, w_000_518, w_000_519);
  or2  I004_170(w_004_170, w_003_035, w_000_056);
  nand2 I004_171(w_004_171, w_003_008, w_000_409);
  or2  I004_172(w_004_172, w_003_024, w_002_056);
  nand2 I004_173(w_004_173, w_002_298, w_002_616);
  not1 I004_174(w_004_174, w_002_070);
  or2  I004_175(w_004_175, w_001_006, w_001_033);
  not1 I004_176(w_004_176, w_002_328);
  and2 I004_177(w_004_177, w_001_036, w_000_345);
  or2  I004_178(w_004_178, w_000_520, w_001_024);
  not1 I004_179(w_004_179, w_000_324);
  or2  I004_180(w_004_180, w_001_007, w_003_021);
  or2  I004_181(w_004_181, w_000_249, w_003_053);
  not1 I004_182(w_004_182, w_001_036);
  and2 I004_183(w_004_183, w_003_005, w_002_703);
  or2  I004_184(w_004_184, w_003_074, w_001_023);
  not1 I004_185(w_004_185, w_001_036);
  nand2 I004_186(w_004_186, w_002_024, w_000_318);
  or2  I004_187(w_004_187, w_001_026, w_001_022);
  nand2 I004_188(w_004_188, w_001_012, w_003_066);
  not1 I004_190(w_004_190, w_001_019);
  nand2 I004_191(w_004_191, w_001_011, w_001_005);
  or2  I004_192(w_004_192, w_002_296, w_001_004);
  and2 I004_193(w_004_193, w_001_026, w_002_194);
  or2  I004_194(w_004_194, w_003_076, w_001_035);
  nand2 I004_195(w_004_195, w_000_521, w_002_028);
  and2 I004_196(w_004_196, w_002_315, w_003_010);
  or2  I004_197(w_004_197, w_002_572, w_001_021);
  not1 I004_198(w_004_198, w_002_022);
  not1 I004_199(w_004_199, w_003_038);
  nand2 I004_200(w_004_200, w_000_182, w_001_035);
  and2 I004_201(w_004_201, w_000_432, w_001_027);
  nand2 I004_202(w_004_202, w_001_024, w_002_549);
  nand2 I004_203(w_004_203, w_000_416, w_002_495);
  or2  I004_204(w_004_204, w_001_028, w_002_212);
  not1 I004_205(w_004_205, w_001_035);
  or2  I004_206(w_004_206, w_000_522, w_000_245);
  and2 I004_207(w_004_207, w_001_017, w_000_385);
  and2 I004_208(w_004_208, w_001_001, w_003_020);
  and2 I004_209(w_004_209, w_001_032, w_003_053);
  nand2 I004_210(w_004_210, w_002_101, w_000_447);
  or2  I004_211(w_004_211, w_003_041, w_003_039);
  not1 I004_212(w_004_212, w_000_160);
  nand2 I004_213(w_004_213, w_000_523, w_003_053);
  or2  I004_214(w_004_214, w_003_063, w_001_011);
  nand2 I004_215(w_004_215, w_000_178, w_003_061);
  or2  I004_216(w_004_216, w_003_041, w_000_069);
  and2 I004_217(w_004_217, w_001_031, w_001_003);
  nand2 I004_218(w_004_218, w_001_019, w_001_001);
  and2 I004_219(w_004_219, w_001_009, w_002_000);
  nand2 I004_220(w_004_220, w_003_065, w_002_696);
  and2 I004_221(w_004_221, w_001_023, w_003_022);
  not1 I004_222(w_004_222, w_000_008);
  not1 I004_223(w_004_223, w_001_022);
  not1 I004_224(w_004_224, w_002_497);
  and2 I004_225(w_004_225, w_002_328, w_001_030);
  not1 I004_226(w_004_226, w_002_686);
  nand2 I004_227(w_004_227, w_000_056, w_003_034);
  nand2 I004_228(w_004_228, w_003_032, w_003_011);
  nand2 I004_229(w_004_229, w_000_027, w_000_524);
  nand2 I004_230(w_004_230, w_000_204, w_000_473);
  nand2 I004_231(w_004_231, w_002_522, w_003_000);
  nand2 I004_232(w_004_232, w_000_366, w_001_004);
  nand2 I004_235(w_004_235, w_000_525, w_002_009);
  nand2 I004_236(w_004_236, w_001_025, w_003_045);
  nand2 I004_237(w_004_237, w_002_496, w_001_004);
  or2  I004_238(w_004_238, w_000_526, w_003_079);
  and2 I004_239(w_004_239, w_000_527, w_003_082);
  or2  I004_240(w_004_240, w_002_015, w_000_451);
  nand2 I004_241(w_004_241, w_003_018, w_000_029);
  and2 I004_242(w_004_242, w_003_082, w_002_594);
  and2 I004_243(w_004_243, w_001_025, w_001_034);
  not1 I004_244(w_004_244, w_002_651);
  and2 I004_245(w_004_245, w_001_033, w_000_462);
  not1 I004_246(w_004_246, w_003_011);
  nand2 I004_247(w_004_247, w_001_003, w_003_080);
  not1 I004_248(w_004_248, w_002_415);
  not1 I004_249(w_004_249, w_003_077);
  or2  I004_250(w_004_250, w_001_002, w_000_194);
  or2  I004_252(w_004_252, w_000_395, w_002_589);
  nand2 I004_253(w_004_253, w_000_035, w_002_656);
  not1 I004_254(w_004_254, w_003_064);
  or2  I004_255(w_004_255, w_003_006, w_003_083);
  and2 I004_256(w_004_256, w_002_307, w_002_003);
  or2  I004_257(w_004_257, w_002_109, w_000_083);
  not1 I004_259(w_004_259, w_000_399);
  or2  I004_260(w_004_260, w_000_434, w_000_001);
  and2 I004_261(w_004_261, w_003_065, w_001_015);
  not1 I004_262(w_004_262, w_000_390);
  nand2 I004_263(w_004_263, w_002_697, w_001_001);
  not1 I004_264(w_004_264, w_003_079);
  not1 I004_265(w_004_265, w_002_075);
  nand2 I004_266(w_004_266, w_000_145, w_001_010);
  or2  I004_267(w_004_267, w_000_400, w_001_015);
  and2 I004_268(w_004_268, w_002_374, w_003_002);
  nand2 I004_269(w_004_269, w_002_537, w_003_047);
  and2 I004_270(w_004_270, w_001_029, w_001_023);
  nand2 I004_271(w_004_271, w_000_528, w_001_030);
  or2  I004_272(w_004_272, w_001_004, w_002_622);
  or2  I004_273(w_004_273, w_003_060, w_001_015);
  or2  I004_274(w_004_274, w_001_003, w_000_405);
  not1 I004_275(w_004_275, w_003_062);
  and2 I004_276(w_004_276, w_003_037, w_000_456);
  or2  I004_277(w_004_277, w_002_059, w_001_024);
  or2  I004_278(w_004_278, w_002_065, w_003_057);
  and2 I004_279(w_004_279, w_001_032, w_001_035);
  or2  I004_280(w_004_280, w_003_031, w_002_016);
  or2  I004_281(w_004_281, w_002_685, w_000_186);
  or2  I004_282(w_004_282, w_000_177, w_001_035);
  or2  I004_283(w_004_283, w_002_342, w_001_001);
  or2  I004_284(w_004_284, w_002_222, w_002_101);
  or2  I004_285(w_004_285, w_002_391, w_003_012);
  and2 I004_286(w_004_286, w_000_026, w_002_583);
  nand2 I004_287(w_004_287, w_003_073, w_000_287);
  nand2 I004_288(w_004_288, w_001_008, w_000_346);
  and2 I004_289(w_004_289, w_002_065, w_002_127);
  and2 I004_290(w_004_290, w_003_081, w_002_517);
  nand2 I004_291(w_004_291, w_000_529, w_002_231);
  nand2 I004_292(w_004_292, w_002_104, w_001_027);
  nand2 I004_293(w_004_293, w_000_235, w_000_441);
  nand2 I004_294(w_004_294, w_000_530, w_002_684);
  or2  I004_295(w_004_295, w_002_302, w_002_053);
  or2  I004_296(w_004_296, w_002_516, w_003_059);
  not1 I004_297(w_004_297, w_002_057);
  and2 I004_299(w_004_299, w_002_418, w_003_008);
  not1 I004_301(w_004_301, w_003_021);
  nand2 I004_302(w_004_302, w_001_020, w_001_036);
  or2  I004_304(w_004_304, w_001_005, w_002_601);
  not1 I004_305(w_004_305, w_003_030);
  not1 I004_307(w_004_307, w_003_024);
  not1 I004_308(w_004_308, w_003_049);
  not1 I004_309(w_004_309, w_001_012);
  not1 I004_310(w_004_310, w_000_533);
  or2  I004_311(w_004_311, w_001_005, w_002_584);
  and2 I004_314(w_004_314, w_000_468, w_003_021);
  or2  I004_315(w_004_315, w_001_022, w_000_151);
  nand2 I004_316(w_004_316, w_000_493, w_000_418);
  nand2 I004_317(w_004_317, w_000_202, w_001_035);
  nand2 I004_319(w_004_319, w_001_030, w_000_146);
  not1 I004_320(w_004_320, w_000_534);
  nand2 I004_321(w_004_321, w_001_016, w_003_045);
  or2  I004_322(w_004_322, w_003_081, w_002_543);
  not1 I004_325(w_004_325, w_002_547);
  or2  I004_326(w_004_326, w_000_535, w_001_034);
  or2  I004_328(w_004_328, w_002_509, w_002_017);
  nand2 I004_329(w_004_329, w_000_112, w_003_026);
  and2 I004_330(w_004_330, w_002_340, w_002_146);
  or2  I004_331(w_004_331, w_001_014, w_003_020);
  and2 I004_332(w_004_332, w_001_010, w_002_498);
  not1 I004_333(w_004_333, w_001_014);
  and2 I004_335(w_004_335, w_000_175, w_003_024);
  nand2 I004_336(w_004_336, w_002_657, w_000_536);
  or2  I004_337(w_004_337, w_002_467, w_003_056);
  and2 I004_338(w_004_338, w_002_211, w_001_028);
  not1 I004_340(w_004_340, w_002_120);
  or2  I004_341(w_004_341, w_000_278, w_001_006);
  not1 I004_343(w_004_343, w_001_026);
  nand2 I004_344(w_004_344, w_003_027, w_002_638);
  nand2 I004_345(w_004_345, w_001_032, w_000_228);
  or2  I004_346(w_004_346, w_003_000, w_003_067);
  and2 I004_347(w_004_347, w_001_016, w_001_006);
  nand2 I004_348(w_004_348, w_002_618, w_000_366);
  nand2 I004_349(w_004_349, w_001_017, w_001_025);
  and2 I004_350(w_004_350, w_000_538, w_003_025);
  and2 I004_351(w_004_351, w_003_045, w_002_543);
  and2 I004_352(w_004_352, w_003_031, w_003_058);
  nand2 I004_353(w_004_353, w_003_035, w_003_053);
  not1 I004_354(w_004_354, w_002_227);
  and2 I004_355(w_004_355, w_003_061, w_003_029);
  and2 I004_357(w_004_357, w_003_081, w_000_486);
  and2 I004_359(w_004_359, w_003_076, w_003_067);
  and2 I004_360(w_004_360, w_003_012, w_002_361);
  nand2 I004_361(w_004_361, w_003_074, w_001_007);
  or2  I004_362(w_004_362, w_000_227, w_000_256);
  and2 I004_363(w_004_363, w_000_027, w_000_449);
  or2  I004_364(w_004_364, w_000_143, w_002_580);
  or2  I004_365(w_004_365, w_003_060, w_002_250);
  nand2 I004_366(w_004_366, w_002_017, w_003_033);
  nand2 I004_367(w_004_367, w_002_304, w_003_054);
  not1 I004_368(w_004_368, w_000_156);
  or2  I004_369(w_004_369, w_000_540, w_001_002);
  nand2 I004_370(w_004_370, w_001_021, w_000_101);
  or2  I004_371(w_004_371, w_003_064, w_003_012);
  not1 I004_372(w_004_372, w_001_028);
  or2  I004_373(w_004_373, w_003_084, w_000_004);
  or2  I004_374(w_004_374, w_002_660, w_000_286);
  nand2 I004_375(w_004_375, w_001_018, w_000_069);
  nand2 I004_376(w_004_376, w_002_030, w_003_008);
  and2 I004_377(w_004_377, w_003_037, w_002_678);
  nand2 I004_378(w_004_378, w_001_030, w_001_017);
  or2  I004_379(w_004_379, w_002_173, w_003_052);
  not1 I004_380(w_004_380, w_000_541);
  or2  I004_382(w_004_382, w_001_026, w_002_031);
  or2  I004_383(w_004_383, w_000_325, w_000_403);
  not1 I004_384(w_004_384, w_000_320);
  and2 I004_386(w_004_386, w_003_016, w_002_112);
  nand2 I004_387(w_004_387, w_000_290, w_003_015);
  or2  I004_388(w_004_388, w_003_065, w_002_061);
  not1 I004_389(w_004_389, w_000_268);
  nand2 I004_390(w_004_390, w_000_542, w_000_192);
  nand2 I004_391(w_004_391, w_000_064, w_003_003);
  and2 I004_392(w_004_392, w_000_349, w_000_299);
  or2  I004_393(w_004_393, w_003_084, w_000_543);
  not1 I004_394(w_004_394, w_003_003);
  nand2 I004_395(w_004_395, w_003_033, w_002_016);
  not1 I004_396(w_004_396, w_002_636);
  not1 I004_397(w_004_397, w_003_016);
  not1 I004_398(w_004_398, w_003_008);
  not1 I004_399(w_004_399, w_003_036);
  and2 I004_400(w_004_400, w_003_022, w_002_128);
  and2 I004_401(w_004_401, w_003_023, w_000_544);
  not1 I004_402(w_004_402, w_003_061);
  not1 I004_405(w_004_405, w_000_545);
  and2 I004_406(w_004_406, w_002_149, w_001_035);
  and2 I004_407(w_004_407, w_001_018, w_000_202);
  not1 I004_408(w_004_408, w_000_331);
  not1 I004_409(w_004_409, w_003_083);
  not1 I004_410(w_004_410, w_001_026);
  or2  I004_411(w_004_411, w_000_357, w_000_508);
  not1 I004_413(w_004_413, w_002_613);
  and2 I004_414(w_004_414, w_003_015, w_000_546);
  nand2 I004_415(w_004_415, w_000_547, w_002_327);
  and2 I004_416(w_004_416, w_001_009, w_003_024);
  and2 I004_418(w_004_418, w_000_253, w_001_023);
  nand2 I004_419(w_004_419, w_002_564, w_001_007);
  or2  I004_420(w_004_420, w_001_013, w_003_056);
  and2 I004_421(w_004_421, w_002_421, w_000_248);
  not1 I004_423(w_004_423, w_000_003);
  or2  I004_424(w_004_424, w_001_011, w_001_026);
  or2  I004_425(w_004_425, w_002_600, w_000_548);
  and2 I004_426(w_004_426, w_001_004, w_001_024);
  or2  I004_427(w_004_427, w_000_549, w_001_029);
  or2  I004_428(w_004_428, w_001_032, w_001_002);
  or2  I004_429(w_004_429, w_003_029, w_003_046);
  not1 I004_431(w_004_431, w_001_015);
  not1 I004_432(w_004_432, w_002_396);
  nand2 I004_433(w_004_433, w_003_049, w_000_002);
  not1 I004_434(w_004_434, w_001_015);
  nand2 I004_435(w_004_435, w_000_094, w_000_507);
  and2 I004_436(w_004_436, w_001_029, w_003_045);
  nand2 I004_437(w_004_437, w_002_684, w_003_039);
  and2 I004_438(w_004_438, w_000_429, w_002_668);
  nand2 I004_439(w_004_439, w_000_264, w_002_127);
  or2  I004_440(w_004_440, w_003_044, w_003_017);
  nand2 I004_441(w_004_441, w_002_176, w_001_002);
  and2 I004_443(w_004_443, w_003_068, w_000_143);
  not1 I004_444(w_004_444, w_001_018);
  nand2 I004_445(w_004_445, w_003_071, w_002_439);
  nand2 I004_446(w_004_446, w_001_007, w_000_550);
  and2 I004_447(w_004_447, w_003_030, w_003_058);
  and2 I004_448(w_004_448, w_000_163, w_003_021);
  not1 I004_449(w_004_449, w_003_019);
  not1 I004_450(w_004_450, w_003_002);
  nand2 I004_451(w_004_451, w_002_039, w_000_337);
  not1 I004_452(w_004_452, w_003_069);
  or2  I004_453(w_004_453, w_002_296, w_002_000);
  or2  I004_454(w_004_454, w_002_512, w_000_390);
  nand2 I004_455(w_004_455, w_002_658, w_000_551);
  or2  I004_456(w_004_456, w_002_048, w_001_018);
  not1 I004_457(w_004_457, w_000_482);
  and2 I004_459(w_004_459, w_000_552, w_001_034);
  or2  I004_460(w_004_460, w_003_051, w_002_341);
  or2  I004_462(w_004_462, w_003_070, w_002_357);
  not1 I004_463(w_004_463, w_003_083);
  and2 I004_464(w_004_464, w_003_020, w_002_229);
  or2  I004_465(w_004_465, w_003_052, w_001_020);
  or2  I004_466(w_004_466, w_002_082, w_002_657);
  or2  I004_468(w_004_468, w_000_403, w_002_323);
  or2  I004_469(w_004_469, w_000_232, w_003_069);
  or2  I004_470(w_004_470, w_000_553, w_001_017);
  or2  I004_471(w_004_471, w_002_425, w_002_599);
  or2  I004_472(w_004_472, w_003_000, w_000_554);
  not1 I004_473(w_004_473, w_001_029);
  and2 I004_474(w_004_474, w_002_369, w_001_035);
  or2  I004_476(w_004_476, w_002_043, w_003_065);
  nand2 I004_477(w_004_477, w_000_484, w_000_555);
  or2  I004_478(w_004_478, w_002_085, w_003_062);
  not1 I004_479(w_004_479, w_003_054);
  and2 I004_480(w_004_480, w_000_556, w_000_223);
  nand2 I004_482(w_004_482, w_003_030, w_000_289);
  nand2 I004_484(w_004_484, w_002_461, w_000_132);
  and2 I004_486(w_004_486, w_002_481, w_000_558);
  nand2 I004_487(w_004_487, w_000_150, w_002_593);
  nand2 I004_488(w_004_488, w_003_031, w_002_078);
  or2  I004_489(w_004_489, w_003_024, w_000_462);
  not1 I004_490(w_004_490, w_002_190);
  or2  I004_491(w_004_491, w_000_559, w_001_009);
  not1 I004_492(w_004_492, w_001_031);
  not1 I004_493(w_004_493, w_003_031);
  and2 I004_495(w_004_495, w_001_033, w_003_069);
  not1 I004_496(w_004_496, w_001_000);
  or2  I004_497(w_004_497, w_000_560, w_000_561);
  or2  I004_498(w_004_498, w_002_175, w_001_020);
  and2 I004_499(w_004_499, w_001_011, w_001_014);
  not1 I004_500(w_004_500, w_001_018);
  or2  I004_501(w_004_501, w_003_062, w_000_060);
  nand2 I004_502(w_004_502, w_001_019, w_002_340);
  not1 I004_503(w_004_503, w_003_073);
  and2 I004_505(w_004_505, w_002_252, w_002_459);
  and2 I004_506(w_004_506, w_003_020, w_002_114);
  or2  I004_507(w_004_507, w_003_064, w_002_282);
  nand2 I004_508(w_004_508, w_002_342, w_002_340);
  nand2 I005_000(w_005_000, w_000_273, w_004_032);
  or2  I005_001(w_005_001, w_001_026, w_002_243);
  or2  I005_002(w_005_002, w_003_013, w_000_253);
  or2  I005_003(w_005_003, w_002_226, w_004_071);
  and2 I005_004(w_005_004, w_002_162, w_000_441);
  and2 I005_005(w_005_005, w_002_240, w_003_052);
  or2  I005_006(w_005_006, w_003_067, w_003_084);
  or2  I005_007(w_005_007, w_003_075, w_002_402);
  nand2 I005_008(w_005_008, w_003_040, w_003_015);
  not1 I005_009(w_005_009, w_001_023);
  and2 I005_010(w_005_010, w_000_563, w_003_007);
  or2  I005_011(w_005_011, w_000_001, w_001_010);
  or2  I005_012(w_005_012, w_004_246, w_001_010);
  and2 I005_013(w_005_013, w_001_031, w_004_029);
  or2  I005_014(w_005_014, w_003_056, w_000_426);
  or2  I005_015(w_005_015, w_001_023, w_004_237);
  and2 I005_016(w_005_016, w_002_207, w_002_457);
  nand2 I005_017(w_005_017, w_004_089, w_003_031);
  and2 I005_018(w_005_018, w_004_150, w_004_227);
  or2  I005_019(w_005_019, w_004_343, w_000_144);
  not1 I005_020(w_005_020, w_003_057);
  nand2 I005_021(w_005_021, w_003_036, w_001_032);
  and2 I005_022(w_005_022, w_001_016, w_001_007);
  not1 I005_023(w_005_023, w_003_032);
  or2  I005_024(w_005_024, w_000_438, w_003_071);
  not1 I005_025(w_005_025, w_004_283);
  and2 I005_026(w_005_026, w_001_031, w_001_020);
  or2  I005_027(w_005_027, w_000_098, w_001_035);
  or2  I005_028(w_005_028, w_001_016, w_004_293);
  and2 I005_029(w_005_029, w_000_531, w_001_020);
  or2  I005_030(w_005_030, w_002_406, w_001_027);
  and2 I005_031(w_005_031, w_001_012, w_000_425);
  or2  I005_032(w_005_032, w_000_098, w_004_249);
  not1 I005_033(w_005_033, w_004_411);
  and2 I005_034(w_005_034, w_000_564, w_000_403);
  nand2 I005_035(w_005_035, w_000_565, w_004_432);
  and2 I005_036(w_005_036, w_001_005, w_001_021);
  and2 I005_037(w_005_037, w_003_022, w_003_026);
  and2 I005_038(w_005_038, w_000_417, w_000_566);
  nand2 I005_039(w_005_039, w_001_025, w_004_090);
  not1 I005_040(w_005_040, w_001_011);
  not1 I005_041(w_005_041, w_004_096);
  or2  I005_042(w_005_042, w_001_011, w_003_040);
  and2 I005_043(w_005_043, w_004_167, w_001_000);
  not1 I005_044(w_005_044, w_001_007);
  nand2 I005_046(w_005_046, w_001_004, w_002_383);
  and2 I005_047(w_005_047, w_002_594, w_003_002);
  and2 I005_048(w_005_048, w_002_608, w_004_045);
  and2 I005_049(w_005_049, w_002_681, w_004_503);
  not1 I005_050(w_005_050, w_002_577);
  and2 I005_051(w_005_051, w_000_395, w_002_354);
  or2  I005_052(w_005_052, w_001_032, w_004_282);
  nand2 I005_053(w_005_053, w_001_033, w_001_004);
  and2 I005_054(w_005_054, w_004_039, w_000_567);
  or2  I005_055(w_005_055, w_004_239, w_002_664);
  not1 I005_056(w_005_056, w_001_016);
  or2  I005_057(w_005_057, w_000_049, w_002_575);
  and2 I005_058(w_005_058, w_002_129, w_000_435);
  not1 I005_059(w_005_059, w_004_269);
  or2  I005_060(w_005_060, w_002_487, w_004_354);
  nand2 I005_061(w_005_061, w_001_030, w_001_017);
  or2  I005_062(w_005_062, w_003_056, w_000_537);
  not1 I005_063(w_005_063, w_003_031);
  nand2 I005_064(w_005_064, w_003_080, w_004_193);
  not1 I005_065(w_005_065, w_001_015);
  and2 I005_066(w_005_066, w_001_005, w_001_024);
  or2  I005_067(w_005_067, w_000_568, w_002_074);
  or2  I005_068(w_005_068, w_000_090, w_000_569);
  and2 I005_069(w_005_069, w_003_072, w_003_062);
  nand2 I005_070(w_005_070, w_002_059, w_003_027);
  and2 I005_071(w_005_071, w_002_538, w_003_009);
  nand2 I005_072(w_005_072, w_000_432, w_002_293);
  not1 I005_073(w_005_073, w_000_570);
  and2 I005_074(w_005_074, w_000_264, w_002_048);
  not1 I005_075(w_005_075, w_004_096);
  not1 I005_076(w_005_076, w_000_571);
  not1 I005_077(w_005_077, w_002_026);
  and2 I005_078(w_005_078, w_001_019, w_002_045);
  not1 I005_079(w_005_079, w_000_215);
  not1 I005_080(w_005_080, w_003_043);
  nand2 I005_081(w_005_081, w_001_032, w_003_036);
  nand2 I005_083(w_005_083, w_001_005, w_002_154);
  nand2 I005_084(w_005_084, w_002_600, w_004_232);
  and2 I005_085(w_005_085, w_003_035, w_004_170);
  and2 I005_086(w_005_086, w_000_385, w_002_150);
  nand2 I005_087(w_005_087, w_003_031, w_004_451);
  not1 I005_088(w_005_088, w_000_405);
  and2 I005_089(w_005_089, w_000_572, w_004_476);
  nand2 I005_090(w_005_090, w_001_034, w_003_048);
  not1 I005_091(w_005_091, w_003_052);
  not1 I005_092(w_005_092, w_003_002);
  or2  I005_093(w_005_093, w_003_058, w_001_002);
  and2 I005_094(w_005_094, w_003_061, w_003_080);
  not1 I005_095(w_005_095, w_001_015);
  not1 I005_096(w_005_096, w_001_018);
  nand2 I005_097(w_005_097, w_001_017, w_000_005);
  or2  I005_098(w_005_098, w_003_021, w_004_132);
  nand2 I005_099(w_005_099, w_001_012, w_004_449);
  and2 I005_100(w_005_100, w_004_252, w_000_573);
  not1 I005_101(w_005_101, w_003_045);
  and2 I005_102(w_005_102, w_000_257, w_000_362);
  nand2 I005_103(w_005_103, w_004_192, w_001_027);
  or2  I005_104(w_005_104, w_002_287, w_004_050);
  nand2 I005_105(w_005_105, w_003_074, w_004_227);
  nand2 I005_106(w_005_106, w_003_058, w_002_522);
  and2 I005_107(w_005_107, w_002_059, w_001_019);
  not1 I005_108(w_005_108, w_002_551);
  and2 I005_109(w_005_109, w_002_466, w_003_033);
  not1 I005_110(w_005_110, w_000_473);
  nand2 I005_111(w_005_111, w_002_313, w_003_004);
  and2 I005_112(w_005_112, w_004_248, w_001_009);
  and2 I005_113(w_005_113, w_001_021, w_003_066);
  or2  I005_114(w_005_114, w_003_040, w_004_071);
  and2 I005_115(w_005_115, w_003_004, w_000_574);
  not1 I005_116(w_005_116, w_004_186);
  and2 I005_117(w_005_117, w_004_211, w_004_098);
  not1 I005_118(w_005_118, w_000_102);
  nand2 I005_119(w_005_119, w_004_192, w_004_042);
  not1 I005_120(w_005_120, w_000_563);
  not1 I005_121(w_005_121, w_003_026);
  or2  I005_122(w_005_122, w_003_067, w_003_065);
  and2 I005_123(w_005_123, w_002_212, w_002_165);
  and2 I005_124(w_005_124, w_003_045, w_002_642);
  or2  I005_125(w_005_125, w_000_076, w_002_094);
  nand2 I005_126(w_005_126, w_003_032, w_000_567);
  nand2 I005_127(w_005_127, w_003_075, w_001_004);
  not1 I005_128(w_005_128, w_000_445);
  or2  I005_129(w_005_129, w_000_317, w_002_603);
  or2  I005_130(w_005_130, w_004_320, w_001_031);
  or2  I005_131(w_005_131, w_003_047, w_001_016);
  and2 I005_132(w_005_132, w_000_295, w_000_575);
  and2 I005_133(w_005_133, w_002_400, w_002_605);
  not1 I005_134(w_005_134, w_000_576);
  and2 I005_135(w_005_135, w_001_015, w_002_676);
  or2  I005_136(w_005_136, w_004_031, w_000_544);
  nand2 I005_137(w_005_137, w_003_046, w_001_003);
  not1 I005_138(w_005_138, w_004_070);
  not1 I005_139(w_005_139, w_000_365);
  not1 I005_140(w_005_140, w_000_210);
  and2 I005_141(w_005_141, w_001_026, w_000_577);
  nand2 I005_142(w_005_142, w_002_581, w_002_488);
  not1 I005_143(w_005_143, w_001_020);
  or2  I005_144(w_005_144, w_002_092, w_001_018);
  and2 I005_145(w_005_145, w_002_256, w_001_004);
  nand2 I005_146(w_005_146, w_001_023, w_000_057);
  not1 I005_147(w_005_147, w_001_008);
  not1 I005_148(w_005_148, w_004_141);
  nand2 I005_149(w_005_149, w_004_292, w_003_032);
  and2 I005_150(w_005_150, w_001_002, w_001_021);
  and2 I005_151(w_005_151, w_000_502, w_001_028);
  not1 I005_152(w_005_152, w_000_578);
  and2 I005_153(w_005_153, w_002_262, w_002_060);
  or2  I005_154(w_005_154, w_001_029, w_000_579);
  and2 I005_155(w_005_155, w_001_029, w_001_001);
  or2  I005_156(w_005_156, w_004_165, w_001_011);
  and2 I005_157(w_005_157, w_002_102, w_002_204);
  and2 I005_158(w_005_158, w_000_580, w_004_345);
  or2  I005_159(w_005_159, w_002_502, w_001_025);
  nand2 I005_160(w_005_160, w_001_035, w_001_006);
  not1 I005_161(w_005_161, w_002_045);
  nand2 I005_162(w_005_162, w_000_581, w_003_049);
  nand2 I005_163(w_005_163, w_001_030, w_003_000);
  or2  I005_164(w_005_164, w_000_374, w_002_306);
  or2  I005_165(w_005_165, w_001_018, w_004_335);
  not1 I005_166(w_005_166, w_002_190);
  or2  I005_167(w_005_167, w_000_582, w_001_026);
  nand2 I005_168(w_005_168, w_000_404, w_002_610);
  not1 I005_169(w_005_169, w_000_296);
  or2  I005_170(w_005_170, w_003_027, w_000_453);
  and2 I005_171(w_005_171, w_003_028, w_000_196);
  or2  I005_172(w_005_172, w_004_399, w_003_074);
  or2  I005_173(w_005_173, w_003_071, w_004_078);
  and2 I005_174(w_005_174, w_003_024, w_002_233);
  or2  I005_175(w_005_175, w_004_396, w_002_097);
  and2 I005_176(w_005_176, w_002_380, w_001_020);
  not1 I005_177(w_005_177, w_004_432);
  not1 I005_178(w_005_178, w_002_628);
  or2  I005_180(w_005_180, w_002_376, w_004_117);
  and2 I005_181(w_005_181, w_002_107, w_001_024);
  and2 I005_182(w_005_182, w_003_065, w_000_583);
  nand2 I005_183(w_005_183, w_002_180, w_001_005);
  not1 I005_184(w_005_184, w_003_061);
  and2 I005_185(w_005_185, w_002_036, w_001_020);
  and2 I005_186(w_005_186, w_000_584, w_003_049);
  not1 I005_187(w_005_187, w_004_178);
  nand2 I005_188(w_005_188, w_003_030, w_000_585);
  and2 I005_189(w_005_189, w_003_033, w_002_130);
  nand2 I005_190(w_005_190, w_004_153, w_001_007);
  or2  I005_191(w_005_191, w_004_400, w_000_286);
  or2  I005_192(w_005_192, w_001_006, w_002_598);
  nand2 I005_193(w_005_193, w_000_017, w_002_061);
  or2  I005_194(w_005_194, w_001_009, w_003_077);
  not1 I005_195(w_005_195, w_000_202);
  not1 I005_196(w_005_196, w_002_685);
  or2  I005_197(w_005_197, w_003_038, w_001_018);
  or2  I005_198(w_005_198, w_003_063, w_004_116);
  and2 I005_199(w_005_199, w_002_345, w_001_000);
  and2 I005_200(w_005_200, w_002_124, w_002_490);
  not1 I005_201(w_005_201, w_004_255);
  nand2 I005_202(w_005_202, w_003_022, w_002_692);
  or2  I005_204(w_005_204, w_002_273, w_000_232);
  and2 I005_205(w_005_205, w_004_349, w_000_586);
  not1 I005_206(w_005_206, w_002_459);
  not1 I005_207(w_005_207, w_001_025);
  nand2 I005_208(w_005_208, w_001_033, w_002_428);
  or2  I005_209(w_005_209, w_002_597, w_001_006);
  and2 I005_210(w_005_210, w_004_147, w_004_353);
  nand2 I005_211(w_005_211, w_004_116, w_000_351);
  nand2 I005_212(w_005_212, w_001_030, w_002_440);
  not1 I005_213(w_005_213, w_001_008);
  and2 I005_214(w_005_214, w_004_078, w_001_015);
  not1 I005_215(w_005_215, w_000_346);
  nand2 I005_216(w_005_216, w_003_071, w_000_065);
  or2  I005_218(w_005_218, w_003_057, w_001_014);
  and2 I005_219(w_005_219, w_003_049, w_002_328);
  not1 I005_220(w_005_220, w_000_332);
  nand2 I005_221(w_005_221, w_000_472, w_003_038);
  or2  I005_223(w_005_223, w_000_142, w_003_010);
  nand2 I005_224(w_005_224, w_004_285, w_001_036);
  not1 I005_225(w_005_225, w_001_023);
  not1 I005_226(w_005_226, w_004_014);
  not1 I005_227(w_005_227, w_003_038);
  not1 I005_228(w_005_228, w_003_039);
  nand2 I005_229(w_005_229, w_003_016, w_001_017);
  and2 I005_230(w_005_230, w_001_014, w_000_587);
  not1 I005_231(w_005_231, w_000_588);
  and2 I005_232(w_005_232, w_002_272, w_001_004);
  nand2 I005_233(w_005_233, w_001_018, w_000_174);
  nand2 I005_234(w_005_234, w_001_023, w_003_025);
  not1 I005_235(w_005_235, w_003_006);
  or2  I005_236(w_005_236, w_001_022, w_004_166);
  not1 I005_237(w_005_237, w_000_589);
  and2 I005_238(w_005_238, w_004_192, w_000_247);
  or2  I005_239(w_005_239, w_004_072, w_000_590);
  nand2 I005_240(w_005_240, w_001_013, w_004_020);
  nand2 I005_242(w_005_242, w_002_155, w_004_065);
  or2  I005_243(w_005_243, w_003_038, w_002_640);
  nand2 I005_244(w_005_244, w_000_155, w_002_013);
  not1 I005_245(w_005_245, w_003_007);
  not1 I005_246(w_005_246, w_003_013);
  or2  I005_247(w_005_247, w_002_130, w_004_164);
  nand2 I005_248(w_005_248, w_002_307, w_000_514);
  not1 I005_249(w_005_249, w_002_222);
  not1 I005_250(w_005_250, w_004_241);
  and2 I005_251(w_005_251, w_002_171, w_003_026);
  nand2 I005_252(w_005_252, w_000_591, w_003_038);
  not1 I005_254(w_005_254, w_001_029);
  or2  I005_255(w_005_255, w_000_137, w_003_067);
  and2 I005_256(w_005_256, w_000_525, w_004_147);
  and2 I005_257(w_005_257, w_003_025, w_001_028);
  not1 I005_259(w_005_259, w_001_015);
  not1 I005_260(w_005_260, w_003_038);
  not1 I005_261(w_005_261, w_004_040);
  and2 I005_262(w_005_262, w_002_070, w_000_039);
  and2 I005_263(w_005_263, w_004_201, w_002_370);
  not1 I005_266(w_005_266, w_003_043);
  not1 I005_267(w_005_267, w_004_276);
  and2 I005_268(w_005_268, w_003_006, w_004_117);
  and2 I005_270(w_005_270, w_000_592, w_003_036);
  nand2 I005_271(w_005_271, w_003_019, w_004_013);
  not1 I005_272(w_005_272, w_001_005);
  and2 I005_273(w_005_273, w_001_001, w_001_032);
  and2 I005_274(w_005_274, w_000_014, w_004_140);
  or2  I005_275(w_005_275, w_000_029, w_001_016);
  or2  I005_276(w_005_276, w_003_027, w_003_078);
  not1 I005_277(w_005_277, w_001_014);
  not1 I005_278(w_005_278, w_001_017);
  not1 I005_279(w_005_279, w_004_211);
  or2  I005_280(w_005_280, w_000_449, w_001_003);
  or2  I005_281(w_005_281, w_000_593, w_002_051);
  nand2 I005_282(w_005_282, w_000_304, w_004_011);
  and2 I005_283(w_005_283, w_003_004, w_001_004);
  and2 I005_285(w_005_285, w_003_044, w_000_594);
  or2  I005_286(w_005_286, w_001_005, w_001_010);
  or2  I005_287(w_005_287, w_004_397, w_002_679);
  and2 I005_288(w_005_288, w_001_024, w_002_316);
  nand2 I005_289(w_005_289, w_003_073, w_002_176);
  and2 I005_290(w_005_290, w_003_047, w_004_314);
  and2 I005_291(w_005_291, w_003_005, w_001_006);
  and2 I005_292(w_005_292, w_004_421, w_001_010);
  nand2 I005_293(w_005_293, w_001_019, w_001_030);
  and2 I005_294(w_005_294, w_002_471, w_001_004);
  and2 I005_295(w_005_295, w_002_270, w_000_174);
  nand2 I005_296(w_005_296, w_004_284, w_001_017);
  nand2 I005_297(w_005_297, w_001_029, w_001_014);
  nand2 I005_298(w_005_298, w_004_123, w_004_136);
  nand2 I005_299(w_005_299, w_002_324, w_003_053);
  or2  I005_300(w_005_300, w_001_029, w_002_274);
  or2  I005_301(w_005_301, w_002_477, w_003_012);
  nand2 I005_302(w_005_302, w_002_085, w_003_023);
  and2 I005_303(w_005_303, w_001_002, w_001_016);
  nand2 I005_304(w_005_304, w_004_231, w_003_013);
  nand2 I005_305(w_005_305, w_000_177, w_000_519);
  not1 I005_306(w_005_306, w_001_023);
  nand2 I005_307(w_005_307, w_004_047, w_004_281);
  not1 I005_308(w_005_308, w_002_526);
  or2  I005_309(w_005_309, w_002_075, w_002_110);
  nand2 I005_310(w_005_310, w_003_002, w_003_022);
  and2 I005_311(w_005_311, w_002_026, w_003_067);
  or2  I005_312(w_005_312, w_003_075, w_003_079);
  nand2 I005_313(w_005_313, w_001_011, w_002_370);
  nand2 I005_314(w_005_314, w_001_019, w_004_035);
  not1 I005_315(w_005_315, w_003_072);
  or2  I005_316(w_005_316, w_003_013, w_002_048);
  nand2 I005_317(w_005_317, w_000_581, w_004_359);
  nand2 I005_318(w_005_318, w_004_256, w_001_034);
  or2  I006_000(w_006_000, w_002_374, w_001_027);
  and2 I006_001(w_006_001, w_003_076, w_000_595);
  not1 I006_002(w_006_002, w_004_069);
  or2  I006_003(w_006_003, w_005_136, w_003_026);
  and2 I006_004(w_006_004, w_001_001, w_003_045);
  and2 I006_005(w_006_005, w_000_289, w_004_221);
  not1 I006_006(w_006_006, w_003_057);
  nand2 I006_007(w_006_007, w_004_409, w_000_564);
  or2  I006_008(w_006_008, w_002_278, w_000_145);
  and2 I006_009(w_006_009, w_002_013, w_001_004);
  or2  I006_010(w_006_010, w_002_529, w_002_220);
  or2  I006_011(w_006_011, w_005_064, w_001_022);
  and2 I006_012(w_006_012, w_004_027, w_004_059);
  or2  I006_013(w_006_013, w_003_060, w_000_596);
  not1 I006_014(w_006_014, w_004_184);
  and2 I006_015(w_006_015, w_004_329, w_000_000);
  not1 I006_016(w_006_016, w_000_597);
  and2 I006_017(w_006_017, w_002_436, w_004_148);
  not1 I006_018(w_006_018, w_001_014);
  nand2 I006_019(w_006_019, w_005_276, w_001_015);
  or2  I006_020(w_006_020, w_001_022, w_002_042);
  and2 I006_021(w_006_021, w_004_134, w_004_008);
  and2 I006_022(w_006_022, w_000_400, w_001_001);
  not1 I006_023(w_006_023, w_001_020);
  not1 I006_024(w_006_024, w_001_008);
  and2 I006_025(w_006_025, w_000_598, w_000_599);
  not1 I006_026(w_006_026, w_005_138);
  nand2 I006_027(w_006_027, w_002_643, w_000_446);
  or2  I006_028(w_006_028, w_003_027, w_000_303);
  nand2 I006_029(w_006_029, w_002_580, w_005_038);
  or2  I006_030(w_006_030, w_002_597, w_002_304);
  nand2 I006_031(w_006_031, w_001_016, w_002_331);
  nand2 I006_032(w_006_032, w_000_600, w_003_049);
  and2 I006_033(w_006_033, w_004_159, w_001_011);
  nand2 I006_034(w_006_034, w_003_034, w_002_513);
  nand2 I006_035(w_006_035, w_001_022, w_005_313);
  not1 I006_036(w_006_036, w_000_601);
  nand2 I006_037(w_006_037, w_000_272, w_000_116);
  or2  I006_038(w_006_038, w_000_447, w_002_636);
  not1 I006_039(w_006_039, w_005_226);
  not1 I006_040(w_006_040, w_001_021);
  not1 I006_041(w_006_041, w_004_253);
  nand2 I006_042(w_006_042, w_002_113, w_002_534);
  not1 I006_043(w_006_043, w_003_022);
  not1 I006_044(w_006_044, w_003_043);
  nand2 I006_045(w_006_045, w_000_362, w_005_140);
  not1 I006_047(w_006_047, w_002_622);
  and2 I006_048(w_006_048, w_005_048, w_000_447);
  nand2 I006_049(w_006_049, w_002_485, w_000_603);
  nand2 I006_051(w_006_051, w_005_289, w_002_001);
  nand2 I006_052(w_006_052, w_003_021, w_000_476);
  not1 I006_053(w_006_053, w_001_013);
  and2 I006_054(w_006_054, w_001_006, w_000_281);
  nand2 I006_055(w_006_055, w_005_280, w_001_000);
  or2  I006_056(w_006_056, w_005_104, w_005_065);
  not1 I006_057(w_006_057, w_005_162);
  or2  I006_058(w_006_058, w_005_003, w_002_032);
  or2  I006_059(w_006_059, w_003_065, w_000_139);
  nand2 I006_060(w_006_060, w_005_152, w_003_078);
  and2 I006_061(w_006_061, w_004_239, w_001_019);
  nand2 I006_062(w_006_062, w_002_010, w_003_023);
  or2  I006_063(w_006_063, w_000_065, w_004_122);
  nand2 I006_064(w_006_064, w_005_274, w_004_111);
  or2  I006_065(w_006_065, w_003_064, w_004_311);
  or2  I006_066(w_006_066, w_003_034, w_004_102);
  or2  I006_067(w_006_067, w_002_204, w_000_085);
  nand2 I006_068(w_006_068, w_000_144, w_002_693);
  and2 I006_069(w_006_069, w_005_133, w_005_139);
  or2  I006_070(w_006_070, w_004_253, w_002_090);
  and2 I006_071(w_006_071, w_004_354, w_001_010);
  or2  I006_072(w_006_072, w_002_563, w_000_374);
  nand2 I006_073(w_006_073, w_005_046, w_002_029);
  not1 I006_074(w_006_074, w_003_005);
  not1 I006_075(w_006_075, w_005_130);
  not1 I006_076(w_006_076, w_003_029);
  nand2 I006_077(w_006_077, w_004_099, w_003_037);
  not1 I006_078(w_006_078, w_000_604);
  not1 I006_079(w_006_079, w_002_445);
  and2 I006_080(w_006_080, w_001_031, w_001_025);
  and2 I006_081(w_006_081, w_000_270, w_004_072);
  and2 I006_082(w_006_082, w_000_286, w_001_030);
  nand2 I006_083(w_006_083, w_002_266, w_002_322);
  or2  I006_084(w_006_084, w_005_135, w_003_029);
  nand2 I006_085(w_006_085, w_001_001, w_003_023);
  or2  I006_086(w_006_086, w_001_007, w_005_108);
  not1 I006_087(w_006_087, w_003_038);
  and2 I006_088(w_006_088, w_001_023, w_002_090);
  nand2 I006_089(w_006_089, w_004_036, w_003_084);
  or2  I006_090(w_006_090, w_005_149, w_002_168);
  or2  I006_091(w_006_091, w_005_304, w_001_033);
  nand2 I006_092(w_006_092, w_002_577, w_005_093);
  not1 I006_093(w_006_093, w_004_010);
  and2 I006_094(w_006_094, w_001_035, w_002_694);
  or2  I006_095(w_006_095, w_003_019, w_002_079);
  nand2 I006_096(w_006_096, w_005_225, w_004_281);
  or2  I006_097(w_006_097, w_000_159, w_000_058);
  not1 I006_098(w_006_098, w_001_013);
  not1 I006_099(w_006_099, w_004_050);
  nand2 I006_100(w_006_100, w_000_605, w_001_010);
  and2 I006_101(w_006_101, w_000_606, w_004_034);
  nand2 I006_102(w_006_102, w_005_081, w_001_023);
  and2 I006_103(w_006_103, w_001_022, w_002_522);
  not1 I006_104(w_006_104, w_002_681);
  or2  I006_105(w_006_105, w_004_216, w_002_345);
  not1 I006_106(w_006_106, w_004_237);
  or2  I006_107(w_006_107, w_002_615, w_000_031);
  nand2 I006_108(w_006_108, w_004_277, w_001_024);
  and2 I006_109(w_006_109, w_001_013, w_001_024);
  nand2 I006_110(w_006_110, w_000_491, w_003_079);
  or2  I006_111(w_006_111, w_000_607, w_000_146);
  not1 I006_112(w_006_112, w_001_006);
  and2 I006_113(w_006_113, w_003_025, w_001_028);
  or2  I006_114(w_006_114, w_005_314, w_002_291);
  not1 I006_115(w_006_115, w_002_029);
  not1 I006_116(w_006_116, w_001_025);
  or2  I006_117(w_006_117, w_004_272, w_000_473);
  and2 I006_118(w_006_118, w_002_391, w_004_490);
  or2  I006_119(w_006_119, w_000_196, w_002_596);
  and2 I006_120(w_006_120, w_004_076, w_001_004);
  and2 I006_121(w_006_121, w_000_129, w_000_249);
  nand2 I006_122(w_006_122, w_000_543, w_005_007);
  and2 I006_123(w_006_123, w_004_118, w_000_518);
  or2  I006_124(w_006_124, w_000_271, w_004_330);
  or2  I006_125(w_006_125, w_004_083, w_000_334);
  nand2 I006_126(w_006_126, w_000_028, w_005_097);
  and2 I006_127(w_006_127, w_003_034, w_001_001);
  and2 I006_128(w_006_128, w_000_162, w_001_020);
  and2 I006_129(w_006_129, w_005_034, w_000_608);
  not1 I006_130(w_006_130, w_001_005);
  or2  I006_131(w_006_131, w_004_238, w_003_079);
  or2  I006_132(w_006_132, w_001_001, w_004_183);
  nand2 I006_133(w_006_133, w_002_151, w_005_020);
  not1 I006_134(w_006_134, w_001_007);
  not1 I006_135(w_006_135, w_005_036);
  or2  I006_136(w_006_136, w_001_026, w_004_363);
  and2 I006_137(w_006_137, w_003_062, w_001_007);
  nand2 I006_138(w_006_138, w_005_279, w_004_105);
  nand2 I006_139(w_006_139, w_003_036, w_004_122);
  or2  I006_140(w_006_140, w_004_116, w_000_493);
  and2 I006_141(w_006_141, w_001_034, w_004_103);
  nand2 I006_142(w_006_142, w_003_084, w_005_128);
  or2  I006_143(w_006_143, w_005_098, w_004_216);
  not1 I006_144(w_006_144, w_005_042);
  and2 I006_145(w_006_145, w_001_010, w_003_017);
  or2  I006_146(w_006_146, w_001_013, w_004_051);
  nand2 I006_147(w_006_147, w_005_255, w_005_108);
  not1 I006_148(w_006_148, w_003_041);
  or2  I006_149(w_006_149, w_004_005, w_000_609);
  not1 I006_150(w_006_150, w_003_008);
  or2  I006_151(w_006_151, w_003_006, w_002_519);
  nand2 I006_152(w_006_152, w_002_567, w_005_033);
  and2 I006_153(w_006_153, w_000_009, w_001_022);
  and2 I006_154(w_006_154, w_004_495, w_005_087);
  or2  I006_155(w_006_155, w_000_610, w_004_252);
  nand2 I006_156(w_006_156, w_002_127, w_002_101);
  or2  I006_157(w_006_157, w_005_102, w_000_553);
  and2 I006_158(w_006_158, w_002_123, w_005_139);
  and2 I006_159(w_006_159, w_001_006, w_001_034);
  and2 I006_160(w_006_160, w_004_361, w_001_032);
  not1 I006_161(w_006_161, w_005_067);
  not1 I006_162(w_006_162, w_004_449);
  not1 I006_163(w_006_163, w_004_040);
  nand2 I006_164(w_006_164, w_003_066, w_001_009);
  nand2 I006_165(w_006_165, w_001_021, w_002_070);
  not1 I006_166(w_006_166, w_003_008);
  and2 I006_167(w_006_167, w_004_393, w_000_592);
  not1 I006_168(w_006_168, w_003_056);
  nand2 I006_169(w_006_169, w_005_113, w_001_015);
  or2  I006_170(w_006_170, w_004_162, w_001_017);
  or2  I006_171(w_006_171, w_003_005, w_004_042);
  or2  I006_172(w_006_172, w_000_310, w_005_094);
  or2  I006_173(w_006_173, w_000_611, w_003_030);
  and2 I006_174(w_006_174, w_003_078, w_002_334);
  and2 I006_175(w_006_175, w_003_023, w_001_028);
  and2 I006_176(w_006_176, w_002_665, w_002_601);
  and2 I006_177(w_006_177, w_001_011, w_002_475);
  not1 I006_178(w_006_178, w_003_062);
  or2  I006_179(w_006_179, w_002_594, w_004_286);
  and2 I006_180(w_006_180, w_001_027, w_002_618);
  and2 I006_181(w_006_181, w_002_504, w_004_262);
  and2 I006_182(w_006_182, w_005_033, w_004_121);
  or2  I006_183(w_006_183, w_000_433, w_003_010);
  nand2 I006_184(w_006_184, w_003_026, w_004_016);
  and2 I006_185(w_006_185, w_005_093, w_004_049);
  nand2 I006_186(w_006_186, w_001_030, w_002_407);
  not1 I006_187(w_006_187, w_004_028);
  not1 I006_188(w_006_188, w_002_062);
  nand2 I006_189(w_006_189, w_000_414, w_005_095);
  and2 I006_190(w_006_190, w_000_080, w_003_053);
  and2 I006_191(w_006_191, w_001_023, w_004_443);
  or2  I006_192(w_006_192, w_003_056, w_001_001);
  nand2 I006_193(w_006_193, w_000_586, w_005_122);
  and2 I006_194(w_006_194, w_003_042, w_002_421);
  not1 I006_195(w_006_195, w_001_015);
  and2 I006_196(w_006_196, w_001_019, w_002_411);
  or2  I006_197(w_006_197, w_000_186, w_005_099);
  nand2 I006_198(w_006_198, w_003_032, w_004_508);
  not1 I006_199(w_006_199, w_005_246);
  or2  I006_200(w_006_200, w_000_384, w_000_612);
  and2 I006_201(w_006_201, w_003_055, w_003_022);
  not1 I006_202(w_006_202, w_002_236);
  not1 I006_203(w_006_203, w_003_036);
  nand2 I006_204(w_006_204, w_000_439, w_003_002);
  and2 I006_205(w_006_205, w_002_210, w_002_206);
  not1 I006_206(w_006_206, w_004_357);
  or2  I006_207(w_006_207, w_003_026, w_005_140);
  or2  I006_208(w_006_208, w_003_072, w_004_455);
  nand2 I006_209(w_006_209, w_003_008, w_005_103);
  and2 I006_210(w_006_210, w_001_025, w_001_035);
  not1 I006_211(w_006_211, w_004_072);
  nand2 I006_212(w_006_212, w_000_613, w_003_065);
  and2 I006_213(w_006_213, w_005_059, w_004_498);
  not1 I006_214(w_006_214, w_003_000);
  nand2 I006_215(w_006_215, w_001_014, w_001_020);
  or2  I006_216(w_006_216, w_005_119, w_002_133);
  not1 I006_217(w_006_217, w_003_058);
  or2  I006_218(w_006_218, w_001_023, w_003_043);
  not1 I006_219(w_006_219, w_001_012);
  or2  I006_220(w_006_220, w_003_032, w_002_167);
  and2 I006_221(w_006_221, w_003_060, w_000_577);
  and2 I006_222(w_006_222, w_005_272, w_001_031);
  and2 I006_223(w_006_223, w_004_465, w_004_005);
  nand2 I006_224(w_006_224, w_000_586, w_002_217);
  or2  I006_225(w_006_225, w_005_293, w_005_148);
  not1 I006_226(w_006_226, w_002_094);
  or2  I006_227(w_006_227, w_002_613, w_005_248);
  not1 I006_228(w_006_228, w_005_025);
  not1 I006_229(w_006_229, w_002_135);
  nand2 I006_230(w_006_230, w_002_271, w_004_005);
  and2 I006_231(w_006_231, w_005_032, w_000_419);
  nand2 I006_232(w_006_232, w_005_072, w_003_054);
  nand2 I006_233(w_006_233, w_001_004, w_001_030);
  nand2 I006_234(w_006_234, w_004_036, w_002_275);
  and2 I006_235(w_006_235, w_000_172, w_002_010);
  nand2 I006_236(w_006_236, w_000_060, w_005_211);
  and2 I006_237(w_006_237, w_005_044, w_005_210);
  nand2 I006_238(w_006_238, w_002_396, w_005_061);
  nand2 I006_239(w_006_239, w_005_187, w_001_001);
  and2 I006_240(w_006_240, w_002_190, w_001_020);
  not1 I006_241(w_006_241, w_003_020);
  not1 I006_242(w_006_242, w_004_347);
  or2  I006_243(w_006_243, w_004_250, w_004_110);
  and2 I006_244(w_006_244, w_001_025, w_003_001);
  and2 I006_245(w_006_245, w_003_022, w_002_065);
  and2 I006_246(w_006_246, w_001_030, w_003_041);
  and2 I006_247(w_006_247, w_004_124, w_003_010);
  not1 I006_248(w_006_248, w_005_101);
  and2 I006_249(w_006_249, w_003_064, w_003_063);
  nand2 I006_250(w_006_250, w_002_683, w_001_015);
  and2 I006_251(w_006_251, w_002_330, w_003_045);
  not1 I006_252(w_006_252, w_005_046);
  nand2 I006_253(w_006_255, w_003_077, w_006_254);
  and2 I006_254(w_006_256, w_006_255, w_001_031);
  and2 I006_255(w_006_254, w_003_040, w_006_256);
  and2 I007_000(w_007_000, w_004_154, w_000_093);
  not1 I007_001(w_007_001, w_003_079);
  or2  I007_002(w_007_002, w_006_208, w_006_222);
  or2  I007_003(w_007_003, w_006_002, w_006_060);
  nand2 I007_004(w_007_004, w_001_002, w_005_031);
  not1 I007_005(w_007_005, w_003_065);
  not1 I007_006(w_007_006, w_002_183);
  nand2 I007_007(w_007_007, w_006_069, w_002_227);
  or2  I007_008(w_007_008, w_006_081, w_002_286);
  not1 I007_009(w_007_009, w_002_494);
  nand2 I007_010(w_007_010, w_006_194, w_006_019);
  or2  I007_011(w_007_011, w_004_247, w_005_132);
  not1 I007_012(w_007_012, w_006_059);
  and2 I007_013(w_007_013, w_005_083, w_002_230);
  not1 I007_014(w_007_014, w_000_005);
  not1 I007_015(w_007_015, w_004_106);
  and2 I007_016(w_007_016, w_006_052, w_003_074);
  nand2 I007_017(w_007_017, w_003_064, w_000_400);
  and2 I007_018(w_007_018, w_004_064, w_000_600);
  and2 I007_019(w_007_019, w_001_026, w_006_112);
  nand2 I007_020(w_007_020, w_003_023, w_000_541);
  nand2 I007_021(w_007_021, w_005_098, w_002_170);
  or2  I007_022(w_007_022, w_001_014, w_004_154);
  and2 I007_023(w_007_023, w_005_298, w_005_031);
  or2  I007_025(w_007_025, w_001_027, w_002_516);
  or2  I007_026(w_007_026, w_002_027, w_005_315);
  and2 I007_027(w_007_027, w_006_099, w_002_078);
  not1 I007_028(w_007_028, w_005_035);
  not1 I007_029(w_007_029, w_000_614);
  not1 I007_031(w_007_031, w_004_267);
  or2  I007_032(w_007_032, w_005_290, w_001_025);
  or2  I007_033(w_007_033, w_005_038, w_001_007);
  nand2 I007_034(w_007_034, w_002_202, w_004_027);
  or2  I007_035(w_007_035, w_004_040, w_005_147);
  and2 I007_036(w_007_036, w_005_236, w_001_015);
  or2  I007_037(w_007_037, w_002_390, w_002_575);
  nand2 I007_038(w_007_038, w_004_055, w_002_406);
  and2 I007_039(w_007_039, w_001_034, w_006_193);
  or2  I007_040(w_007_040, w_006_121, w_004_456);
  or2  I007_041(w_007_041, w_004_405, w_005_123);
  not1 I007_042(w_007_042, w_003_044);
  nand2 I007_043(w_007_043, w_002_522, w_005_106);
  or2  I007_044(w_007_044, w_000_233, w_001_007);
  or2  I007_045(w_007_045, w_002_557, w_005_047);
  or2  I007_046(w_007_046, w_004_074, w_002_367);
  not1 I007_047(w_007_047, w_006_023);
  nand2 I007_049(w_007_049, w_001_014, w_001_017);
  nand2 I007_050(w_007_050, w_006_200, w_006_221);
  not1 I007_051(w_007_051, w_006_119);
  nand2 I007_052(w_007_052, w_001_019, w_001_003);
  nand2 I007_053(w_007_053, w_004_116, w_001_007);
  not1 I007_054(w_007_054, w_006_032);
  or2  I007_055(w_007_055, w_001_006, w_004_448);
  and2 I007_056(w_007_056, w_003_041, w_004_244);
  or2  I007_057(w_007_057, w_001_000, w_001_006);
  or2  I007_058(w_007_058, w_000_616, w_004_325);
  and2 I007_059(w_007_059, w_005_019, w_005_157);
  or2  I007_060(w_007_060, w_000_617, w_006_031);
  nand2 I007_061(w_007_061, w_004_093, w_006_164);
  nand2 I007_062(w_007_062, w_002_025, w_006_232);
  nand2 I007_063(w_007_063, w_001_017, w_003_043);
  not1 I007_064(w_007_064, w_003_081);
  and2 I007_065(w_007_065, w_005_031, w_001_013);
  or2  I007_066(w_007_066, w_006_065, w_000_549);
  or2  I007_067(w_007_067, w_005_132, w_005_200);
  nand2 I007_068(w_007_068, w_002_488, w_002_207);
  or2  I007_069(w_007_069, w_001_014, w_001_021);
  nand2 I007_070(w_007_070, w_002_277, w_003_033);
  nand2 I007_071(w_007_071, w_003_031, w_004_449);
  and2 I007_072(w_007_072, w_001_025, w_000_374);
  not1 I007_073(w_007_073, w_000_196);
  nand2 I007_074(w_007_074, w_003_012, w_006_001);
  and2 I007_076(w_007_076, w_002_647, w_003_072);
  or2  I007_077(w_007_077, w_000_422, w_002_030);
  or2  I007_078(w_007_078, w_006_032, w_001_021);
  or2  I007_079(w_007_079, w_001_022, w_005_308);
  not1 I007_080(w_007_080, w_002_489);
  not1 I007_081(w_007_081, w_002_031);
  not1 I007_082(w_007_082, w_001_016);
  nand2 I007_083(w_007_083, w_002_312, w_005_073);
  nand2 I007_084(w_007_084, w_003_048, w_000_004);
  or2  I007_085(w_007_085, w_002_605, w_003_032);
  nand2 I007_086(w_007_086, w_000_344, w_000_090);
  nand2 I007_087(w_007_087, w_000_618, w_006_236);
  not1 I007_088(w_007_088, w_001_007);
  and2 I007_089(w_007_089, w_000_619, w_000_097);
  and2 I007_090(w_007_090, w_003_021, w_006_191);
  or2  I007_091(w_007_091, w_000_196, w_003_067);
  or2  I007_092(w_007_092, w_000_354, w_005_211);
  not1 I007_093(w_007_093, w_006_048);
  or2  I007_094(w_007_094, w_004_253, w_005_290);
  or2  I007_096(w_007_096, w_002_349, w_000_620);
  not1 I007_097(w_007_097, w_006_045);
  and2 I007_098(w_007_098, w_006_241, w_002_507);
  nand2 I007_099(w_007_099, w_000_413, w_004_464);
  nand2 I007_100(w_007_100, w_001_025, w_003_039);
  nand2 I007_101(w_007_101, w_001_010, w_001_012);
  or2  I007_102(w_007_102, w_005_204, w_003_016);
  and2 I007_103(w_007_103, w_003_075, w_004_380);
  nand2 I007_104(w_007_104, w_003_020, w_004_117);
  and2 I007_105(w_007_105, w_001_020, w_000_621);
  nand2 I007_106(w_007_106, w_004_231, w_002_358);
  not1 I007_107(w_007_107, w_000_410);
  nand2 I007_108(w_007_108, w_001_011, w_006_010);
  and2 I007_109(w_007_109, w_001_026, w_003_070);
  and2 I007_110(w_007_110, w_005_131, w_000_622);
  nand2 I007_111(w_007_111, w_004_292, w_000_081);
  nand2 I007_112(w_007_112, w_000_064, w_002_313);
  nand2 I007_113(w_007_113, w_002_223, w_004_026);
  not1 I007_114(w_007_114, w_001_020);
  nand2 I007_115(w_007_115, w_000_585, w_006_108);
  and2 I007_116(w_007_116, w_000_531, w_002_385);
  or2  I007_117(w_007_117, w_002_560, w_000_623);
  and2 I007_118(w_007_118, w_005_019, w_001_009);
  nand2 I007_119(w_007_119, w_001_022, w_006_134);
  or2  I007_120(w_007_120, w_003_038, w_000_285);
  not1 I007_121(w_007_121, w_005_108);
  nand2 I007_122(w_007_122, w_002_087, w_000_299);
  not1 I007_123(w_007_123, w_003_066);
  and2 I007_124(w_007_124, w_005_158, w_006_201);
  or2  I007_125(w_007_125, w_005_154, w_001_029);
  nand2 I007_126(w_007_126, w_002_361, w_005_039);
  not1 I007_127(w_007_127, w_006_162);
  or2  I007_128(w_007_128, w_002_412, w_005_104);
  nand2 I007_129(w_007_129, w_000_062, w_001_035);
  or2  I007_130(w_007_130, w_002_530, w_000_463);
  nand2 I007_131(w_007_131, w_006_216, w_002_213);
  not1 I007_132(w_007_132, w_001_020);
  or2  I007_134(w_007_134, w_006_010, w_000_570);
  not1 I007_135(w_007_135, w_005_226);
  or2  I007_136(w_007_136, w_003_012, w_000_475);
  and2 I007_137(w_007_137, w_002_206, w_000_455);
  or2  I007_138(w_007_138, w_000_124, w_001_007);
  not1 I007_139(w_007_139, w_000_186);
  and2 I007_140(w_007_140, w_001_023, w_001_035);
  not1 I007_141(w_007_141, w_005_078);
  or2  I007_142(w_007_142, w_004_371, w_000_624);
  and2 I007_143(w_007_143, w_004_124, w_000_625);
  and2 I007_144(w_007_144, w_002_195, w_000_515);
  and2 I007_145(w_007_145, w_005_192, w_001_009);
  not1 I007_146(w_007_146, w_001_010);
  not1 I007_147(w_007_147, w_002_436);
  not1 I007_148(w_007_148, w_005_040);
  nand2 I007_149(w_007_149, w_006_208, w_005_277);
  or2  I007_150(w_007_150, w_000_622, w_000_615);
  nand2 I007_151(w_007_151, w_004_270, w_001_022);
  not1 I007_152(w_007_152, w_001_032);
  nand2 I007_153(w_007_153, w_003_049, w_003_020);
  or2  I007_154(w_007_154, w_004_332, w_000_626);
  not1 I007_155(w_007_155, w_005_008);
  or2  I007_156(w_007_156, w_003_026, w_006_227);
  or2  I007_157(w_007_157, w_005_107, w_000_179);
  not1 I007_158(w_007_158, w_004_001);
  not1 I007_159(w_007_159, w_005_099);
  or2  I007_160(w_007_160, w_002_576, w_000_627);
  or2  I007_161(w_007_161, w_001_012, w_000_413);
  and2 I007_162(w_007_162, w_006_155, w_003_069);
  or2  I007_163(w_007_163, w_004_037, w_001_002);
  not1 I007_164(w_007_164, w_006_190);
  not1 I007_165(w_007_165, w_005_155);
  not1 I007_166(w_007_166, w_003_052);
  nand2 I007_167(w_007_167, w_002_520, w_004_144);
  and2 I007_168(w_007_168, w_002_327, w_006_022);
  and2 I007_169(w_007_169, w_002_024, w_006_205);
  not1 I007_170(w_007_170, w_000_116);
  and2 I007_171(w_007_171, w_003_035, w_002_046);
  nand2 I007_172(w_007_172, w_004_006, w_006_094);
  not1 I007_173(w_007_173, w_000_628);
  and2 I007_175(w_007_175, w_006_120, w_006_138);
  or2  I007_176(w_007_176, w_002_668, w_000_389);
  not1 I007_177(w_007_177, w_005_057);
  not1 I007_178(w_007_178, w_006_154);
  or2  I007_179(w_007_179, w_005_245, w_006_218);
  or2  I007_180(w_007_180, w_006_230, w_004_139);
  and2 I007_181(w_007_181, w_004_211, w_000_005);
  and2 I007_182(w_007_182, w_005_159, w_000_470);
  nand2 I007_183(w_007_183, w_000_629, w_005_110);
  and2 I007_184(w_007_184, w_003_061, w_001_027);
  or2  I007_185(w_007_185, w_002_698, w_000_075);
  not1 I007_186(w_007_186, w_004_057);
  and2 I007_187(w_007_187, w_001_000, w_006_093);
  not1 I007_188(w_007_188, w_005_033);
  not1 I007_189(w_007_189, w_003_030);
  or2  I007_190(w_007_190, w_003_076, w_006_003);
  nand2 I007_191(w_007_191, w_000_240, w_006_184);
  not1 I007_192(w_007_192, w_006_025);
  or2  I007_193(w_007_193, w_004_269, w_004_287);
  or2  I007_194(w_007_194, w_002_401, w_005_145);
  not1 I007_195(w_007_195, w_006_006);
  and2 I007_196(w_007_196, w_000_372, w_004_191);
  or2  I007_197(w_007_197, w_000_352, w_000_354);
  nand2 I007_198(w_007_198, w_005_275, w_004_149);
  and2 I007_199(w_007_199, w_003_053, w_005_226);
  nand2 I007_200(w_007_200, w_002_303, w_006_037);
  not1 I007_201(w_007_201, w_002_448);
  and2 I007_202(w_007_202, w_003_003, w_000_415);
  or2  I007_203(w_007_203, w_000_161, w_004_341);
  nand2 I007_204(w_007_204, w_000_563, w_000_388);
  nand2 I007_205(w_007_205, w_001_018, w_000_518);
  not1 I007_206(w_007_206, w_005_297);
  or2  I007_207(w_007_207, w_005_281, w_002_351);
  not1 I007_208(w_007_208, w_002_351);
  nand2 I007_209(w_007_209, w_005_161, w_003_067);
  nand2 I007_210(w_007_210, w_003_070, w_002_464);
  nand2 I007_211(w_007_211, w_002_227, w_004_200);
  not1 I007_212(w_007_212, w_003_007);
  nand2 I007_213(w_007_213, w_006_051, w_006_171);
  or2  I007_214(w_007_214, w_002_029, w_003_025);
  nand2 I007_215(w_007_215, w_005_035, w_006_016);
  nand2 I007_216(w_007_216, w_002_141, w_001_033);
  not1 I007_217(w_007_217, w_003_056);
  or2  I007_218(w_007_218, w_006_214, w_000_276);
  nand2 I007_219(w_007_219, w_001_016, w_003_083);
  not1 I007_220(w_007_220, w_001_023);
  and2 I007_221(w_007_221, w_003_001, w_005_065);
  or2  I007_222(w_007_222, w_003_058, w_005_071);
  or2  I007_223(w_007_223, w_006_213, w_000_587);
  nand2 I007_224(w_007_224, w_003_048, w_004_293);
  and2 I007_225(w_007_225, w_004_122, w_005_067);
  and2 I007_226(w_007_226, w_002_361, w_005_148);
  not1 I007_227(w_007_227, w_000_529);
  nand2 I007_228(w_007_228, w_003_028, w_006_067);
  or2  I007_230(w_007_230, w_003_001, w_005_030);
  or2  I007_231(w_007_231, w_002_514, w_006_094);
  and2 I007_232(w_007_232, w_005_285, w_006_165);
  not1 I007_233(w_007_233, w_004_019);
  and2 I007_234(w_007_234, w_002_548, w_003_051);
  not1 I007_235(w_007_235, w_002_542);
  or2  I007_236(w_007_236, w_005_167, w_006_025);
  nand2 I007_237(w_007_237, w_000_279, w_001_036);
  and2 I007_238(w_007_238, w_001_032, w_004_038);
  not1 I007_239(w_007_239, w_002_323);
  not1 I007_240(w_007_240, w_005_170);
  not1 I007_241(w_007_241, w_004_072);
  nand2 I007_244(w_007_244, w_002_097, w_004_425);
  and2 I007_245(w_007_245, w_000_538, w_000_353);
  and2 I007_246(w_007_246, w_005_005, w_005_318);
  or2  I007_247(w_007_247, w_003_007, w_002_098);
  not1 I007_248(w_007_248, w_000_591);
  and2 I007_249(w_007_249, w_001_018, w_000_486);
  and2 I007_250(w_007_250, w_002_292, w_006_191);
  or2  I007_251(w_007_251, w_003_079, w_006_097);
  and2 I007_252(w_007_252, w_006_002, w_004_314);
  or2  I007_253(w_007_253, w_000_504, w_000_036);
  nand2 I007_254(w_007_254, w_002_134, w_006_201);
  not1 I007_255(w_007_255, w_000_020);
  or2  I007_256(w_007_256, w_005_187, w_006_022);
  not1 I007_257(w_007_257, w_003_012);
  nand2 I007_258(w_007_258, w_005_014, w_000_320);
  and2 I007_259(w_007_259, w_000_323, w_003_065);
  and2 I007_260(w_007_260, w_003_036, w_006_071);
  nand2 I007_261(w_007_261, w_002_263, w_001_013);
  or2  I007_262(w_007_262, w_006_244, w_004_024);
  nand2 I007_263(w_007_263, w_001_034, w_001_015);
  not1 I007_264(w_007_264, w_002_423);
  not1 I007_265(w_007_265, w_003_040);
  not1 I007_266(w_007_266, w_001_022);
  nand2 I007_267(w_007_267, w_001_025, w_005_318);
  not1 I007_268(w_007_268, w_001_007);
  and2 I007_269(w_007_269, w_003_008, w_005_186);
  and2 I007_270(w_007_270, w_005_256, w_006_040);
  and2 I007_271(w_007_271, w_002_039, w_005_242);
  or2  I007_272(w_007_272, w_006_176, w_005_231);
  nand2 I007_273(w_007_273, w_004_211, w_005_036);
  and2 I007_274(w_007_274, w_003_014, w_001_008);
  nand2 I007_275(w_007_275, w_004_116, w_004_016);
  not1 I007_276(w_007_276, w_000_554);
  not1 I007_277(w_007_277, w_004_399);
  not1 I007_278(w_007_278, w_006_098);
  not1 I007_279(w_007_279, w_001_030);
  or2  I007_280(w_007_280, w_002_023, w_004_009);
  or2  I007_281(w_007_281, w_000_406, w_001_017);
  and2 I007_282(w_007_282, w_000_427, w_000_107);
  not1 I007_283(w_007_283, w_006_166);
  not1 I007_284(w_007_284, w_006_021);
  and2 I007_285(w_007_285, w_001_023, w_000_191);
  and2 I007_286(w_007_286, w_003_043, w_000_183);
  nand2 I007_287(w_007_287, w_000_558, w_004_328);
  nand2 I007_288(w_007_288, w_004_286, w_002_389);
  not1 I007_289(w_007_289, w_002_016);
  not1 I007_291(w_007_291, w_002_293);
  and2 I007_292(w_007_292, w_005_084, w_006_070);
  not1 I007_293(w_007_293, w_001_010);
  or2  I007_294(w_007_294, w_001_026, w_001_028);
  or2  I007_295(w_007_295, w_004_099, w_000_317);
  nand2 I007_296(w_007_296, w_006_081, w_006_195);
  not1 I007_297(w_007_297, w_001_023);
  not1 I007_299(w_007_299, w_005_204);
  and2 I007_300(w_007_300, w_004_042, w_002_469);
  and2 I007_303(w_007_303, w_005_088, w_006_112);
  nand2 I007_304(w_007_304, w_000_630, w_002_617);
  not1 I007_306(w_007_306, w_001_001);
  and2 I007_307(w_007_307, w_004_188, w_004_228);
  nand2 I007_308(w_007_308, w_003_081, w_002_247);
  nand2 I007_309(w_007_309, w_000_214, w_005_226);
  not1 I007_310(w_007_310, w_002_633);
  or2  I007_312(w_007_312, w_006_019, w_005_271);
  not1 I007_313(w_007_313, w_006_015);
  not1 I007_314(w_007_314, w_001_018);
  not1 I007_315(w_007_315, w_003_008);
  nand2 I007_316(w_007_316, w_006_130, w_005_068);
  not1 I007_318(w_007_318, w_000_043);
  not1 I007_319(w_007_319, w_003_074);
  and2 I007_320(w_007_320, w_006_229, w_001_018);
  or2  I007_321(w_007_321, w_001_022, w_002_597);
  not1 I007_323(w_007_323, w_004_067);
  and2 I007_324(w_007_324, w_000_536, w_003_046);
  not1 I007_325(w_007_325, w_002_352);
  nand2 I007_327(w_007_327, w_003_017, w_004_055);
  and2 I007_328(w_007_328, w_005_268, w_001_002);
  nand2 I007_330(w_007_330, w_005_147, w_004_084);
  not1 I007_331(w_007_331, w_000_632);
  and2 I007_332(w_007_332, w_000_545, w_000_424);
  and2 I007_333(w_007_333, w_004_129, w_000_254);
  and2 I007_334(w_007_334, w_004_019, w_006_036);
  nand2 I007_336(w_007_336, w_000_590, w_004_174);
  and2 I007_337(w_007_337, w_001_034, w_002_288);
  or2  I007_339(w_007_339, w_006_030, w_003_031);
  nand2 I007_340(w_007_340, w_001_016, w_001_009);
  not1 I007_342(w_007_342, w_003_030);
  and2 I007_343(w_007_343, w_005_169, w_006_014);
  or2  I007_345(w_007_345, w_002_181, w_005_299);
  not1 I007_346(w_007_346, w_001_025);
  or2  I007_347(w_007_347, w_002_263, w_005_304);
  nand2 I007_348(w_007_348, w_003_006, w_000_365);
  not1 I007_349(w_007_349, w_001_018);
  not1 I007_350(w_007_350, w_006_218);
  nand2 I007_351(w_007_351, w_005_124, w_000_061);
  and2 I007_353(w_007_353, w_000_634, w_005_295);
  nand2 I007_354(w_007_354, w_005_110, w_002_230);
  and2 I007_356(w_007_356, w_005_292, w_000_218);
  not1 I007_357(w_007_357, w_006_242);
  nand2 I007_359(w_007_359, w_004_497, w_002_304);
  or2  I007_360(w_007_360, w_001_007, w_002_438);
  or2  I007_361(w_007_361, w_000_549, w_003_058);
  nand2 I007_362(w_007_362, w_006_020, w_006_175);
  not1 I007_363(w_007_363, w_006_199);
  and2 I007_364(w_007_364, w_003_076, w_003_054);
  or2  I007_365(w_007_365, w_006_056, w_004_124);
  nand2 I007_367(w_007_367, w_006_250, w_001_016);
  or2  I007_368(w_007_368, w_006_215, w_002_600);
  nand2 I007_371(w_007_371, w_004_191, w_002_216);
  and2 I007_372(w_007_372, w_000_051, w_005_051);
  or2  I007_373(w_007_373, w_004_174, w_000_309);
  nand2 I007_374(w_007_374, w_006_244, w_005_024);
  or2  I007_377(w_007_377, w_006_216, w_001_010);
  not1 I007_378(w_007_378, w_003_016);
  or2  I007_379(w_007_379, w_001_011, w_006_144);
  and2 I007_380(w_007_380, w_006_200, w_003_023);
  nand2 I007_381(w_007_381, w_001_012, w_003_032);
  not1 I007_382(w_007_382, w_000_313);
  or2  I007_384(w_007_384, w_005_201, w_003_058);
  not1 I007_385(w_007_385, w_006_248);
  and2 I007_386(w_007_386, w_005_127, w_001_018);
  not1 I007_387(w_007_387, w_000_254);
  or2  I007_389(w_007_389, w_005_089, w_000_299);
  nand2 I007_390(w_007_390, w_004_444, w_002_658);
  not1 I007_391(w_007_391, w_004_289);
  and2 I007_392(w_007_392, w_002_673, w_000_385);
  and2 I007_393(w_007_393, w_004_179, w_000_482);
  and2 I007_394(w_007_394, w_002_409, w_005_180);
  nand2 I007_395(w_007_395, w_000_489, w_004_090);
  not1 I007_396(w_007_396, w_003_049);
  or2  I007_397(w_007_397, w_005_066, w_003_041);
  and2 I007_398(w_007_398, w_005_188, w_003_024);
  nand2 I007_400(w_007_400, w_004_032, w_000_603);
  and2 I007_403(w_007_403, w_003_064, w_006_052);
  nand2 I007_405(w_007_405, w_004_079, w_001_010);
  and2 I007_407(w_007_407, w_004_055, w_001_017);
  and2 I007_408(w_007_408, w_004_302, w_006_147);
  and2 I007_410(w_007_410, w_004_212, w_006_120);
  nand2 I007_413(w_007_413, w_006_075, w_004_309);
  nand2 I007_414(w_007_414, w_005_152, w_006_094);
  or2  I007_415(w_007_415, w_003_068, w_004_359);
  not1 I007_416(w_007_416, w_002_300);
  not1 I007_418(w_007_418, w_005_295);
  not1 I007_419(w_007_419, w_002_021);
  not1 I007_420(w_007_420, w_004_033);
  nand2 I007_421(w_007_421, w_003_071, w_004_235);
  not1 I007_422(w_007_422, w_005_213);
  or2  I007_423(w_007_423, w_002_308, w_006_196);
  and2 I007_424(w_007_424, w_002_261, w_002_247);
  or2  I007_425(w_007_425, w_000_403, w_001_025);
  nand2 I007_426(w_007_426, w_000_097, w_006_182);
  nand2 I007_427(w_007_427, w_002_468, w_002_465);
  or2  I007_428(w_007_428, w_006_003, w_005_144);
  nand2 I007_429(w_007_429, w_003_037, w_002_684);
  not1 I007_431(w_007_431, w_002_190);
  or2  I007_432(w_007_432, w_002_289, w_001_036);
  or2  I007_434(w_007_434, w_001_007, w_003_017);
  or2  I007_436(w_007_436, w_002_344, w_006_026);
  and2 I007_437(w_007_437, w_004_054, w_006_013);
  and2 I007_438(w_007_438, w_006_203, w_006_045);
  or2  I007_439(w_007_439, w_005_307, w_005_232);
  not1 I007_440(w_007_440, w_000_039);
  not1 I007_441(w_007_441, w_001_034);
  nand2 I007_443(w_007_443, w_004_115, w_000_055);
  and2 I007_444(w_007_444, w_002_461, w_003_056);
  or2  I007_445(w_007_445, w_000_637, w_003_009);
  or2  I007_447(w_007_447, w_006_035, w_003_019);
  nand2 I007_448(w_007_448, w_000_589, w_006_184);
  or2  I007_449(w_007_449, w_000_312, w_004_431);
  nand2 I007_450(w_007_450, w_006_139, w_006_011);
  not1 I007_451(w_007_451, w_003_009);
  or2  I007_452(w_007_452, w_006_192, w_005_086);
  or2  I007_453(w_007_453, w_006_181, w_006_045);
  not1 I007_454(w_007_454, w_000_549);
  or2  I007_455(w_007_455, w_000_639, w_005_026);
  and2 I007_456(w_007_456, w_004_147, w_005_053);
  not1 I007_459(w_007_459, w_002_043);
  and2 I007_460(w_007_460, w_006_029, w_003_033);
  nand2 I007_461(w_007_461, w_003_050, w_000_575);
  not1 I007_462(w_007_462, w_004_472);
  not1 I007_463(w_007_463, w_001_016);
  not1 I007_464(w_007_464, w_003_010);
  or2  I007_469(w_007_469, w_006_223, w_003_048);
  nand2 I007_470(w_007_470, w_004_282, w_001_004);
  not1 I007_471(w_007_471, w_003_033);
  or2  I007_472(w_007_472, w_002_377, w_005_077);
  and2 I007_473(w_007_473, w_003_076, w_003_051);
  and2 I007_474(w_007_474, w_004_124, w_004_319);
  or2  I007_475(w_007_475, w_001_034, w_002_021);
  nand2 I007_477(w_007_477, w_001_002, w_006_073);
  or2  I007_478(w_007_478, w_003_003, w_001_033);
  nand2 I007_480(w_007_480, w_003_042, w_004_146);
  and2 I007_482(w_006_258, w_000_657, w_006_254);
  or2  I008_001(w_008_001, w_006_096, w_002_081);
  and2 I008_003(w_008_003, w_007_008, w_006_091);
  or2  I008_004(w_008_004, w_007_361, w_005_267);
  and2 I008_005(w_008_005, w_006_220, w_001_006);
  and2 I008_008(w_008_008, w_002_414, w_005_088);
  and2 I008_009(w_008_009, w_001_035, w_003_061);
  and2 I008_010(w_008_010, w_004_161, w_005_042);
  or2  I008_011(w_008_011, w_001_032, w_005_123);
  or2  I008_012(w_008_012, w_000_533, w_002_013);
  or2  I008_013(w_008_013, w_002_103, w_004_420);
  nand2 I008_014(w_008_014, w_000_414, w_001_015);
  not1 I008_015(w_008_015, w_002_198);
  or2  I008_016(w_008_016, w_005_111, w_001_008);
  or2  I008_017(w_008_017, w_006_150, w_006_095);
  not1 I008_018(w_008_018, w_003_004);
  and2 I008_019(w_008_019, w_003_028, w_006_123);
  and2 I008_020(w_008_020, w_000_031, w_004_150);
  not1 I008_021(w_008_021, w_004_117);
  and2 I008_022(w_008_022, w_001_016, w_006_190);
  not1 I008_023(w_008_023, w_003_083);
  nand2 I008_024(w_008_024, w_004_021, w_005_064);
  or2  I008_025(w_008_025, w_004_482, w_004_215);
  not1 I008_026(w_008_026, w_007_100);
  and2 I008_027(w_008_027, w_007_141, w_004_288);
  or2  I008_028(w_008_028, w_000_056, w_006_222);
  and2 I008_029(w_008_029, w_007_228, w_002_503);
  not1 I008_030(w_008_030, w_005_062);
  or2  I008_031(w_008_031, w_002_112, w_006_188);
  or2  I008_032(w_008_032, w_002_123, w_005_312);
  or2  I008_033(w_008_033, w_004_254, w_005_228);
  or2  I008_034(w_008_034, w_001_023, w_003_054);
  not1 I008_035(w_008_035, w_001_014);
  not1 I008_036(w_008_036, w_000_640);
  or2  I008_037(w_008_037, w_000_180, w_006_152);
  not1 I008_038(w_008_038, w_000_518);
  and2 I008_039(w_008_039, w_002_575, w_007_397);
  or2  I008_040(w_008_040, w_007_021, w_001_033);
  and2 I008_041(w_008_041, w_005_038, w_006_140);
  and2 I008_042(w_008_042, w_000_352, w_001_025);
  nand2 I008_043(w_008_043, w_001_023, w_000_641);
  and2 I008_044(w_008_044, w_006_173, w_002_271);
  or2  I008_045(w_008_045, w_006_039, w_004_349);
  not1 I008_046(w_008_046, w_001_025);
  or2  I008_047(w_008_047, w_003_026, w_002_592);
  or2  I008_048(w_008_048, w_000_642, w_005_256);
  nand2 I008_049(w_008_049, w_006_219, w_006_231);
  or2  I008_050(w_008_050, w_006_252, w_001_013);
  and2 I008_051(w_008_051, w_003_029, w_005_146);
  and2 I008_052(w_008_052, w_001_034, w_003_026);
  nand2 I008_053(w_008_053, w_000_046, w_003_039);
  not1 I008_054(w_008_054, w_000_394);
  and2 I008_055(w_008_055, w_005_202, w_003_057);
  and2 I008_056(w_008_056, w_001_015, w_005_192);
  or2  I008_059(w_008_059, w_007_045, w_005_063);
  and2 I008_061(w_008_061, w_006_065, w_007_185);
  not1 I008_062(w_008_062, w_007_289);
  or2  I008_063(w_008_063, w_004_034, w_001_001);
  not1 I008_064(w_008_064, w_005_028);
  or2  I008_067(w_008_067, w_006_074, w_000_345);
  and2 I008_068(w_008_068, w_002_179, w_005_135);
  or2  I008_069(w_008_069, w_004_024, w_002_118);
  and2 I008_071(w_008_071, w_003_070, w_001_013);
  and2 I008_072(w_008_072, w_007_297, w_006_040);
  not1 I008_073(w_008_073, w_007_219);
  not1 I008_074(w_008_074, w_000_599);
  nand2 I008_076(w_008_076, w_004_207, w_005_154);
  and2 I008_077(w_008_077, w_003_041, w_005_068);
  or2  I008_078(w_008_078, w_000_337, w_002_590);
  not1 I008_079(w_008_079, w_001_015);
  nand2 I008_082(w_008_082, w_006_056, w_002_027);
  nand2 I008_083(w_008_083, w_000_445, w_004_253);
  nand2 I008_084(w_008_084, w_001_017, w_004_066);
  nand2 I008_085(w_008_085, w_007_208, w_005_017);
  or2  I008_088(w_008_088, w_000_544, w_005_270);
  and2 I008_089(w_008_089, w_007_079, w_000_527);
  nand2 I008_090(w_008_090, w_004_490, w_002_013);
  nand2 I008_093(w_008_093, w_001_025, w_007_227);
  nand2 I008_094(w_008_094, w_005_276, w_000_490);
  not1 I008_095(w_008_095, w_000_257);
  nand2 I008_096(w_008_096, w_000_337, w_002_452);
  nand2 I008_097(w_008_097, w_004_220, w_004_069);
  not1 I008_099(w_008_099, w_004_147);
  not1 I008_100(w_008_100, w_005_030);
  not1 I008_103(w_008_103, w_006_125);
  or2  I008_105(w_008_105, w_005_127, w_004_447);
  and2 I008_107(w_008_107, w_003_048, w_005_177);
  not1 I008_108(w_008_108, w_003_070);
  or2  I008_110(w_008_110, w_006_092, w_003_040);
  or2  I008_111(w_008_111, w_002_708, w_000_293);
  or2  I008_112(w_008_112, w_006_233, w_001_031);
  not1 I008_114(w_008_114, w_001_029);
  nand2 I008_115(w_008_115, w_002_212, w_002_056);
  nand2 I008_117(w_008_117, w_004_113, w_002_212);
  not1 I008_118(w_008_118, w_005_154);
  or2  I008_121(w_008_121, w_007_377, w_004_123);
  or2  I008_122(w_008_122, w_007_153, w_004_091);
  and2 I008_124(w_008_124, w_004_484, w_006_159);
  or2  I008_125(w_008_125, w_005_068, w_003_046);
  or2  I008_126(w_008_126, w_003_062, w_004_009);
  and2 I008_127(w_008_127, w_002_624, w_005_046);
  or2  I008_128(w_008_128, w_003_042, w_003_022);
  and2 I008_129(w_008_129, w_006_194, w_007_424);
  not1 I008_130(w_008_130, w_007_060);
  not1 I008_131(w_008_131, w_005_088);
  not1 I008_133(w_008_133, w_002_290);
  nand2 I008_134(w_008_134, w_003_046, w_001_005);
  nand2 I008_135(w_008_135, w_007_477, w_006_147);
  and2 I008_136(w_008_136, w_006_133, w_006_038);
  and2 I008_137(w_008_137, w_006_210, w_003_020);
  and2 I008_138(w_008_138, w_001_035, w_003_058);
  or2  I008_140(w_008_140, w_004_077, w_004_431);
  or2  I008_142(w_008_142, w_003_071, w_001_017);
  nand2 I008_143(w_008_143, w_000_354, w_003_009);
  not1 I008_145(w_008_145, w_000_644);
  or2  I008_147(w_008_147, w_006_073, w_002_379);
  or2  I008_149(w_008_149, w_004_284, w_000_284);
  not1 I008_150(w_008_150, w_003_015);
  not1 I008_152(w_008_152, w_000_126);
  nand2 I008_153(w_008_153, w_003_069, w_005_073);
  nand2 I008_156(w_008_156, w_007_086, w_007_395);
  or2  I008_157(w_008_157, w_002_206, w_000_646);
  and2 I008_159(w_008_159, w_000_238, w_004_275);
  nand2 I008_161(w_008_161, w_005_014, w_006_246);
  or2  I008_162(w_008_162, w_005_011, w_001_016);
  nand2 I008_164(w_008_164, w_002_082, w_003_028);
  and2 I008_167(w_008_167, w_005_143, w_000_647);
  not1 I008_168(w_008_168, w_006_071);
  and2 I008_169(w_008_169, w_007_201, w_004_151);
  nand2 I008_170(w_008_170, w_004_027, w_002_086);
  or2  I008_171(w_008_171, w_005_302, w_001_002);
  nand2 I008_172(w_008_172, w_006_059, w_000_648);
  not1 I008_173(w_008_173, w_006_176);
  nand2 I008_175(w_008_175, w_000_066, w_005_306);
  not1 I008_178(w_008_178, w_007_443);
  and2 I008_179(w_008_179, w_004_210, w_001_024);
  and2 I008_180(w_008_180, w_005_292, w_004_341);
  not1 I008_181(w_008_181, w_006_209);
  nand2 I008_182(w_008_182, w_005_136, w_002_076);
  nand2 I008_183(w_008_183, w_004_161, w_001_008);
  or2  I008_184(w_008_184, w_003_056, w_000_197);
  or2  I008_186(w_008_186, w_001_025, w_001_013);
  and2 I008_188(w_008_188, w_004_007, w_003_051);
  not1 I008_189(w_008_189, w_006_101);
  not1 I008_190(w_008_190, w_002_262);
  nand2 I008_191(w_008_191, w_005_148, w_002_450);
  nand2 I008_192(w_008_192, w_007_469, w_003_027);
  or2  I008_193(w_008_193, w_007_105, w_007_191);
  not1 I008_194(w_008_194, w_005_089);
  nand2 I008_196(w_008_196, w_005_270, w_001_030);
  nand2 I008_198(w_008_198, w_006_101, w_006_080);
  and2 I008_199(w_008_199, w_001_029, w_005_154);
  not1 I008_200(w_008_200, w_004_217);
  and2 I008_202(w_008_202, w_005_244, w_003_021);
  not1 I008_205(w_008_205, w_005_125);
  not1 I008_206(w_008_206, w_007_450);
  and2 I008_207(w_008_207, w_007_303, w_004_041);
  not1 I008_208(w_008_208, w_006_185);
  nand2 I008_209(w_008_209, w_001_024, w_000_636);
  and2 I008_210(w_008_210, w_002_222, w_000_326);
  and2 I008_211(w_008_211, w_000_650, w_005_168);
  or2  I008_212(w_008_212, w_005_106, w_006_160);
  or2  I008_213(w_008_213, w_005_030, w_005_310);
  or2  I008_214(w_008_214, w_001_000, w_007_056);
  nand2 I008_215(w_008_215, w_002_129, w_001_027);
  not1 I008_216(w_008_216, w_005_124);
  and2 I008_217(w_008_217, w_006_002, w_000_182);
  and2 I008_218(w_008_218, w_005_031, w_005_059);
  or2  I008_220(w_008_220, w_002_182, w_006_151);
  and2 I008_221(w_008_221, w_006_207, w_004_194);
  or2  I008_222(w_008_222, w_005_316, w_003_079);
  nand2 I008_223(w_008_223, w_007_272, w_002_631);
  and2 I008_225(w_008_225, w_004_047, w_005_113);
  and2 I008_226(w_008_226, w_002_337, w_005_046);
  and2 I008_227(w_008_227, w_003_004, w_004_145);
  or2  I008_228(w_008_228, w_000_050, w_002_677);
  and2 I008_230(w_008_230, w_006_008, w_007_325);
  or2  I008_232(w_008_232, w_000_651, w_005_044);
  and2 I008_236(w_008_236, w_005_135, w_006_213);
  nand2 I008_237(w_008_237, w_004_141, w_001_029);
  and2 I008_239(w_008_239, w_000_400, w_002_035);
  nand2 I008_240(w_008_240, w_004_227, w_005_003);
  and2 I008_241(w_008_241, w_004_042, w_002_044);
  not1 I008_243(w_008_243, w_005_061);
  nand2 I008_244(w_008_244, w_006_028, w_000_077);
  or2  I008_246(w_008_246, w_000_300, w_000_636);
  nand2 I008_247(w_008_247, w_005_192, w_004_076);
  or2  I008_248(w_008_248, w_006_036, w_004_433);
  nand2 I008_249(w_008_249, w_006_030, w_005_107);
  and2 I008_250(w_008_250, w_000_652, w_007_230);
  or2  I008_252(w_008_252, w_000_334, w_005_256);
  and2 I008_254(w_008_254, w_003_033, w_006_159);
  and2 I008_255(w_008_255, w_005_246, w_003_018);
  nand2 I008_257(w_008_257, w_002_011, w_003_079);
  not1 I008_258(w_008_258, w_004_222);
  or2  I008_261(w_008_261, w_003_024, w_006_246);
  not1 I008_262(w_008_262, w_001_021);
  nand2 I008_264(w_008_264, w_005_180, w_003_043);
  not1 I008_266(w_008_266, w_001_011);
  nand2 I008_268(w_008_268, w_005_275, w_000_155);
  not1 I008_269(w_008_269, w_000_257);
  and2 I008_271(w_008_271, w_005_200, w_004_122);
  and2 I008_272(w_008_272, w_004_222, w_004_039);
  or2  I008_273(w_008_273, w_002_494, w_003_048);
  nand2 I008_274(w_008_274, w_004_179, w_006_197);
  not1 I008_275(w_008_275, w_004_277);
  not1 I008_277(w_008_277, w_000_653);
  and2 I008_278(w_008_278, w_002_249, w_006_005);
  or2  I008_281(w_008_281, w_006_157, w_007_103);
  nand2 I008_282(w_008_282, w_007_028, w_006_240);
  and2 I008_283(w_008_283, w_000_313, w_006_099);
  and2 I008_284(w_008_284, w_001_024, w_000_363);
  not1 I008_285(w_008_285, w_003_079);
  and2 I008_287(w_008_287, w_007_110, w_005_069);
  not1 I008_288(w_008_288, w_005_016);
  or2  I008_289(w_008_289, w_004_206, w_003_029);
  or2  I008_290(w_008_290, w_003_065, w_003_018);
  nand2 I008_291(w_008_291, w_004_212, w_004_119);
  not1 I008_292(w_008_292, w_007_154);
  and2 I008_295(w_008_295, w_004_239, w_005_283);
  or2  I008_298(w_008_298, w_004_207, w_005_156);
  nand2 I008_299(w_008_299, w_004_311, w_005_154);
  not1 I008_300(w_008_300, w_005_047);
  or2  I008_301(w_008_301, w_005_084, w_001_002);
  not1 I008_302(w_008_302, w_007_396);
  or2  I008_304(w_008_304, w_003_073, w_007_473);
  or2  I008_307(w_008_307, w_006_067, w_007_018);
  nand2 I008_309(w_008_309, w_005_297, w_006_101);
  nand2 I008_310(w_008_310, w_007_054, w_004_068);
  not1 I008_312(w_008_312, w_004_199);
  not1 I008_314(w_008_314, w_006_167);
  or2  I008_315(w_008_315, w_007_072, w_006_078);
  not1 I008_316(w_008_316, w_004_370);
  or2  I008_317(w_008_317, w_003_073, w_006_213);
  not1 I008_318(w_008_318, w_005_065);
  and2 I008_319(w_008_319, w_001_014, w_006_035);
  nand2 I008_320(w_008_320, w_005_043, w_006_223);
  and2 I008_322(w_008_322, w_002_282, w_000_589);
  nand2 I008_325(w_008_325, w_005_147, w_003_073);
  not1 I008_327(w_008_327, w_006_132);
  nand2 I008_329(w_008_329, w_005_306, w_007_330);
  nand2 I008_331(w_008_331, w_007_004, w_007_192);
  not1 I008_332(w_008_332, w_001_012);
  nand2 I008_333(w_008_333, w_004_184, w_001_028);
  nand2 I008_334(w_008_334, w_005_121, w_006_201);
  or2  I008_335(w_008_335, w_004_184, w_007_113);
  and2 I008_336(w_008_336, w_004_453, w_007_084);
  and2 I008_337(w_008_337, w_005_044, w_007_324);
  not1 I008_338(w_008_338, w_006_010);
  and2 I008_339(w_008_339, w_007_157, w_003_050);
  not1 I008_341(w_008_341, w_003_017);
  nand2 I008_342(w_008_342, w_007_372, w_002_570);
  and2 I008_343(w_008_343, w_007_224, w_003_009);
  and2 I008_344(w_008_344, w_001_023, w_007_381);
  and2 I008_345(w_008_345, w_005_098, w_004_188);
  or2  I008_346(w_008_346, w_000_654, w_007_099);
  and2 I008_347(w_008_347, w_004_057, w_002_103);
  not1 I008_348(w_008_348, w_005_207);
  not1 I008_349(w_008_349, w_000_296);
  not1 I008_350(w_008_350, w_007_072);
  not1 I008_351(w_008_351, w_004_274);
  nand2 I008_352(w_008_352, w_006_135, w_004_506);
  and2 I008_353(w_008_353, w_006_174, w_000_216);
  not1 I008_354(w_008_354, w_007_143);
  nand2 I008_355(w_008_355, w_004_299, w_002_646);
  not1 I008_356(w_008_356, w_005_062);
  and2 I008_357(w_008_357, w_003_057, w_000_438);
  nand2 I008_358(w_008_358, w_001_036, w_007_385);
  or2  I008_360(w_008_360, w_006_033, w_006_145);
  and2 I008_361(w_008_361, w_005_093, w_000_625);
  and2 I008_362(w_008_362, w_002_472, w_002_295);
  or2  I008_364(w_008_364, w_003_052, w_005_090);
  nand2 I008_366(w_008_366, w_003_046, w_005_202);
  nand2 I008_367(w_008_367, w_002_703, w_000_626);
  nand2 I008_370(w_008_370, w_000_655, w_002_501);
  not1 I008_371(w_008_371, w_007_269);
  or2  I008_374(w_008_374, w_001_010, w_006_193);
  not1 I008_376(w_008_376, w_001_007);
  nand2 I008_377(w_008_377, w_005_027, w_003_004);
  not1 I008_378(w_008_378, w_003_056);
  nand2 I008_381(w_008_381, w_007_200, w_000_497);
  not1 I008_382(w_008_382, w_003_025);
  or2  I008_383(w_008_383, w_003_020, w_006_086);
  and2 I008_384(w_008_384, w_003_008, w_000_376);
  or2  I008_386(w_008_386, w_007_351, w_001_008);
  nand2 I008_387(w_008_387, w_006_211, w_007_086);
  and2 I008_388(w_008_388, w_007_101, w_002_099);
  not1 I008_389(w_008_389, w_007_238);
  nand2 I008_390(w_008_390, w_005_038, w_004_067);
  or2  I008_391(w_008_391, w_004_153, w_001_008);
  or2  I008_394(w_008_394, w_005_303, w_004_037);
  and2 I008_396(w_008_396, w_005_118, w_004_075);
  or2  I008_397(w_008_397, w_000_652, w_007_188);
  or2  I008_398(w_008_398, w_000_155, w_005_236);
  not1 I008_399(w_008_399, w_002_175);
  or2  I008_402(w_008_402, w_004_039, w_001_017);
  not1 I008_403(w_008_403, w_005_254);
  nand2 I008_404(w_008_404, w_005_139, w_002_321);
  not1 I008_405(w_008_405, w_002_028);
  not1 I008_407(w_008_407, w_007_289);
  and2 I008_408(w_008_408, w_006_159, w_006_158);
  nand2 I008_409(w_008_409, w_004_021, w_007_113);
  not1 I008_411(w_008_411, w_002_215);
  and2 I008_413(w_008_413, w_002_406, w_006_216);
  or2  I008_414(w_008_414, w_005_057, w_001_006);
  or2  I008_416(w_008_416, w_003_044, w_000_348);
  and2 I008_417(w_008_417, w_002_551, w_004_088);
  or2  I008_418(w_008_418, w_006_150, w_006_178);
  or2  I008_419(w_008_419, w_002_554, w_006_132);
  and2 I008_420(w_008_420, w_004_190, w_005_185);
  or2  I008_421(w_008_421, w_006_076, w_003_003);
  and2 I008_423(w_008_423, w_000_391, w_003_019);
  nand2 I008_424(w_008_424, w_001_019, w_007_359);
  or2  I008_425(w_008_425, w_005_011, w_007_313);
  or2  I008_426(w_008_426, w_000_231, w_001_013);
  or2  I008_428(w_008_428, w_003_079, w_002_444);
  and2 I008_429(w_008_429, w_006_124, w_003_018);
  not1 I008_431(w_008_431, w_002_231);
  and2 I008_432(w_008_432, w_002_578, w_001_014);
  or2  I008_433(w_008_433, w_003_002, w_001_022);
  nand2 I008_434(w_008_434, w_005_036, w_005_056);
  nand2 I008_435(w_008_435, w_007_018, w_007_155);
  or2  I008_436(w_008_436, w_002_655, w_002_645);
  not1 I008_437(w_008_437, w_007_197);
  and2 I008_439(w_008_439, w_002_510, w_001_019);
  and2 I008_441(w_008_441, w_006_213, w_007_291);
  and2 I008_442(w_008_442, w_007_128, w_005_018);
  and2 I008_444(w_008_444, w_007_413, w_001_012);
  nand2 I008_446(w_008_446, w_004_084, w_000_054);
  or2  I008_449(w_008_449, w_004_099, w_004_039);
  or2  I008_453(w_008_453, w_006_075, w_005_075);
  not1 I008_454(w_008_454, w_004_197);
  nand2 I008_457(w_008_457, w_002_053, w_001_015);
  and2 I008_459(w_008_459, w_005_023, w_001_033);
  not1 I008_460(w_008_460, w_000_333);
  nand2 I008_461(w_008_461, w_001_007, w_007_148);
  or2  I008_463(w_008_463, w_007_363, w_005_095);
  nand2 I008_466(w_008_466, w_004_094, w_004_113);
  or2  I008_467(w_008_467, w_003_025, w_005_304);
  nand2 I008_468(w_008_468, w_006_206, w_002_378);
  not1 I008_469(w_008_469, w_003_057);
  or2  I008_471(w_008_471, w_004_078, w_001_028);
  not1 I008_472(w_008_472, w_006_190);
  or2  I008_473(w_008_473, w_002_599, w_001_027);
  and2 I008_474(w_008_474, w_004_237, w_002_349);
  not1 I008_475(w_008_475, w_000_360);
  not1 I008_477(w_008_477, w_007_309);
  not1 I008_478(w_008_478, w_001_022);
  not1 I008_479(w_008_479, w_000_656);
  or2  I008_480(w_008_480, w_006_108, w_000_083);
  and2 I008_482(w_008_482, w_000_657, w_005_310);
  not1 I008_483(w_008_483, w_006_178);
  or2  I008_484(w_008_484, w_004_070, w_004_186);
  nand2 I008_485(w_008_485, w_001_004, w_005_184);
  nand2 I008_486(w_008_486, w_005_152, w_001_035);
  not1 I008_487(w_008_487, w_001_003);
  nand2 I008_488(w_008_488, w_001_026, w_003_014);
  not1 I008_489(w_008_489, w_003_001);
  and2 I008_490(w_008_490, w_002_105, w_006_215);
  or2  I008_493(w_008_493, w_003_035, w_006_108);
  and2 I008_494(w_008_494, w_000_428, w_007_239);
  not1 I008_495(w_008_495, w_002_542);
  and2 I008_496(w_008_496, w_006_207, w_000_120);
  or2  I008_498(w_008_498, w_001_003, w_004_184);
  and2 I008_499(w_008_499, w_005_288, w_006_193);
  nand2 I008_501(w_008_501, w_004_109, w_006_027);
  or2  I008_502(w_008_502, w_001_016, w_001_028);
  and2 I008_504(w_008_504, w_004_369, w_007_102);
  nand2 I008_505(w_008_505, w_007_189, w_007_203);
  nand2 I008_506(w_008_506, w_005_262, w_003_057);
  or2  I008_509(w_008_509, w_003_048, w_001_025);
  and2 I008_510(w_008_510, w_007_019, w_000_659);
  nand2 I008_511(w_008_511, w_000_484, w_006_015);
  or2  I008_514(w_008_514, w_001_026, w_003_048);
  or2  I008_515(w_008_515, w_000_446, w_006_052);
  nand2 I008_516(w_008_516, w_006_168, w_000_279);
  and2 I008_517(w_008_517, w_007_447, w_000_574);
  not1 I008_518(w_008_518, w_001_005);
  nand2 I008_519(w_008_519, w_006_239, w_007_382);
  nand2 I008_520(w_008_520, w_006_258, w_004_145);
  and2 I008_521(w_008_521, w_007_340, w_002_367);
  not1 I008_522(w_008_522, w_000_224);
  or2  I008_523(w_008_523, w_007_392, w_006_182);
  and2 I008_524(w_008_524, w_005_310, w_004_283);
  nand2 I008_525(w_008_525, w_006_245, w_007_162);
  not1 I008_526(w_008_526, w_006_227);
  and2 I008_528(w_008_528, w_004_222, w_002_491);
  and2 I008_530(w_008_530, w_002_660, w_002_608);
  or2  I008_533(w_008_533, w_005_218, w_002_635);
  not1 I008_534(w_008_534, w_000_227);
  nand2 I008_535(w_008_535, w_004_159, w_001_023);
  nand2 I008_538(w_008_538, w_005_096, w_004_152);
  and2 I008_539(w_008_539, w_003_058, w_001_002);
  and2 I008_541(w_008_541, w_004_471, w_007_240);
  and2 I008_543(w_008_543, w_005_124, w_005_156);
  nand2 I008_544(w_008_544, w_001_028, w_003_046);
  not1 I008_545(w_008_545, w_000_490);
  and2 I008_548(w_008_548, w_003_033, w_004_244);
  nand2 I008_550(w_008_550, w_005_111, w_000_449);
  nand2 I008_552(w_008_552, w_007_198, w_007_083);
  and2 I008_553(w_008_553, w_001_031, w_001_003);
  and2 I008_555(w_008_555, w_006_011, w_004_210);
  nand2 I008_556(w_008_556, w_000_057, w_002_045);
  not1 I008_557(w_008_557, w_003_069);
  or2  I008_558(w_008_558, w_007_155, w_004_230);
  nand2 I008_559(w_008_559, w_004_285, w_003_045);
  not1 I008_560(w_008_560, w_004_081);
  nand2 I008_561(w_008_561, w_005_089, w_002_560);
  or2  I008_562(w_008_562, w_000_278, w_005_154);
  or2  I008_563(w_008_563, w_006_149, w_000_419);
  or2  I008_565(w_008_565, w_006_001, w_000_610);
  and2 I008_566(w_008_566, w_003_060, w_007_040);
  or2  I008_567(w_008_567, w_006_093, w_002_344);
  not1 I008_568(w_008_568, w_004_416);
  and2 I008_569(w_008_569, w_001_020, w_001_026);
  nand2 I008_571(w_008_571, w_004_445, w_004_137);
  not1 I008_572(w_008_572, w_002_648);
  not1 I008_573(w_008_573, w_004_038);
  or2  I008_574(w_008_574, w_004_267, w_005_205);
  or2  I008_575(w_008_575, w_003_050, w_001_006);
  nand2 I008_576(w_008_576, w_001_009, w_005_044);
  not1 I008_577(w_008_577, w_004_148);
  and2 I008_580(w_008_580, w_003_030, w_006_213);
  nand2 I008_581(w_008_581, w_003_051, w_005_190);
  nand2 I008_582(w_008_582, w_006_202, w_007_270);
  and2 I008_583(w_008_583, w_004_186, w_003_050);
  not1 I008_584(w_008_584, w_003_075);
  not1 I008_585(w_008_585, w_007_074);
  and2 I008_587(w_008_587, w_006_249, w_003_059);
  or2  I008_588(w_008_588, w_002_674, w_005_008);
  nand2 I008_589(w_008_589, w_003_010, w_005_228);
  or2  I008_590(w_008_590, w_005_184, w_005_056);
  not1 I008_591(w_008_591, w_005_072);
  or2  I008_592(w_008_592, w_005_205, w_005_132);
  not1 I008_594(w_008_594, w_006_091);
  not1 I008_595(w_008_595, w_005_114);
  or2  I008_598(w_008_598, w_006_244, w_005_076);
  and2 I008_601(w_008_601, w_000_186, w_005_081);
  and2 I008_602(w_008_602, w_005_001, w_005_231);
  or2  I008_603(w_008_603, w_004_246, w_000_370);
  or2  I008_604(w_008_604, w_005_230, w_006_118);
  nand2 I008_605(w_008_605, w_003_063, w_007_059);
  and2 I008_608(w_008_608, w_002_656, w_004_129);
  or2  I008_610(w_008_610, w_007_033, w_006_031);
  nand2 I008_611(w_008_611, w_005_208, w_006_003);
  not1 I008_612(w_008_612, w_005_029);
  or2  I008_613(w_008_613, w_003_000, w_002_084);
  or2  I008_614(w_008_614, w_007_021, w_001_012);
  or2  I008_615(w_008_615, w_006_031, w_006_038);
  and2 I008_616(w_008_616, w_004_048, w_005_052);
  or2  I008_619(w_008_619, w_004_285, w_000_254);
  or2  I008_620(w_008_620, w_006_078, w_006_213);
  nand2 I008_621(w_008_621, w_003_057, w_000_609);
  or2  I008_622(w_008_622, w_000_262, w_004_288);
  or2  I008_623(w_008_623, w_003_007, w_001_021);
  nand2 I008_624(w_008_624, w_001_036, w_004_152);
  and2 I008_625(w_008_625, w_001_007, w_006_208);
  not1 I008_626(w_008_626, w_007_296);
  or2  I008_628(w_008_628, w_000_139, w_002_233);
  or2  I008_629(w_008_629, w_006_231, w_002_050);
  or2  I008_636(w_008_636, w_006_107, w_006_096);
  nand2 I008_637(w_008_637, w_002_344, w_002_562);
  or2  I008_638(w_008_638, w_005_213, w_007_022);
  and2 I008_639(w_008_639, w_003_038, w_004_015);
  or2  I008_640(w_008_640, w_000_372, w_005_145);
  not1 I008_644(w_008_644, w_002_423);
  nand2 I008_645(w_008_645, w_001_020, w_003_071);
  nand2 I008_646(w_008_646, w_000_524, w_000_560);
  and2 I008_647(w_008_647, w_005_224, w_001_011);
  and2 I008_648(w_008_648, w_000_337, w_001_012);
  not1 I008_650(w_008_650, w_006_115);
  and2 I008_651(w_008_651, w_000_090, w_003_084);
  not1 I008_653(w_008_653, w_003_058);
  not1 I008_654(w_008_654, w_001_034);
  and2 I008_656(w_008_656, w_007_228, w_006_221);
  or2  I008_657(w_008_657, w_007_045, w_003_059);
  and2 I008_658(w_008_658, w_003_076, w_003_016);
  or2  I008_659(w_008_659, w_002_044, w_000_009);
  or2  I008_661(w_008_661, w_004_072, w_004_157);
  nand2 I008_662(w_008_662, w_000_379, w_000_439);
  nand2 I008_663(w_008_663, w_006_213, w_004_055);
  and2 I008_664(w_008_664, w_007_176, w_004_244);
  not1 I008_665(w_008_665, w_000_056);
  nand2 I008_666(w_008_666, w_002_012, w_003_052);
  nand2 I008_668(w_008_668, w_003_060, w_000_661);
  and2 I008_669(w_008_669, w_000_662, w_000_503);
  and2 I008_674(w_008_674, w_006_078, w_007_473);
  and2 I008_676(w_008_676, w_005_176, w_000_123);
  nand2 I008_677(w_008_677, w_004_302, w_004_463);
  not1 I008_678(w_008_678, w_002_477);
  and2 I008_679(w_008_679, w_007_098, w_001_035);
  and2 I008_680(w_008_680, w_001_012, w_000_256);
  and2 I008_681(w_008_681, w_007_247, w_001_021);
  or2  I008_682(w_008_682, w_006_129, w_001_010);
  or2  I008_683(w_008_683, w_002_462, w_001_010);
  nand2 I008_685(w_008_685, w_003_058, w_005_103);
  not1 I008_686(w_008_686, w_001_009);
  not1 I008_688(w_008_688, w_001_006);
  not1 I008_692(w_008_692, w_001_034);
  not1 I008_693(w_008_693, w_004_365);
  or2  I008_694(w_008_694, w_001_029, w_007_155);
  or2  I008_696(w_008_696, w_007_108, w_005_288);
  nand2 I008_697(w_008_697, w_004_204, w_003_076);
  nand2 I008_698(w_008_698, w_001_022, w_002_116);
  nand2 I008_699(w_008_699, w_003_053, w_001_005);
  not1 I008_700(w_008_700, w_002_088);
  and2 I008_701(w_008_701, w_002_595, w_005_003);
  and2 I008_702(w_008_702, w_004_021, w_005_157);
  or2  I008_703(w_008_703, w_003_028, w_005_097);
  or2  I008_704(w_008_704, w_000_666, w_004_020);
  or2  I008_707(w_008_707, w_002_345, w_004_025);
  or2  I008_708(w_008_708, w_004_459, w_000_610);
  not1 I008_709(w_008_709, w_001_009);
  or2  I008_710(w_008_710, w_006_234, w_007_005);
  nand2 I008_711(w_008_711, w_003_059, w_007_000);
  and2 I008_713(w_008_713, w_000_423, w_005_107);
  and2 I008_714(w_008_714, w_001_013, w_005_111);
  not1 I008_715(w_008_715, w_005_240);
  or2  I008_718(w_008_718, w_003_011, w_004_021);
  not1 I008_719(w_008_719, w_007_203);
  not1 I008_720(w_008_720, w_007_178);
  nand2 I008_721(w_008_721, w_002_628, w_000_629);
  not1 I008_722(w_008_722, w_006_230);
  or2  I008_724(w_008_724, w_004_214, w_002_040);
  and2 I008_725(w_008_725, w_003_038, w_003_031);
  not1 I008_726(w_008_726, w_001_006);
  or2  I008_727(w_008_727, w_006_131, w_001_008);
  and2 I008_728(w_008_728, w_003_007, w_005_216);
  and2 I008_729(w_008_729, w_003_019, w_000_066);
  nand2 I008_730(w_008_730, w_006_157, w_000_170);
  not1 I008_733(w_008_733, w_003_082);
  not1 I008_735(w_008_735, w_007_425);
  or2  I008_737(w_008_737, w_005_152, w_003_032);
  and2 I008_738(w_008_738, w_001_022, w_007_027);
  nand2 I008_740(w_008_740, w_005_175, w_002_044);
  not1 I008_742(w_008_742, w_003_040);
  and2 I008_743(w_008_743, w_005_283, w_001_006);
  and2 I008_745(w_008_745, w_003_020, w_000_229);
  not1 I008_746(w_008_746, w_002_216);
  not1 I008_747(w_008_747, w_007_263);
  and2 I008_748(w_008_748, w_004_090, w_004_053);
  and2 I008_749(w_008_749, w_002_055, w_007_284);
  nand2 I008_750(w_008_750, w_004_120, w_000_094);
  and2 I008_751(w_008_751, w_005_129, w_005_156);
  nand2 I008_753(w_008_753, w_007_438, w_005_015);
  and2 I008_755(w_008_755, w_004_488, w_007_323);
  nand2 I008_757(w_008_757, w_006_061, w_007_266);
  nand2 I008_758(w_008_758, w_004_423, w_004_103);
  or2  I008_760(w_008_760, w_004_376, w_007_333);
  nand2 I008_762(w_008_762, w_002_494, w_001_028);
  or2  I008_763(w_008_763, w_000_255, w_002_552);
  not1 I008_766(w_008_768, w_008_767);
  or2  I008_767(w_008_769, w_002_073, w_008_768);
  nand2 I008_768(w_008_770, w_008_769, w_008_786);
  nand2 I008_769(w_008_771, w_008_770, w_006_092);
  or2  I008_770(w_008_772, w_008_771, w_006_085);
  and2 I008_771(w_008_773, w_001_032, w_008_772);
  or2  I008_772(w_008_767, w_007_180, w_008_773);
  or2  I008_773(w_008_778, w_008_777, w_001_006);
  and2 I008_774(w_008_779, w_004_215, w_008_778);
  not1 I008_775(w_008_780, w_008_779);
  not1 I008_776(w_008_781, w_008_780);
  or2  I008_777(w_008_782, w_008_781, w_001_013);
  or2  I008_778(w_008_783, w_008_782, w_001_031);
  and2 I008_779(w_008_784, w_004_473, w_008_783);
  not1 I008_780(w_008_777, w_008_770);
  and2 I008_781(w_008_786, w_005_143, w_008_784);
  not1 I009_000(w_009_000, w_008_650);
  or2  I009_001(w_009_001, w_008_357, w_002_042);
  not1 I009_003(w_009_003, w_007_256);
  nand2 I009_004(w_009_004, w_007_012, w_004_230);
  not1 I009_005(w_009_005, w_005_122);
  and2 I009_006(w_009_006, w_003_042, w_005_123);
  and2 I009_007(w_009_007, w_005_048, w_008_167);
  not1 I009_009(w_009_009, w_008_740);
  or2  I009_010(w_009_010, w_005_042, w_008_662);
  or2  I009_011(w_009_011, w_006_169, w_000_358);
  or2  I009_012(w_009_012, w_004_319, w_004_449);
  not1 I009_013(w_009_013, w_007_280);
  not1 I009_014(w_009_014, w_003_002);
  and2 I009_015(w_009_015, w_005_167, w_000_603);
  nand2 I009_016(w_009_016, w_002_033, w_003_031);
  not1 I009_017(w_009_017, w_007_017);
  and2 I009_018(w_009_018, w_007_004, w_001_012);
  or2  I009_019(w_009_019, w_004_069, w_008_118);
  not1 I009_020(w_009_020, w_004_054);
  nand2 I009_021(w_009_021, w_004_200, w_003_068);
  nand2 I009_022(w_009_022, w_008_725, w_004_029);
  and2 I009_023(w_009_023, w_007_124, w_003_042);
  not1 I009_024(w_009_024, w_008_348);
  not1 I009_025(w_009_025, w_005_067);
  nand2 I009_026(w_009_026, w_007_100, w_005_225);
  nand2 I009_027(w_009_027, w_006_134, w_007_424);
  nand2 I009_028(w_009_028, w_002_686, w_006_210);
  or2  I009_029(w_009_029, w_003_046, w_007_028);
  or2  I009_030(w_009_030, w_005_152, w_008_076);
  not1 I009_031(w_009_031, w_006_172);
  or2  I009_032(w_009_032, w_002_330, w_004_185);
  and2 I009_033(w_009_033, w_007_120, w_008_686);
  and2 I009_035(w_009_035, w_003_013, w_000_589);
  not1 I009_036(w_009_036, w_007_135);
  nand2 I009_037(w_009_037, w_001_025, w_000_507);
  nand2 I009_038(w_009_038, w_004_484, w_002_008);
  not1 I009_040(w_009_040, w_002_016);
  or2  I009_041(w_009_041, w_006_029, w_006_014);
  nand2 I009_042(w_009_042, w_004_115, w_008_524);
  or2  I009_043(w_009_043, w_005_271, w_006_001);
  not1 I009_044(w_009_044, w_007_192);
  or2  I009_045(w_009_045, w_003_057, w_004_408);
  not1 I009_046(w_009_046, w_008_008);
  not1 I009_047(w_009_047, w_004_453);
  or2  I009_048(w_009_048, w_005_036, w_006_101);
  and2 I009_049(w_009_049, w_001_033, w_008_587);
  nand2 I009_050(w_009_050, w_007_134, w_000_574);
  or2  I009_051(w_009_051, w_003_018, w_003_066);
  not1 I009_052(w_009_052, w_006_235);
  and2 I009_053(w_009_053, w_005_129, w_001_031);
  and2 I009_054(w_009_054, w_005_161, w_003_074);
  not1 I009_055(w_009_055, w_000_260);
  not1 I009_056(w_009_056, w_008_552);
  not1 I009_058(w_009_058, w_001_032);
  not1 I009_059(w_009_059, w_000_071);
  and2 I009_060(w_009_060, w_000_164, w_006_090);
  and2 I009_061(w_009_061, w_000_108, w_005_261);
  nand2 I009_062(w_009_062, w_005_063, w_004_120);
  not1 I009_064(w_009_064, w_004_223);
  nand2 I009_065(w_009_065, w_004_223, w_003_058);
  and2 I009_066(w_009_066, w_004_214, w_004_466);
  or2  I009_068(w_009_068, w_004_213, w_006_219);
  nand2 I009_070(w_009_070, w_004_192, w_007_209);
  and2 I009_071(w_009_071, w_000_667, w_008_318);
  not1 I009_072(w_009_072, w_001_005);
  not1 I009_073(w_009_073, w_003_022);
  not1 I009_074(w_009_074, w_005_121);
  nand2 I009_075(w_009_075, w_005_297, w_002_661);
  or2  I009_076(w_009_076, w_008_390, w_004_042);
  or2  I009_077(w_009_077, w_001_024, w_008_626);
  and2 I009_078(w_009_078, w_004_222, w_003_061);
  not1 I009_079(w_009_079, w_008_683);
  and2 I009_080(w_009_080, w_007_221, w_004_038);
  nand2 I009_081(w_009_081, w_000_188, w_007_400);
  or2  I009_082(w_009_082, w_007_131, w_001_020);
  nand2 I009_083(w_009_083, w_006_101, w_001_020);
  and2 I009_084(w_009_084, w_000_605, w_000_036);
  and2 I009_085(w_009_085, w_003_024, w_001_030);
  and2 I009_086(w_009_086, w_002_389, w_006_024);
  or2  I009_087(w_009_087, w_000_543, w_005_137);
  nand2 I009_088(w_009_088, w_001_013, w_000_349);
  not1 I009_089(w_009_089, w_005_182);
  or2  I009_090(w_009_090, w_004_128, w_004_372);
  not1 I009_091(w_009_091, w_004_250);
  not1 I009_092(w_009_092, w_005_090);
  and2 I009_093(w_009_093, w_006_235, w_007_379);
  not1 I009_094(w_009_094, w_004_068);
  not1 I009_095(w_009_095, w_008_298);
  or2  I009_096(w_009_096, w_006_212, w_000_387);
  or2  I009_097(w_009_097, w_000_355, w_005_263);
  and2 I009_098(w_009_098, w_007_166, w_006_075);
  or2  I009_099(w_009_099, w_003_010, w_008_613);
  nand2 I009_100(w_009_100, w_005_235, w_008_506);
  and2 I009_101(w_009_101, w_003_042, w_008_078);
  or2  I009_102(w_009_102, w_006_157, w_006_031);
  and2 I009_103(w_009_103, w_005_163, w_005_117);
  not1 I009_104(w_009_104, w_006_159);
  not1 I009_105(w_009_105, w_003_035);
  and2 I009_106(w_009_106, w_004_130, w_003_001);
  nand2 I009_107(w_009_107, w_006_028, w_007_460);
  nand2 I009_108(w_009_108, w_001_032, w_000_068);
  and2 I009_109(w_009_109, w_004_067, w_002_685);
  not1 I009_110(w_009_110, w_007_238);
  not1 I009_111(w_009_111, w_007_088);
  not1 I009_113(w_009_113, w_005_052);
  not1 I009_114(w_009_114, w_003_009);
  nand2 I009_115(w_009_115, w_003_036, w_007_278);
  and2 I009_116(w_009_116, w_008_751, w_008_298);
  nand2 I009_117(w_009_117, w_004_190, w_002_692);
  or2  I009_118(w_009_118, w_008_501, w_005_063);
  nand2 I009_119(w_009_119, w_008_103, w_005_096);
  or2  I009_120(w_009_120, w_001_000, w_000_582);
  nand2 I009_121(w_009_121, w_005_279, w_005_161);
  not1 I009_122(w_009_122, w_006_077);
  or2  I009_123(w_009_123, w_005_056, w_005_234);
  nand2 I009_124(w_009_124, w_005_159, w_001_009);
  not1 I009_125(w_009_125, w_004_058);
  or2  I009_126(w_009_126, w_002_513, w_003_043);
  not1 I009_127(w_009_127, w_002_086);
  or2  I009_128(w_009_128, w_005_154, w_005_232);
  and2 I009_129(w_009_129, w_008_343, w_008_676);
  and2 I009_130(w_009_130, w_004_093, w_004_434);
  nand2 I009_131(w_009_131, w_000_432, w_000_668);
  not1 I009_132(w_009_132, w_002_290);
  and2 I009_133(w_009_133, w_004_003, w_006_217);
  or2  I009_134(w_009_134, w_008_469, w_006_032);
  not1 I009_135(w_009_135, w_002_058);
  nand2 I009_136(w_009_136, w_008_665, w_000_024);
  not1 I009_137(w_009_137, w_003_033);
  nand2 I009_138(w_009_138, w_005_259, w_003_064);
  nand2 I009_139(w_009_139, w_003_037, w_002_362);
  or2  I009_140(w_009_140, w_007_235, w_003_043);
  nand2 I009_141(w_009_141, w_002_489, w_007_073);
  and2 I009_142(w_009_142, w_008_044, w_006_182);
  or2  I009_143(w_009_143, w_006_207, w_003_080);
  and2 I009_144(w_009_144, w_006_250, w_000_390);
  not1 I009_145(w_009_145, w_000_461);
  nand2 I009_146(w_009_146, w_002_375, w_005_129);
  or2  I009_147(w_009_147, w_006_092, w_004_242);
  or2  I009_149(w_009_149, w_002_020, w_003_084);
  and2 I009_150(w_009_150, w_004_469, w_003_007);
  or2  I009_151(w_009_151, w_001_033, w_002_629);
  or2  I009_152(w_009_152, w_008_760, w_005_301);
  not1 I009_153(w_009_153, w_008_588);
  and2 I009_154(w_009_154, w_003_007, w_008_025);
  not1 I009_155(w_009_155, w_003_035);
  nand2 I009_156(w_009_156, w_003_055, w_000_493);
  and2 I009_158(w_009_158, w_001_004, w_003_003);
  nand2 I009_159(w_009_159, w_003_061, w_006_215);
  not1 I009_160(w_009_160, w_004_256);
  not1 I009_161(w_009_161, w_005_063);
  or2  I009_162(w_009_162, w_000_371, w_003_006);
  not1 I009_163(w_009_163, w_007_066);
  or2  I009_164(w_009_164, w_006_022, w_002_574);
  nand2 I009_166(w_009_166, w_008_073, w_001_000);
  or2  I009_167(w_009_167, w_005_287, w_007_156);
  or2  I009_168(w_009_168, w_003_057, w_007_010);
  and2 I009_169(w_009_169, w_001_019, w_006_168);
  and2 I009_172(w_009_172, w_000_138, w_000_337);
  and2 I009_173(w_009_173, w_003_067, w_005_090);
  nand2 I009_175(w_009_175, w_001_005, w_006_075);
  or2  I009_176(w_009_176, w_001_013, w_007_235);
  or2  I009_177(w_009_177, w_002_024, w_003_084);
  not1 I009_180(w_009_180, w_006_017);
  nand2 I009_181(w_009_181, w_006_191, w_008_381);
  and2 I009_182(w_009_182, w_003_007, w_008_399);
  not1 I009_183(w_009_183, w_004_317);
  nand2 I009_184(w_009_184, w_006_099, w_008_152);
  nand2 I009_185(w_009_185, w_004_126, w_006_049);
  not1 I009_186(w_009_186, w_007_342);
  not1 I009_189(w_009_189, w_002_571);
  and2 I009_190(w_009_190, w_002_340, w_005_027);
  nand2 I009_191(w_009_191, w_002_696, w_008_290);
  and2 I009_193(w_009_193, w_003_042, w_003_044);
  nand2 I009_194(w_009_194, w_003_033, w_007_068);
  nand2 I009_196(w_009_196, w_006_214, w_002_635);
  and2 I009_197(w_009_197, w_005_000, w_004_099);
  or2  I009_198(w_009_198, w_006_126, w_007_474);
  nand2 I009_199(w_009_199, w_003_007, w_000_445);
  nand2 I009_200(w_009_200, w_008_459, w_003_015);
  not1 I009_208(w_009_208, w_000_613);
  or2  I009_209(w_009_209, w_008_419, w_004_281);
  and2 I009_210(w_009_210, w_006_032, w_003_019);
  not1 I009_211(w_009_211, w_006_212);
  nand2 I009_213(w_009_213, w_007_136, w_006_083);
  and2 I009_214(w_009_214, w_003_056, w_004_204);
  or2  I009_215(w_009_215, w_003_017, w_003_079);
  or2  I009_216(w_009_216, w_008_240, w_000_030);
  nand2 I009_217(w_009_217, w_004_134, w_003_078);
  nand2 I009_219(w_009_219, w_008_225, w_002_685);
  or2  I009_220(w_009_220, w_008_346, w_002_196);
  not1 I009_221(w_009_221, w_003_024);
  nand2 I009_222(w_009_222, w_007_420, w_005_004);
  and2 I009_223(w_009_223, w_006_100, w_004_273);
  not1 I009_224(w_009_224, w_007_221);
  or2  I009_226(w_009_226, w_006_231, w_008_762);
  nand2 I009_228(w_009_228, w_001_015, w_001_012);
  not1 I009_229(w_009_229, w_004_371);
  not1 I009_230(w_009_230, w_007_480);
  or2  I009_231(w_009_231, w_001_007, w_000_165);
  nand2 I009_232(w_009_232, w_007_124, w_007_209);
  nand2 I009_233(w_009_233, w_007_066, w_007_118);
  not1 I009_234(w_009_234, w_004_222);
  not1 I009_235(w_009_235, w_002_193);
  and2 I009_236(w_009_236, w_003_021, w_004_074);
  nand2 I009_237(w_009_237, w_005_213, w_000_436);
  or2  I009_238(w_009_238, w_001_032, w_007_098);
  or2  I009_239(w_009_239, w_004_256, w_008_023);
  nand2 I009_240(w_009_240, w_006_065, w_001_014);
  or2  I009_241(w_009_241, w_004_384, w_007_059);
  nand2 I009_243(w_009_243, w_004_165, w_007_437);
  or2  I009_244(w_009_244, w_005_073, w_000_437);
  nand2 I009_245(w_009_245, w_006_029, w_002_590);
  nand2 I009_246(w_009_246, w_001_021, w_005_103);
  and2 I009_247(w_009_247, w_005_104, w_003_078);
  and2 I009_248(w_009_248, w_001_019, w_001_005);
  not1 I009_249(w_009_249, w_007_041);
  nand2 I009_250(w_009_250, w_004_160, w_007_178);
  or2  I009_251(w_009_251, w_005_297, w_000_349);
  and2 I009_253(w_009_253, w_001_024, w_006_144);
  not1 I009_255(w_009_255, w_005_305);
  nand2 I009_258(w_009_258, w_000_658, w_005_193);
  or2  I009_259(w_009_259, w_001_035, w_005_093);
  or2  I009_260(w_009_260, w_002_490, w_001_027);
  not1 I009_264(w_009_264, w_006_247);
  and2 I009_265(w_009_265, w_008_220, w_003_064);
  and2 I009_267(w_009_267, w_004_176, w_005_211);
  not1 I009_268(w_009_268, w_007_202);
  or2  I009_270(w_009_270, w_006_216, w_006_215);
  or2  I009_271(w_009_271, w_001_009, w_008_711);
  nand2 I009_272(w_009_272, w_002_327, w_001_007);
  or2  I009_273(w_009_273, w_001_017, w_006_154);
  or2  I009_274(w_009_274, w_003_066, w_006_134);
  and2 I009_279(w_009_279, w_001_012, w_007_308);
  or2  I009_281(w_009_281, w_001_023, w_000_257);
  nand2 I009_283(w_009_283, w_001_032, w_000_461);
  nand2 I009_284(w_009_284, w_008_196, w_006_033);
  or2  I009_288(w_009_288, w_008_504, w_007_288);
  or2  I009_293(w_009_293, w_002_400, w_004_051);
  nand2 I009_294(w_009_294, w_003_082, w_001_035);
  not1 I009_295(w_009_295, w_006_199);
  nand2 I009_296(w_009_296, w_005_216, w_002_264);
  and2 I009_297(w_009_297, w_005_294, w_000_665);
  nand2 I009_300(w_009_300, w_003_074, w_000_675);
  or2  I009_301(w_009_301, w_008_331, w_005_087);
  nand2 I009_302(w_009_302, w_006_169, w_002_246);
  not1 I009_303(w_009_303, w_008_644);
  or2  I009_305(w_009_305, w_006_062, w_003_067);
  and2 I009_308(w_009_308, w_000_175, w_004_259);
  nand2 I009_310(w_009_310, w_000_607, w_006_017);
  nand2 I009_313(w_009_313, w_007_185, w_000_431);
  not1 I009_314(w_009_314, w_006_158);
  or2  I009_315(w_009_315, w_002_127, w_004_193);
  nand2 I009_316(w_009_316, w_008_621, w_008_498);
  and2 I009_317(w_009_317, w_004_067, w_007_092);
  nand2 I009_318(w_009_318, w_007_091, w_004_277);
  nand2 I009_320(w_009_320, w_004_440, w_005_037);
  not1 I009_321(w_009_321, w_003_006);
  or2  I009_322(w_009_322, w_005_156, w_005_137);
  not1 I009_325(w_009_325, w_002_267);
  nand2 I009_326(w_009_326, w_004_279, w_003_084);
  and2 I009_328(w_009_328, w_005_227, w_004_241);
  or2  I009_329(w_009_329, w_001_027, w_002_673);
  nand2 I009_330(w_009_330, w_000_587, w_006_237);
  or2  I009_331(w_009_331, w_005_223, w_007_272);
  and2 I009_333(w_009_333, w_005_238, w_008_099);
  nand2 I009_335(w_009_335, w_002_091, w_000_367);
  or2  I009_336(w_009_336, w_003_070, w_007_361);
  nand2 I009_337(w_009_337, w_005_018, w_001_017);
  nand2 I009_338(w_009_338, w_008_656, w_006_239);
  not1 I009_340(w_009_340, w_007_246);
  nand2 I009_341(w_009_341, w_003_068, w_003_078);
  or2  I009_342(w_009_342, w_004_105, w_004_460);
  and2 I009_343(w_009_343, w_003_021, w_007_114);
  or2  I009_344(w_009_344, w_006_245, w_004_289);
  not1 I009_345(w_009_345, w_001_006);
  not1 I009_350(w_009_350, w_001_013);
  or2  I009_351(w_009_351, w_000_575, w_008_484);
  or2  I009_353(w_009_353, w_005_004, w_000_097);
  nand2 I009_354(w_009_354, w_004_244, w_003_066);
  and2 I009_357(w_009_357, w_001_016, w_003_041);
  nand2 I009_359(w_009_359, w_005_032, w_004_375);
  and2 I009_360(w_009_360, w_004_472, w_007_002);
  not1 I009_361(w_009_361, w_001_010);
  nand2 I009_362(w_009_362, w_003_081, w_006_155);
  not1 I009_363(w_009_363, w_006_028);
  not1 I009_364(w_009_364, w_008_657);
  nand2 I009_365(w_009_365, w_007_074, w_001_023);
  nand2 I009_366(w_009_366, w_002_316, w_003_016);
  and2 I009_368(w_009_368, w_008_485, w_003_031);
  and2 I009_369(w_009_369, w_005_054, w_008_446);
  and2 I009_370(w_009_370, w_004_022, w_002_043);
  or2  I009_371(w_009_371, w_005_232, w_008_031);
  and2 I009_372(w_009_372, w_006_232, w_002_695);
  not1 I009_373(w_009_373, w_000_377);
  not1 I009_374(w_009_374, w_000_532);
  not1 I009_375(w_009_375, w_006_217);
  or2  I009_376(w_009_376, w_004_015, w_004_118);
  nand2 I009_377(w_009_377, w_002_045, w_008_044);
  nand2 I009_378(w_009_378, w_000_434, w_001_003);
  and2 I009_379(w_009_379, w_005_033, w_007_437);
  or2  I009_380(w_009_380, w_007_091, w_005_227);
  nand2 I009_382(w_009_382, w_001_017, w_004_435);
  or2  I009_383(w_009_383, w_008_747, w_007_321);
  and2 I009_384(w_009_384, w_002_106, w_008_103);
  not1 I009_388(w_009_388, w_004_206);
  nand2 I009_389(w_009_389, w_007_159, w_005_015);
  or2  I009_390(w_009_390, w_001_023, w_007_425);
  not1 I009_391(w_009_391, w_006_023);
  or2  I009_392(w_009_392, w_006_177, w_008_156);
  not1 I009_393(w_009_393, w_002_259);
  and2 I009_394(w_009_394, w_001_035, w_004_040);
  and2 I009_395(w_009_395, w_004_051, w_004_311);
  and2 I009_396(w_009_396, w_002_505, w_006_055);
  not1 I009_397(w_009_397, w_008_516);
  nand2 I009_398(w_009_398, w_002_383, w_001_028);
  and2 I009_399(w_009_399, w_007_166, w_005_085);
  nand2 I009_402(w_009_402, w_000_088, w_004_115);
  or2  I009_403(w_009_403, w_001_022, w_002_006);
  not1 I009_404(w_009_404, w_008_209);
  or2  I009_405(w_009_405, w_000_140, w_008_083);
  nand2 I009_406(w_009_406, w_004_006, w_004_452);
  and2 I009_407(w_009_407, w_005_042, w_001_027);
  nand2 I009_408(w_009_408, w_004_242, w_003_049);
  nand2 I009_411(w_009_411, w_005_080, w_007_064);
  or2  I009_412(w_009_412, w_004_357, w_005_059);
  not1 I009_414(w_009_414, w_008_162);
  or2  I009_415(w_009_415, w_001_022, w_002_622);
  not1 I009_416(w_009_416, w_000_666);
  nand2 I009_417(w_009_417, w_005_077, w_004_199);
  nand2 I009_418(w_009_418, w_005_046, w_000_387);
  nand2 I009_420(w_009_420, w_002_061, w_007_114);
  and2 I009_421(w_009_421, w_007_310, w_000_389);
  and2 I009_422(w_009_422, w_002_212, w_002_648);
  not1 I009_423(w_009_423, w_002_078);
  not1 I009_424(w_009_424, w_006_251);
  not1 I009_426(w_009_426, w_004_040);
  and2 I009_427(w_009_427, w_008_272, w_003_022);
  not1 I009_428(w_009_428, w_002_038);
  or2  I009_430(w_009_430, w_000_229, w_007_154);
  not1 I009_432(w_009_432, w_002_534);
  not1 I009_433(w_009_433, w_003_026);
  not1 I009_435(w_009_435, w_004_104);
  not1 I009_438(w_009_438, w_000_250);
  nand2 I009_439(w_009_439, w_005_086, w_003_038);
  not1 I009_440(w_009_440, w_006_218);
  or2  I009_441(w_009_441, w_008_557, w_000_260);
  and2 I009_442(w_009_442, w_005_088, w_004_145);
  or2  I009_443(w_009_443, w_006_137, w_005_087);
  not1 I009_444(w_009_444, w_004_269);
  or2  I009_445(w_009_445, w_003_066, w_007_014);
  and2 I009_446(w_009_446, w_002_583, w_001_020);
  and2 I009_448(w_009_448, w_008_210, w_007_296);
  and2 I009_449(w_009_449, w_002_186, w_004_188);
  not1 I009_451(w_009_451, w_003_000);
  nand2 I009_452(w_009_452, w_001_000, w_003_071);
  and2 I009_455(w_009_455, w_001_015, w_002_351);
  not1 I009_456(w_009_456, w_005_250);
  not1 I009_460(w_009_460, w_001_031);
  or2  I009_462(w_009_462, w_001_024, w_001_009);
  nand2 I009_463(w_009_463, w_002_243, w_007_180);
  or2  I009_464(w_009_464, w_002_606, w_002_449);
  not1 I009_465(w_009_465, w_002_626);
  not1 I009_468(w_009_468, w_002_042);
  nand2 I009_469(w_009_469, w_002_233, w_005_210);
  and2 I009_470(w_009_470, w_008_454, w_004_001);
  nand2 I009_471(w_009_471, w_004_097, w_001_013);
  or2  I009_472(w_009_472, w_002_061, w_004_296);
  not1 I009_473(w_009_473, w_001_018);
  and2 I009_476(w_009_476, w_004_038, w_002_568);
  not1 I009_478(w_009_478, w_006_028);
  nand2 I009_479(w_009_479, w_007_092, w_008_031);
  or2  I009_480(w_009_480, w_000_099, w_000_383);
  or2  I009_481(w_009_481, w_006_251, w_005_316);
  not1 I009_482(w_009_482, w_005_183);
  not1 I009_483(w_009_483, w_000_283);
  not1 I009_485(w_009_485, w_001_021);
  not1 I009_486(w_009_486, w_001_005);
  not1 I009_487(w_009_487, w_000_074);
  nand2 I009_488(w_009_488, w_008_610, w_001_025);
  or2  I009_489(w_009_489, w_005_138, w_003_078);
  and2 I009_490(w_009_490, w_007_181, w_002_295);
  or2  I009_491(w_009_491, w_004_077, w_007_308);
  nand2 I009_492(w_009_492, w_007_032, w_004_375);
  not1 I009_493(w_009_493, w_006_056);
  and2 I009_497(w_009_497, w_003_024, w_001_020);
  or2  I009_498(w_009_498, w_005_155, w_003_031);
  or2  I009_499(w_009_499, w_002_380, w_002_128);
  nand2 I009_500(w_009_500, w_006_184, w_008_169);
  not1 I009_501(w_009_501, w_004_091);
  and2 I009_502(w_009_502, w_008_035, w_008_047);
  nand2 I009_503(w_009_503, w_006_054, w_001_036);
  and2 I009_504(w_009_504, w_000_440, w_001_019);
  not1 I009_505(w_009_505, w_004_122);
  not1 I009_507(w_009_507, w_008_585);
  or2  I009_508(w_009_508, w_007_182, w_001_007);
  and2 I009_509(w_009_509, w_000_542, w_008_748);
  or2  I009_510(w_009_510, w_004_060, w_003_040);
  and2 I009_512(w_009_512, w_006_235, w_000_069);
  nand2 I009_513(w_009_513, w_002_316, w_008_316);
  not1 I009_515(w_009_515, w_000_182);
  not1 I009_516(w_009_516, w_008_724);
  nand2 I009_517(w_009_517, w_000_325, w_000_602);
  and2 I009_520(w_009_520, w_008_143, w_006_000);
  and2 I009_521(w_009_521, w_006_073, w_004_245);
  not1 I009_522(w_009_522, w_007_142);
  not1 I009_523(w_009_523, w_007_164);
  and2 I009_524(w_009_524, w_005_086, w_007_042);
  not1 I009_525(w_009_525, w_002_688);
  and2 I009_527(w_009_527, w_004_502, w_008_282);
  nand2 I009_528(w_009_528, w_008_398, w_002_043);
  nand2 I009_529(w_009_529, w_007_116, w_004_103);
  not1 I009_531(w_009_531, w_008_589);
  and2 I009_532(w_009_532, w_000_478, w_002_620);
  or2  I009_533(w_009_533, w_004_167, w_007_019);
  and2 I009_536(w_009_536, w_002_113, w_008_029);
  not1 I009_537(w_009_537, w_008_576);
  nand2 I009_539(w_009_539, w_006_033, w_002_005);
  not1 I009_540(w_009_540, w_000_288);
  nand2 I009_541(w_009_541, w_005_174, w_000_187);
  or2  I009_542(w_009_542, w_007_390, w_000_059);
  not1 I009_543(w_009_543, w_000_172);
  not1 I009_545(w_009_545, w_005_193);
  nand2 I009_546(w_009_546, w_002_459, w_007_272);
  and2 I009_547(w_009_547, w_005_178, w_008_090);
  or2  I009_549(w_009_549, w_003_053, w_003_021);
  nand2 I009_550(w_009_550, w_003_024, w_004_221);
  nand2 I009_551(w_009_551, w_002_367, w_001_000);
  nand2 I009_552(w_009_552, w_000_510, w_004_089);
  not1 I009_553(w_009_553, w_002_691);
  and2 I009_554(w_009_554, w_001_005, w_000_270);
  not1 I009_555(w_009_555, w_005_273);
  nand2 I009_556(w_009_556, w_008_218, w_003_083);
  or2  I009_557(w_009_557, w_006_169, w_004_229);
  or2  I009_558(w_009_558, w_006_054, w_002_543);
  or2  I009_560(w_009_560, w_007_139, w_005_081);
  nand2 I009_561(w_009_561, w_004_063, w_001_008);
  or2  I009_562(w_009_562, w_006_166, w_007_396);
  and2 I009_563(w_009_563, w_001_005, w_001_025);
  not1 I009_564(w_009_564, w_005_035);
  nand2 I009_568(w_009_568, w_006_054, w_006_189);
  not1 I009_570(w_009_570, w_007_127);
  and2 I009_571(w_009_571, w_001_000, w_006_156);
  not1 I009_572(w_009_572, w_004_012);
  or2  I009_573(w_009_573, w_004_188, w_002_514);
  or2  I009_574(w_009_574, w_005_188, w_000_630);
  not1 I009_579(w_009_579, w_006_105);
  and2 I009_581(w_009_581, w_000_092, w_007_122);
  and2 I009_583(w_009_583, w_003_084, w_008_413);
  nand2 I009_584(w_009_584, w_003_081, w_000_583);
  or2  I009_591(w_009_591, w_003_007, w_008_743);
  nand2 I009_594(w_009_594, w_005_083, w_001_035);
  or2  I009_597(w_009_597, w_002_017, w_002_054);
  and2 I009_598(w_009_598, w_000_576, w_000_312);
  or2  I009_600(w_009_600, w_001_017, w_000_557);
  nand2 I009_601(w_009_601, w_006_198, w_001_029);
  nand2 I009_602(w_009_602, w_005_009, w_002_061);
  and2 I009_603(w_009_603, w_006_022, w_004_188);
  nand2 I009_604(w_009_604, w_002_677, w_000_602);
  not1 I009_606(w_009_606, w_008_638);
  not1 I009_607(w_009_607, w_007_265);
  not1 I009_609(w_009_609, w_008_645);
  and2 I009_610(w_009_610, w_006_007, w_000_381);
  nand2 I009_611(w_009_611, w_006_010, w_005_131);
  and2 I009_612(w_009_612, w_006_191, w_007_159);
  or2  I009_614(w_009_614, w_004_439, w_006_007);
  or2  I009_616(w_009_616, w_003_041, w_004_466);
  nand2 I009_619(w_009_619, w_002_271, w_002_360);
  and2 I009_621(w_009_621, w_007_405, w_003_049);
  not1 I009_623(w_009_623, w_006_212);
  nand2 I009_625(w_009_625, w_001_001, w_007_259);
  not1 I009_626(w_009_626, w_000_082);
  nand2 I009_627(w_009_627, w_002_243, w_007_316);
  and2 I009_628(w_009_628, w_002_296, w_007_244);
  nand2 I009_629(w_009_629, w_000_674, w_008_169);
  not1 I009_630(w_009_632, w_009_631);
  not1 I009_631(w_009_633, w_009_632);
  not1 I009_632(w_009_634, w_009_633);
  not1 I009_633(w_009_635, w_009_634);
  nand2 I009_634(w_009_636, w_008_168, w_009_635);
  or2  I009_635(w_009_637, w_009_636, w_009_654);
  and2 I009_636(w_009_638, w_004_351, w_009_637);
  not1 I009_637(w_009_631, w_009_638);
  nand2 I009_638(w_009_643, w_009_642, w_008_022);
  not1 I009_639(w_009_644, w_009_643);
  nand2 I009_640(w_009_645, w_009_644, w_003_046);
  or2  I009_641(w_009_646, w_002_282, w_009_645);
  nand2 I009_642(w_009_647, w_009_646, w_002_014);
  nand2 I009_643(w_009_648, w_003_066, w_009_647);
  or2  I009_644(w_009_649, w_009_648, w_003_025);
  or2  I009_645(w_009_650, w_009_649, w_002_518);
  nand2 I009_646(w_009_651, w_009_650, w_004_041);
  and2 I009_647(w_009_652, w_002_363, w_009_651);
  not1 I009_648(w_009_642, w_009_637);
  and2 I009_649(w_009_654, w_005_299, w_009_652);
  not1 I010_000(w_010_000, w_005_176);
  and2 I010_002(w_010_002, w_004_267, w_007_300);
  and2 I010_003(w_010_003, w_002_082, w_008_125);
  and2 I010_004(w_010_004, w_005_169, w_005_054);
  not1 I010_005(w_010_005, w_001_028);
  and2 I010_006(w_010_006, w_007_003, w_006_009);
  and2 I010_008(w_010_008, w_008_679, w_000_172);
  and2 I010_009(w_010_009, w_008_506, w_009_522);
  and2 I010_010(w_010_010, w_007_165, w_004_454);
  or2  I010_011(w_010_011, w_009_028, w_009_172);
  or2  I010_012(w_010_012, w_006_229, w_004_274);
  and2 I010_013(w_010_013, w_007_285, w_009_138);
  not1 I010_014(w_010_014, w_003_076);
  not1 I010_016(w_010_016, w_003_052);
  nand2 I010_017(w_010_017, w_005_061, w_001_010);
  and2 I010_018(w_010_018, w_007_282, w_005_097);
  not1 I010_020(w_010_020, w_005_257);
  nand2 I010_021(w_010_021, w_005_187, w_008_089);
  and2 I010_027(w_010_027, w_004_022, w_006_091);
  and2 I010_031(w_010_031, w_008_248, w_005_005);
  or2  I010_032(w_010_032, w_002_420, w_001_006);
  or2  I010_036(w_010_036, w_009_104, w_006_175);
  nand2 I010_039(w_010_039, w_003_061, w_002_093);
  not1 I010_042(w_010_042, w_003_017);
  nand2 I010_043(w_010_043, w_006_030, w_007_010);
  not1 I010_045(w_010_045, w_000_479);
  not1 I010_049(w_010_049, w_003_027);
  nand2 I010_050(w_010_050, w_002_084, w_007_286);
  or2  I010_051(w_010_051, w_009_501, w_007_049);
  or2  I010_053(w_010_053, w_002_557, w_000_022);
  nand2 I010_054(w_010_054, w_003_078, w_002_113);
  or2  I010_056(w_010_056, w_004_231, w_001_013);
  nand2 I010_057(w_010_057, w_004_085, w_002_151);
  or2  I010_058(w_010_058, w_007_094, w_008_434);
  and2 I010_059(w_010_059, w_009_326, w_009_572);
  and2 I010_060(w_010_060, w_002_017, w_008_646);
  not1 I010_061(w_010_061, w_005_161);
  and2 I010_064(w_010_064, w_009_107, w_006_136);
  nand2 I010_067(w_010_067, w_006_111, w_005_204);
  or2  I010_070(w_010_070, w_002_359, w_001_025);
  not1 I010_073(w_010_073, w_008_110);
  and2 I010_074(w_010_074, w_006_148, w_002_373);
  and2 I010_076(w_010_076, w_004_237, w_006_097);
  not1 I010_077(w_010_077, w_005_114);
  not1 I010_078(w_010_078, w_004_017);
  nand2 I010_080(w_010_080, w_007_039, w_006_003);
  and2 I010_083(w_010_083, w_000_389, w_008_677);
  and2 I010_084(w_010_084, w_004_343, w_004_140);
  not1 I010_085(w_010_085, w_008_135);
  nand2 I010_086(w_010_086, w_009_451, w_008_298);
  not1 I010_087(w_010_087, w_004_007);
  not1 I010_088(w_010_088, w_008_371);
  and2 I010_089(w_010_089, w_008_396, w_003_066);
  or2  I010_091(w_010_091, w_000_135, w_005_185);
  or2  I010_094(w_010_094, w_004_151, w_007_187);
  not1 I010_095(w_010_095, w_006_024);
  and2 I010_097(w_010_097, w_005_257, w_004_196);
  and2 I010_099(w_010_099, w_001_008, w_009_403);
  or2  I010_102(w_010_102, w_007_222, w_000_680);
  not1 I010_105(w_010_105, w_004_271);
  not1 I010_106(w_010_106, w_006_038);
  and2 I010_107(w_010_107, w_001_036, w_007_045);
  nand2 I010_108(w_010_108, w_000_281, w_000_456);
  nand2 I010_109(w_010_109, w_007_230, w_005_014);
  or2  I010_113(w_010_113, w_000_521, w_005_125);
  nand2 I010_114(w_010_114, w_002_171, w_008_284);
  nand2 I010_117(w_010_117, w_002_274, w_003_005);
  not1 I010_118(w_010_118, w_001_000);
  or2  I010_119(w_010_119, w_005_042, w_008_528);
  not1 I010_120(w_010_120, w_005_172);
  or2  I010_121(w_010_121, w_007_343, w_009_522);
  nand2 I010_122(w_010_122, w_000_014, w_009_368);
  nand2 I010_123(w_010_123, w_007_382, w_002_400);
  or2  I010_124(w_010_124, w_004_227, w_004_064);
  or2  I010_125(w_010_125, w_007_320, w_008_733);
  and2 I010_126(w_010_126, w_006_208, w_002_383);
  or2  I010_127(w_010_127, w_003_026, w_000_455);
  nand2 I010_128(w_010_128, w_009_375, w_001_018);
  nand2 I010_129(w_010_129, w_000_548, w_007_384);
  and2 I010_130(w_010_130, w_008_189, w_007_373);
  or2  I010_131(w_010_131, w_005_000, w_005_003);
  nand2 I010_133(w_010_133, w_003_006, w_008_563);
  nand2 I010_134(w_010_134, w_005_224, w_006_063);
  or2  I010_135(w_010_135, w_003_006, w_003_027);
  not1 I010_136(w_010_136, w_004_480);
  nand2 I010_139(w_010_139, w_004_406, w_000_216);
  or2  I010_140(w_010_140, w_003_052, w_004_279);
  or2  I010_144(w_010_144, w_000_681, w_005_169);
  and2 I010_145(w_010_145, w_003_028, w_002_119);
  and2 I010_147(w_010_147, w_000_656, w_008_194);
  and2 I010_148(w_010_148, w_001_028, w_000_680);
  and2 I010_149(w_010_149, w_005_229, w_008_682);
  or2  I010_151(w_010_151, w_006_230, w_006_062);
  not1 I010_154(w_010_154, w_006_076);
  nand2 I010_155(w_010_155, w_000_682, w_003_030);
  nand2 I010_156(w_010_156, w_000_010, w_000_412);
  and2 I010_157(w_010_157, w_005_078, w_008_478);
  not1 I010_158(w_010_158, w_004_415);
  not1 I010_159(w_010_159, w_005_023);
  nand2 I010_161(w_010_161, w_002_692, w_006_194);
  nand2 I010_162(w_010_162, w_008_758, w_000_380);
  or2  I010_163(w_010_163, w_000_390, w_009_594);
  not1 I010_164(w_010_164, w_005_062);
  not1 I010_165(w_010_165, w_003_004);
  nand2 I010_166(w_010_166, w_000_243, w_002_673);
  and2 I010_168(w_010_168, w_001_018, w_000_250);
  and2 I010_169(w_010_169, w_008_208, w_004_268);
  or2  I010_172(w_010_172, w_008_029, w_004_360);
  or2  I010_174(w_010_174, w_002_066, w_004_279);
  and2 I010_177(w_010_177, w_006_015, w_000_444);
  and2 I010_178(w_010_178, w_003_077, w_008_078);
  and2 I010_179(w_010_179, w_000_675, w_006_024);
  and2 I010_181(w_010_181, w_004_113, w_000_683);
  and2 I010_183(w_010_183, w_008_281, w_005_024);
  nand2 I010_185(w_010_185, w_009_138, w_003_042);
  and2 I010_186(w_010_186, w_000_319, w_008_729);
  nand2 I010_187(w_010_187, w_000_222, w_007_385);
  or2  I010_188(w_010_188, w_008_378, w_003_013);
  nand2 I010_190(w_010_190, w_001_017, w_003_015);
  nand2 I010_191(w_010_191, w_004_331, w_000_114);
  nand2 I010_192(w_010_192, w_004_156, w_007_256);
  nand2 I010_193(w_010_193, w_005_185, w_008_056);
  nand2 I010_194(w_010_194, w_006_034, w_004_326);
  and2 I010_196(w_010_196, w_009_097, w_006_224);
  or2  I010_197(w_010_197, w_002_578, w_000_152);
  not1 I010_199(w_010_199, w_008_347);
  and2 I010_201(w_010_201, w_003_052, w_001_017);
  and2 I010_204(w_010_204, w_008_173, w_003_037);
  and2 I010_205(w_010_205, w_003_028, w_008_301);
  and2 I010_207(w_010_207, w_007_237, w_009_019);
  or2  I010_209(w_010_209, w_002_022, w_007_209);
  and2 I010_210(w_010_210, w_003_032, w_006_113);
  or2  I010_211(w_010_211, w_009_235, w_001_023);
  and2 I010_213(w_010_213, w_008_726, w_003_043);
  or2  I010_216(w_010_216, w_009_106, w_009_014);
  not1 I010_217(w_010_217, w_007_127);
  and2 I010_218(w_010_218, w_007_362, w_009_194);
  nand2 I010_219(w_010_219, w_009_032, w_004_219);
  nand2 I010_220(w_010_220, w_004_146, w_004_252);
  and2 I010_221(w_010_221, w_008_291, w_006_185);
  not1 I010_222(w_010_222, w_008_107);
  and2 I010_224(w_010_224, w_008_164, w_002_457);
  not1 I010_225(w_010_225, w_001_022);
  or2  I010_226(w_010_226, w_003_065, w_005_023);
  and2 I010_227(w_010_227, w_000_040, w_000_522);
  and2 I010_228(w_010_228, w_000_366, w_005_074);
  and2 I010_229(w_010_229, w_003_031, w_006_179);
  and2 I010_230(w_010_230, w_008_370, w_008_698);
  and2 I010_232(w_010_232, w_004_048, w_006_183);
  and2 I010_233(w_010_233, w_001_028, w_000_684);
  not1 I010_235(w_010_235, w_007_007);
  not1 I010_236(w_010_236, w_003_060);
  nand2 I010_238(w_010_238, w_000_565, w_003_081);
  and2 I010_240(w_010_240, w_001_010, w_003_072);
  and2 I010_241(w_010_241, w_008_348, w_006_186);
  or2  I010_242(w_010_242, w_004_357, w_008_088);
  not1 I010_243(w_010_243, w_000_578);
  and2 I010_245(w_010_245, w_004_395, w_007_453);
  or2  I010_248(w_010_248, w_003_079, w_004_037);
  and2 I010_249(w_010_249, w_005_158, w_004_445);
  and2 I010_250(w_010_250, w_006_019, w_003_048);
  nand2 I010_255(w_010_255, w_003_033, w_008_518);
  not1 I010_258(w_010_258, w_003_007);
  not1 I010_259(w_010_259, w_000_685);
  or2  I010_260(w_010_260, w_008_629, w_000_142);
  or2  I010_261(w_010_261, w_008_004, w_005_030);
  or2  I010_263(w_010_263, w_009_361, w_003_055);
  or2  I010_264(w_010_264, w_009_066, w_001_019);
  nand2 I010_265(w_010_265, w_001_027, w_004_470);
  and2 I010_268(w_010_268, w_006_223, w_004_142);
  or2  I010_269(w_010_269, w_000_252, w_004_443);
  and2 I010_270(w_010_270, w_004_215, w_000_295);
  and2 I010_272(w_010_272, w_005_292, w_004_091);
  not1 I010_275(w_010_275, w_004_441);
  nand2 I010_276(w_010_276, w_004_245, w_006_161);
  or2  I010_277(w_010_277, w_000_082, w_001_006);
  or2  I010_278(w_010_278, w_004_257, w_003_026);
  or2  I010_280(w_010_280, w_001_014, w_006_207);
  and2 I010_282(w_010_282, w_007_204, w_004_253);
  or2  I010_283(w_010_283, w_002_631, w_000_352);
  not1 I010_285(w_010_285, w_008_718);
  nand2 I010_286(w_010_286, w_008_472, w_001_006);
  not1 I010_288(w_010_288, w_001_016);
  not1 I010_289(w_010_289, w_008_013);
  not1 I010_290(w_010_290, w_002_014);
  and2 I010_291(w_010_291, w_005_238, w_000_602);
  not1 I010_295(w_010_295, w_006_054);
  and2 I010_298(w_010_298, w_002_180, w_002_695);
  or2  I010_300(w_010_300, w_005_150, w_004_140);
  nand2 I010_301(w_010_301, w_007_172, w_009_075);
  or2  I010_303(w_010_303, w_007_147, w_009_166);
  not1 I010_306(w_010_306, w_000_441);
  or2  I010_308(w_010_308, w_000_491, w_008_011);
  nand2 I010_311(w_010_311, w_009_196, w_009_376);
  nand2 I010_312(w_010_312, w_006_096, w_005_312);
  and2 I010_313(w_010_313, w_005_305, w_009_122);
  not1 I010_314(w_010_314, w_002_311);
  nand2 I010_315(w_010_315, w_004_354, w_003_068);
  nand2 I010_317(w_010_317, w_002_526, w_002_563);
  or2  I010_319(w_010_319, w_001_001, w_003_081);
  or2  I010_321(w_010_321, w_004_151, w_004_098);
  and2 I010_322(w_010_322, w_008_024, w_008_517);
  nand2 I010_326(w_010_326, w_000_053, w_007_068);
  and2 I010_327(w_010_327, w_001_031, w_001_014);
  and2 I010_328(w_010_328, w_005_248, w_000_135);
  nand2 I010_331(w_010_331, w_002_362, w_001_010);
  or2  I010_335(w_010_335, w_000_092, w_006_014);
  or2  I010_338(w_010_338, w_002_202, w_002_565);
  and2 I010_339(w_010_339, w_009_300, w_009_444);
  not1 I010_341(w_010_341, w_003_065);
  not1 I010_342(w_010_342, w_005_189);
  not1 I010_343(w_010_343, w_007_294);
  or2  I010_347(w_010_347, w_008_329, w_003_046);
  nand2 I010_348(w_010_348, w_007_039, w_007_205);
  not1 I010_349(w_010_349, w_004_255);
  nand2 I010_350(w_010_350, w_003_028, w_001_030);
  nand2 I010_351(w_010_351, w_004_005, w_002_286);
  or2  I010_352(w_010_352, w_001_004, w_004_175);
  and2 I010_353(w_010_353, w_002_533, w_007_222);
  not1 I010_354(w_010_354, w_002_161);
  or2  I010_355(w_010_355, w_009_234, w_000_459);
  and2 I010_356(w_010_356, w_005_105, w_004_150);
  and2 I010_357(w_010_357, w_005_200, w_003_021);
  nand2 I010_358(w_010_358, w_007_308, w_000_138);
  not1 I010_359(w_010_359, w_006_061);
  not1 I010_360(w_010_360, w_000_399);
  nand2 I010_361(w_010_361, w_003_014, w_001_016);
  nand2 I010_362(w_010_362, w_003_025, w_008_552);
  and2 I010_364(w_010_364, w_001_007, w_003_068);
  nand2 I010_365(w_010_365, w_002_523, w_004_311);
  and2 I010_368(w_010_368, w_000_064, w_004_078);
  and2 I010_369(w_010_369, w_004_253, w_009_581);
  not1 I010_370(w_010_370, w_007_292);
  not1 I010_373(w_010_373, w_008_069);
  not1 I010_375(w_010_375, w_007_266);
  not1 I010_377(w_010_377, w_005_058);
  and2 I010_381(w_010_381, w_001_006, w_002_427);
  not1 I010_382(w_010_382, w_008_474);
  or2  I010_383(w_010_383, w_008_140, w_007_279);
  not1 I010_384(w_010_384, w_004_337);
  or2  I010_385(w_010_385, w_006_201, w_009_011);
  not1 I010_386(w_010_386, w_007_019);
  not1 I010_387(w_010_387, w_009_550);
  and2 I010_388(w_010_388, w_005_063, w_006_089);
  not1 I010_395(w_010_395, w_007_175);
  nand2 I010_396(w_010_396, w_000_124, w_009_245);
  or2  I010_397(w_010_397, w_005_033, w_004_201);
  nand2 I010_398(w_010_398, w_004_066, w_009_144);
  or2  I010_399(w_010_399, w_009_460, w_002_201);
  not1 I010_400(w_010_400, w_006_197);
  or2  I010_403(w_010_403, w_001_006, w_006_153);
  and2 I010_405(w_010_405, w_005_171, w_007_419);
  or2  I010_406(w_010_406, w_008_431, w_005_311);
  or2  I010_407(w_010_407, w_004_085, w_000_309);
  and2 I010_408(w_010_408, w_003_053, w_008_054);
  or2  I010_412(w_010_412, w_003_009, w_000_039);
  nand2 I010_413(w_010_413, w_003_000, w_004_265);
  and2 I010_414(w_010_414, w_007_179, w_009_135);
  nand2 I010_415(w_010_415, w_003_072, w_002_041);
  nand2 I010_416(w_010_416, w_005_080, w_009_209);
  nand2 I010_417(w_010_417, w_008_011, w_001_027);
  and2 I010_418(w_010_418, w_002_146, w_001_005);
  or2  I010_419(w_010_419, w_001_016, w_002_037);
  or2  I010_420(w_010_420, w_006_081, w_006_244);
  or2  I010_421(w_010_421, w_003_020, w_005_236);
  nand2 I010_423(w_010_423, w_009_098, w_002_082);
  and2 I010_425(w_010_425, w_005_019, w_001_011);
  or2  I010_426(w_010_426, w_003_001, w_002_061);
  and2 I010_427(w_010_427, w_008_558, w_006_193);
  or2  I010_428(w_010_428, w_001_008, w_007_092);
  not1 I010_429(w_010_429, w_003_020);
  nand2 I010_431(w_010_431, w_001_003, w_003_012);
  and2 I010_432(w_010_432, w_007_003, w_005_011);
  not1 I010_434(w_010_434, w_006_088);
  or2  I010_437(w_010_437, w_008_237, w_000_687);
  or2  I010_441(w_010_441, w_005_139, w_009_075);
  not1 I010_442(w_010_442, w_003_057);
  nand2 I010_443(w_010_443, w_003_036, w_001_036);
  and2 I010_444(w_010_444, w_009_144, w_004_271);
  or2  I010_446(w_010_446, w_006_171, w_009_283);
  not1 I010_447(w_010_447, w_000_628);
  not1 I010_449(w_010_449, w_004_024);
  or2  I010_450(w_010_450, w_007_365, w_004_162);
  not1 I010_451(w_010_451, w_006_198);
  not1 I010_452(w_010_452, w_009_371);
  not1 I010_453(w_010_453, w_000_688);
  nand2 I010_454(w_010_454, w_000_230, w_008_461);
  or2  I010_455(w_010_455, w_003_081, w_002_213);
  or2  I010_456(w_010_456, w_002_302, w_006_064);
  and2 I010_457(w_010_457, w_002_057, w_006_028);
  nand2 I010_458(w_010_458, w_000_238, w_009_098);
  and2 I010_459(w_010_459, w_008_469, w_003_001);
  not1 I010_460(w_010_460, w_008_001);
  not1 I010_466(w_010_466, w_002_312);
  or2  I010_467(w_010_467, w_005_259, w_003_031);
  nand2 I010_468(w_010_468, w_002_300, w_007_413);
  and2 I010_471(w_010_471, w_008_374, w_008_423);
  and2 I010_472(w_010_472, w_002_266, w_005_297);
  or2  I010_476(w_010_476, w_000_113, w_006_115);
  or2  I010_478(w_010_478, w_000_003, w_008_485);
  and2 I010_479(w_010_479, w_009_106, w_003_010);
  not1 I010_481(w_010_481, w_005_075);
  nand2 I010_482(w_010_482, w_005_246, w_001_000);
  or2  I010_484(w_010_484, w_000_689, w_007_156);
  not1 I010_486(w_010_486, w_006_010);
  or2  I010_487(w_010_487, w_004_089, w_007_408);
  nand2 I010_488(w_010_488, w_008_582, w_001_022);
  or2  I010_489(w_010_489, w_008_250, w_000_653);
  not1 I010_491(w_010_491, w_001_015);
  or2  I010_494(w_010_494, w_006_000, w_001_001);
  not1 I010_496(w_010_496, w_004_124);
  and2 I010_497(w_010_497, w_009_043, w_006_223);
  not1 I010_498(w_010_498, w_004_091);
  nand2 I010_499(w_010_499, w_006_041, w_003_069);
  and2 I010_500(w_010_500, w_000_053, w_008_724);
  nand2 I010_505(w_010_505, w_001_020, w_005_075);
  and2 I010_506(w_010_506, w_001_036, w_005_119);
  or2  I010_507(w_010_507, w_004_226, w_001_004);
  or2  I010_510(w_010_510, w_006_215, w_005_150);
  or2  I010_511(w_010_511, w_002_049, w_006_151);
  and2 I010_513(w_010_513, w_002_018, w_008_226);
  or2  I010_514(w_010_514, w_008_288, w_007_148);
  and2 I010_515(w_010_515, w_003_053, w_008_397);
  or2  I010_516(w_010_516, w_009_583, w_004_064);
  nand2 I010_517(w_010_517, w_009_237, w_003_033);
  not1 I010_518(w_010_518, w_009_236);
  nand2 I010_519(w_010_519, w_002_234, w_009_384);
  or2  I010_520(w_010_520, w_009_610, w_000_088);
  nand2 I010_522(w_010_522, w_001_023, w_008_541);
  not1 I010_525(w_010_525, w_002_424);
  and2 I010_526(w_010_526, w_003_021, w_001_002);
  nand2 I010_528(w_010_528, w_007_264, w_004_099);
  not1 I010_529(w_010_529, w_004_192);
  nand2 I010_530(w_010_530, w_008_411, w_003_013);
  and2 I010_531(w_010_531, w_007_295, w_001_018);
  or2  I010_532(w_010_532, w_003_051, w_001_002);
  or2  I010_533(w_010_533, w_003_060, w_000_690);
  or2  I010_539(w_010_539, w_001_000, w_003_034);
  not1 I010_540(w_010_540, w_004_321);
  or2  I010_542(w_010_542, w_004_452, w_008_271);
  not1 I010_544(w_010_544, w_006_227);
  not1 I010_548(w_010_548, w_005_074);
  and2 I010_550(w_010_550, w_004_282, w_003_038);
  and2 I010_551(w_010_551, w_006_156, w_000_198);
  and2 I010_553(w_010_553, w_008_227, w_006_016);
  or2  I010_554(w_010_554, w_001_033, w_003_016);
  nand2 I010_556(w_010_556, w_002_220, w_004_345);
  nand2 I010_558(w_010_558, w_008_710, w_004_087);
  or2  I010_559(w_010_559, w_009_508, w_007_347);
  nand2 I010_560(w_010_560, w_006_168, w_006_039);
  and2 I010_561(w_010_561, w_009_395, w_000_684);
  and2 I010_563(w_010_563, w_004_489, w_000_662);
  or2  I010_564(w_010_564, w_009_541, w_003_003);
  not1 I010_565(w_010_565, w_005_302);
  not1 I010_566(w_010_566, w_004_201);
  or2  I010_567(w_010_567, w_000_075, w_003_069);
  and2 I010_568(w_010_568, w_005_038, w_002_389);
  and2 I010_569(w_010_569, w_003_071, w_002_469);
  or2  I010_570(w_010_570, w_007_158, w_003_036);
  nand2 I010_571(w_010_571, w_003_044, w_004_148);
  not1 I010_576(w_010_576, w_004_049);
  nand2 I010_577(w_010_577, w_005_193, w_004_288);
  not1 I010_579(w_010_579, w_003_049);
  not1 I010_580(w_010_580, w_008_707);
  or2  I010_581(w_010_581, w_009_142, w_009_123);
  and2 I010_583(w_010_583, w_009_440, w_005_230);
  not1 I010_584(w_010_584, w_006_224);
  not1 I010_585(w_010_585, w_009_369);
  not1 I010_586(w_010_586, w_002_223);
  not1 I010_587(w_010_587, w_008_437);
  nand2 I010_588(w_010_588, w_008_577, w_003_027);
  and2 I010_589(w_010_589, w_007_161, w_002_426);
  not1 I010_591(w_010_591, w_003_026);
  nand2 I010_592(w_010_592, w_008_089, w_002_212);
  and2 I010_593(w_010_593, w_003_044, w_002_276);
  not1 I010_595(w_010_595, w_001_024);
  nand2 I010_596(w_010_596, w_001_015, w_003_032);
  or2  I010_597(w_010_597, w_009_557, w_000_353);
  nand2 I010_598(w_010_598, w_006_103, w_003_009);
  or2  I010_599(w_010_599, w_007_198, w_005_074);
  and2 I010_603(w_010_603, w_004_486, w_007_011);
  nand2 I010_604(w_010_604, w_000_398, w_000_466);
  nand2 I010_606(w_010_606, w_002_650, w_009_456);
  nand2 I010_609(w_010_609, w_001_009, w_003_065);
  and2 I010_610(w_010_610, w_007_346, w_001_024);
  or2  I010_611(w_010_611, w_003_034, w_009_041);
  not1 I010_612(w_010_612, w_005_174);
  or2  I010_613(w_010_613, w_009_065, w_008_386);
  not1 I010_614(w_010_614, w_009_583);
  and2 I010_616(w_010_616, w_008_589, w_005_003);
  nand2 I010_618(w_010_618, w_003_062, w_004_332);
  not1 I010_619(w_010_619, w_006_144);
  not1 I010_622(w_010_622, w_003_042);
  or2  I010_623(w_010_623, w_001_006, w_005_013);
  or2  I010_625(w_010_625, w_001_036, w_002_616);
  nand2 I010_626(w_010_626, w_007_410, w_007_477);
  or2  I010_627(w_010_627, w_009_597, w_005_114);
  and2 I010_628(w_010_628, w_008_133, w_000_093);
  nand2 I010_631(w_010_631, w_003_060, w_005_018);
  or2  I010_632(w_010_632, w_009_153, w_007_426);
  nand2 I010_633(w_010_633, w_006_104, w_008_505);
  and2 I010_635(w_010_635, w_003_039, w_006_057);
  or2  I010_638(w_010_638, w_007_010, w_004_106);
  and2 I010_640(w_010_640, w_006_101, w_001_004);
  and2 I010_641(w_010_641, w_008_383, w_001_030);
  or2  I010_642(w_010_642, w_007_106, w_002_353);
  or2  I010_644(w_010_644, w_007_353, w_009_153);
  nand2 I010_645(w_010_645, w_008_735, w_006_054);
  and2 I010_646(w_010_646, w_006_106, w_003_034);
  and2 I010_649(w_010_649, w_008_664, w_005_001);
  not1 I010_653(w_010_653, w_005_063);
  not1 I010_655(w_010_655, w_006_082);
  or2  I010_656(w_010_656, w_000_481, w_002_366);
  not1 I010_659(w_010_659, w_006_062);
  not1 I010_660(w_010_660, w_004_384);
  nand2 I010_661(w_010_661, w_000_691, w_005_012);
  and2 I010_663(w_010_663, w_006_004, w_008_582);
  and2 I010_667(w_010_667, w_001_024, w_009_374);
  or2  I010_668(w_010_668, w_004_228, w_005_025);
  or2  I010_669(w_010_669, w_001_001, w_009_427);
  not1 I010_670(w_010_670, w_009_561);
  or2  I010_672(w_010_672, w_005_309, w_004_199);
  not1 I010_673(w_010_673, w_000_561);
  not1 I010_674(w_010_674, w_001_026);
  or2  I010_675(w_010_675, w_005_085, w_006_021);
  or2  I010_677(w_010_677, w_009_480, w_003_039);
  or2  I010_678(w_010_678, w_004_136, w_000_281);
  not1 I010_679(w_010_679, w_005_068);
  and2 I010_680(w_010_680, w_006_206, w_009_158);
  not1 I010_681(w_010_681, w_000_438);
  and2 I010_682(w_010_682, w_009_359, w_001_005);
  nand2 I010_684(w_010_684, w_007_416, w_002_158);
  not1 I010_685(w_010_685, w_009_005);
  not1 I010_686(w_010_686, w_002_139);
  nand2 I010_688(w_010_688, w_002_165, w_001_022);
  and2 I010_691(w_010_691, w_007_191, w_007_273);
  or2  I010_692(w_010_692, w_006_001, w_003_078);
  nand2 I010_695(w_010_695, w_000_109, w_007_387);
  nand2 I010_697(w_010_697, w_003_024, w_008_382);
  and2 I010_698(w_010_698, w_009_100, w_002_135);
  and2 I010_700(w_010_700, w_006_151, w_001_036);
  or2  I010_703(w_010_703, w_002_291, w_000_488);
  or2  I010_705(w_010_705, w_008_657, w_001_035);
  nand2 I010_707(w_010_707, w_003_082, w_008_714);
  and2 I010_709(w_010_709, w_007_441, w_008_550);
  nand2 I010_711(w_010_711, w_005_113, w_003_041);
  or2  I010_712(w_010_712, w_007_278, w_000_317);
  or2  I010_713(w_010_713, w_002_092, w_005_282);
  nand2 I010_714(w_010_714, w_005_287, w_009_130);
  not1 I010_715(w_010_715, w_006_127);
  and2 I010_716(w_010_716, w_004_229, w_009_150);
  not1 I010_717(w_010_717, w_001_003);
  not1 I010_718(w_010_718, w_006_011);
  nand2 I010_719(w_010_719, w_005_302, w_008_727);
  and2 I010_720(w_010_720, w_007_303, w_006_235);
  not1 I010_721(w_010_721, w_008_748);
  nand2 I010_722(w_010_722, w_008_680, w_009_394);
  and2 I010_724(w_010_724, w_000_693, w_009_364);
  not1 I010_726(w_010_726, w_008_702);
  nand2 I010_731(w_010_731, w_000_221, w_008_748);
  or2  I010_732(w_010_732, w_006_217, w_004_224);
  not1 I010_733(w_010_733, w_009_521);
  not1 I010_735(w_010_735, w_008_076);
  nand2 I010_736(w_010_736, w_000_645, w_008_490);
  and2 I010_737(w_010_737, w_005_149, w_009_542);
  or2  I010_739(w_010_739, w_005_123, w_003_036);
  nand2 I010_742(w_010_742, w_009_156, w_004_220);
  not1 I010_743(w_010_743, w_004_105);
  or2  I010_745(w_010_745, w_007_067, w_004_137);
  and2 I010_746(w_010_746, w_009_140, w_001_017);
  and2 I010_747(w_010_747, w_005_064, w_009_022);
  and2 I010_748(w_010_748, w_005_218, w_000_231);
  and2 I010_749(w_010_749, w_001_017, w_003_026);
  not1 I010_750(w_010_750, w_009_217);
  and2 I010_751(w_010_751, w_005_098, w_000_044);
  or2  I010_753(w_010_753, w_004_426, w_003_025);
  or2  I010_754(w_010_754, w_004_144, w_005_149);
  and2 I010_756(w_010_756, w_004_172, w_008_534);
  or2  I010_757(w_010_757, w_004_131, w_000_196);
  nand2 I010_758(w_010_758, w_006_047, w_006_165);
  or2  I010_759(w_010_759, w_009_486, w_007_283);
  not1 I010_760(w_010_760, w_008_289);
  nand2 I010_763(w_010_763, w_005_005, w_000_620);
  or2  I010_765(w_010_765, w_001_030, w_008_112);
  not1 I010_766(w_010_766, w_008_077);
  and2 I010_767(w_010_767, w_006_114, w_002_224);
  not1 I010_768(w_010_768, w_009_018);
  or2  I010_769(w_010_769, w_005_035, w_009_078);
  and2 I010_770(w_010_770, w_004_265, w_002_054);
  or2  I010_773(w_010_773, w_001_010, w_009_499);
  and2 I010_775(w_010_775, w_000_694, w_002_597);
  nand2 I010_777(w_010_777, w_000_572, w_005_195);
  or2  I010_779(w_010_779, w_002_657, w_004_273);
  and2 I011_001(w_011_001, w_001_017, w_010_226);
  nand2 I011_002(w_011_002, w_008_350, w_007_171);
  or2  I011_003(w_011_003, w_004_449, w_006_022);
  not1 I011_004(w_011_004, w_010_737);
  and2 I011_005(w_011_005, w_010_005, w_008_137);
  or2  I011_006(w_011_006, w_002_096, w_006_227);
  and2 I011_007(w_011_007, w_006_107, w_001_033);
  not1 I011_009(w_011_009, w_006_037);
  nand2 I011_010(w_011_010, w_000_695, w_007_373);
  and2 I011_011(w_011_011, w_004_311, w_009_015);
  nand2 I011_013(w_011_013, w_000_395, w_003_069);
  and2 I011_014(w_011_014, w_005_072, w_005_021);
  nand2 I011_015(w_011_015, w_004_165, w_002_644);
  not1 I011_016(w_011_016, w_000_489);
  and2 I011_017(w_011_017, w_007_414, w_010_088);
  or2  I011_018(w_011_018, w_006_228, w_001_014);
  or2  I011_020(w_011_020, w_002_667, w_006_019);
  not1 I011_021(w_011_021, w_009_360);
  not1 I011_022(w_011_022, w_000_525);
  and2 I011_023(w_011_023, w_009_239, w_009_128);
  nand2 I011_024(w_011_024, w_004_095, w_008_479);
  and2 I011_025(w_011_025, w_003_073, w_009_531);
  not1 I011_026(w_011_026, w_002_001);
  not1 I011_027(w_011_027, w_009_395);
  not1 I011_028(w_011_028, w_010_285);
  nand2 I011_030(w_011_030, w_007_136, w_007_228);
  and2 I011_031(w_011_031, w_001_033, w_006_202);
  not1 I011_032(w_011_032, w_008_575);
  nand2 I011_033(w_011_033, w_000_274, w_007_004);
  nand2 I011_035(w_011_035, w_010_136, w_007_060);
  and2 I011_036(w_011_036, w_008_237, w_009_007);
  nand2 I011_037(w_011_037, w_003_037, w_010_306);
  and2 I011_039(w_011_039, w_009_169, w_006_149);
  not1 I011_041(w_011_041, w_010_169);
  not1 I011_042(w_011_042, w_005_074);
  nand2 I011_043(w_011_043, w_002_501, w_008_247);
  and2 I011_044(w_011_044, w_000_696, w_009_260);
  and2 I011_045(w_011_045, w_001_007, w_007_245);
  or2  I011_046(w_011_046, w_005_129, w_002_016);
  and2 I011_047(w_011_047, w_010_139, w_009_354);
  or2  I011_048(w_011_048, w_007_042, w_005_185);
  and2 I011_049(w_011_049, w_004_114, w_003_075);
  or2  I011_050(w_011_050, w_001_021, w_001_029);
  and2 I011_051(w_011_051, w_003_018, w_002_579);
  nand2 I011_052(w_011_052, w_010_105, w_003_022);
  or2  I011_054(w_011_054, w_010_452, w_001_036);
  not1 I011_056(w_011_056, w_004_045);
  nand2 I011_057(w_011_057, w_005_266, w_009_532);
  or2  I011_058(w_011_058, w_010_720, w_010_517);
  nand2 I011_059(w_011_059, w_007_141, w_004_468);
  or2  I011_060(w_011_060, w_007_083, w_010_748);
  or2  I011_061(w_011_061, w_000_128, w_005_218);
  or2  I011_062(w_011_062, w_006_038, w_001_033);
  nand2 I011_063(w_011_063, w_009_221, w_001_020);
  or2  I011_064(w_011_064, w_009_032, w_006_135);
  or2  I011_066(w_011_066, w_003_029, w_007_407);
  or2  I011_069(w_011_069, w_009_271, w_010_421);
  not1 I011_070(w_011_070, w_006_194);
  not1 I011_071(w_011_071, w_009_499);
  nand2 I011_072(w_011_072, w_001_017, w_005_116);
  or2  I011_073(w_011_073, w_006_140, w_006_008);
  nand2 I011_075(w_011_075, w_005_053, w_006_060);
  or2  I011_077(w_011_077, w_009_391, w_004_350);
  nand2 I011_078(w_011_078, w_005_078, w_001_033);
  and2 I011_079(w_011_079, w_004_214, w_000_381);
  or2  I011_080(w_011_080, w_006_205, w_007_459);
  not1 I011_081(w_011_081, w_009_246);
  not1 I011_082(w_011_082, w_002_659);
  nand2 I011_083(w_011_083, w_005_094, w_008_496);
  and2 I011_084(w_011_084, w_004_439, w_008_196);
  not1 I011_085(w_011_085, w_003_027);
  not1 I011_086(w_011_086, w_001_016);
  not1 I011_087(w_011_087, w_003_026);
  and2 I011_088(w_011_088, w_005_083, w_004_376);
  not1 I011_089(w_011_089, w_009_079);
  or2  I011_090(w_011_090, w_010_155, w_002_109);
  not1 I011_092(w_011_092, w_003_072);
  or2  I011_093(w_011_093, w_001_005, w_008_760);
  nand2 I011_094(w_011_094, w_007_255, w_003_055);
  not1 I011_095(w_011_095, w_009_158);
  nand2 I011_096(w_011_096, w_008_646, w_003_015);
  not1 I011_097(w_011_097, w_010_685);
  and2 I011_098(w_011_098, w_004_279, w_004_094);
  and2 I011_099(w_011_099, w_005_020, w_002_026);
  not1 I011_102(w_011_102, w_010_386);
  or2  I011_103(w_011_103, w_007_233, w_001_001);
  nand2 I011_104(w_011_104, w_009_220, w_008_009);
  and2 I011_108(w_011_108, w_001_025, w_008_677);
  and2 I011_109(w_011_109, w_006_065, w_008_700);
  or2  I011_110(w_011_110, w_006_210, w_006_213);
  or2  I011_111(w_011_111, w_005_056, w_008_388);
  nand2 I011_112(w_011_112, w_004_024, w_006_141);
  or2  I011_113(w_011_113, w_009_547, w_000_113);
  nand2 I011_114(w_011_114, w_005_156, w_007_035);
  and2 I011_116(w_011_116, w_009_552, w_007_233);
  or2  I011_117(w_011_117, w_001_006, w_000_331);
  and2 I011_118(w_011_118, w_005_097, w_004_024);
  not1 I011_119(w_011_119, w_001_027);
  not1 I011_120(w_011_120, w_010_006);
  or2  I011_121(w_011_121, w_004_352, w_009_279);
  and2 I011_123(w_011_123, w_005_254, w_009_080);
  not1 I011_124(w_011_124, w_008_134);
  not1 I011_125(w_011_125, w_007_264);
  or2  I011_126(w_011_126, w_007_101, w_010_513);
  or2  I011_127(w_011_127, w_002_403, w_004_172);
  and2 I011_128(w_011_128, w_007_104, w_004_009);
  nand2 I011_130(w_011_130, w_010_236, w_009_442);
  and2 I011_131(w_011_131, w_004_084, w_009_012);
  nand2 I011_132(w_011_132, w_005_121, w_008_015);
  not1 I011_133(w_011_133, w_005_046);
  and2 I011_134(w_011_134, w_008_001, w_000_697);
  not1 I011_135(w_011_135, w_007_092);
  or2  I011_136(w_011_136, w_007_040, w_000_596);
  and2 I011_137(w_011_137, w_008_032, w_004_019);
  or2  I011_138(w_011_138, w_007_165, w_009_191);
  and2 I011_139(w_011_139, w_001_021, w_001_025);
  or2  I011_140(w_011_140, w_006_140, w_009_155);
  nand2 I011_141(w_011_141, w_009_325, w_002_264);
  and2 I011_142(w_011_142, w_005_309, w_009_341);
  or2  I011_143(w_011_143, w_004_270, w_008_325);
  or2  I011_144(w_011_144, w_008_504, w_009_040);
  nand2 I011_146(w_011_146, w_005_019, w_008_656);
  or2  I011_147(w_011_147, w_009_146, w_000_278);
  not1 I011_148(w_011_148, w_006_148);
  nand2 I011_149(w_011_149, w_005_294, w_001_033);
  not1 I011_150(w_011_150, w_007_246);
  nand2 I011_151(w_011_151, w_002_072, w_006_246);
  and2 I011_152(w_011_152, w_008_088, w_010_585);
  or2  I011_154(w_011_154, w_002_443, w_004_160);
  not1 I011_155(w_011_155, w_010_114);
  or2  I011_156(w_011_156, w_002_048, w_006_207);
  nand2 I011_157(w_011_157, w_002_193, w_009_051);
  not1 I011_158(w_011_158, w_004_355);
  not1 I011_159(w_011_159, w_010_014);
  and2 I011_160(w_011_160, w_008_019, w_009_175);
  and2 I011_162(w_011_162, w_008_035, w_006_079);
  or2  I011_163(w_011_163, w_006_040, w_010_437);
  and2 I011_164(w_011_164, w_002_631, w_000_636);
  nand2 I011_166(w_011_166, w_005_051, w_006_063);
  not1 I011_167(w_011_167, w_001_006);
  not1 I011_168(w_011_168, w_000_283);
  nand2 I011_169(w_011_169, w_007_319, w_003_044);
  and2 I011_170(w_011_170, w_007_002, w_003_073);
  and2 I011_172(w_011_172, w_008_309, w_004_184);
  and2 I011_173(w_011_173, w_007_297, w_008_442);
  nand2 I011_174(w_011_174, w_009_296, w_005_278);
  nand2 I011_175(w_011_175, w_002_585, w_000_467);
  and2 I011_176(w_011_176, w_004_357, w_007_122);
  or2  I011_177(w_011_177, w_002_050, w_002_000);
  or2  I011_179(w_011_179, w_003_009, w_008_236);
  nand2 I011_180(w_011_180, w_010_777, w_007_254);
  nand2 I011_181(w_011_181, w_006_179, w_002_421);
  and2 I011_182(w_011_182, w_003_072, w_006_129);
  and2 I011_187(w_011_187, w_006_009, w_009_102);
  not1 I011_188(w_011_188, w_004_169);
  nand2 I011_189(w_011_189, w_008_073, w_010_384);
  not1 I011_190(w_011_190, w_007_362);
  or2  I011_191(w_011_191, w_006_138, w_008_697);
  nand2 I011_193(w_011_193, w_009_505, w_006_149);
  not1 I011_194(w_011_194, w_010_117);
  not1 I011_195(w_011_195, w_009_440);
  or2  I011_196(w_011_196, w_010_259, w_000_151);
  nand2 I011_197(w_011_197, w_007_004, w_000_432);
  nand2 I011_198(w_011_198, w_006_023, w_006_146);
  not1 I011_199(w_011_199, w_001_010);
  nand2 I011_201(w_011_201, w_008_381, w_001_000);
  not1 I011_202(w_011_202, w_004_171);
  and2 I011_203(w_011_203, w_002_320, w_001_011);
  not1 I011_204(w_011_204, w_000_361);
  and2 I011_205(w_011_205, w_002_482, w_003_012);
  and2 I011_206(w_011_206, w_004_106, w_007_246);
  nand2 I011_208(w_011_208, w_005_105, w_006_015);
  nand2 I011_209(w_011_209, w_010_011, w_004_283);
  and2 I011_210(w_011_210, w_006_197, w_002_328);
  not1 I011_211(w_011_211, w_003_064);
  nand2 I011_213(w_011_213, w_008_019, w_005_003);
  not1 I011_214(w_011_214, w_001_032);
  or2  I011_215(w_011_215, w_006_022, w_003_081);
  not1 I011_216(w_011_216, w_002_328);
  or2  I011_217(w_011_217, w_010_192, w_001_010);
  and2 I011_219(w_011_219, w_010_415, w_008_651);
  not1 I011_220(w_011_220, w_005_189);
  and2 I011_222(w_011_222, w_001_003, w_003_012);
  and2 I011_224(w_011_224, w_003_029, w_005_040);
  nand2 I011_227(w_011_227, w_007_043, w_004_361);
  not1 I011_228(w_011_228, w_003_061);
  not1 I011_229(w_011_229, w_008_049);
  or2  I011_231(w_011_231, w_010_129, w_009_168);
  and2 I011_232(w_011_232, w_001_026, w_000_368);
  not1 I011_233(w_011_233, w_010_224);
  not1 I011_235(w_011_235, w_003_007);
  nand2 I011_236(w_011_236, w_003_003, w_006_075);
  not1 I011_237(w_011_237, w_007_226);
  or2  I011_239(w_011_239, w_005_128, w_009_325);
  or2  I011_240(w_011_240, w_002_656, w_003_076);
  not1 I011_242(w_011_242, w_007_239);
  or2  I011_243(w_011_243, w_010_361, w_009_314);
  and2 I011_244(w_011_244, w_003_031, w_005_263);
  and2 I011_248(w_011_248, w_010_564, w_009_274);
  or2  I011_249(w_011_249, w_002_260, w_006_251);
  nand2 I011_251(w_011_251, w_009_029, w_003_057);
  nand2 I011_253(w_011_253, w_009_536, w_002_003);
  and2 I011_257(w_011_257, w_003_079, w_001_005);
  not1 I011_260(w_011_260, w_000_698);
  or2  I011_262(w_011_262, w_000_699, w_007_046);
  nand2 I011_263(w_011_263, w_005_084, w_008_461);
  and2 I011_265(w_011_265, w_006_059, w_004_292);
  not1 I011_267(w_011_267, w_010_446);
  or2  I011_268(w_011_268, w_001_001, w_000_626);
  not1 I011_269(w_011_269, w_007_225);
  or2  I011_270(w_011_270, w_000_181, w_007_235);
  and2 I011_271(w_011_271, w_004_263, w_006_184);
  nand2 I011_273(w_011_273, w_006_055, w_001_010);
  nand2 I011_276(w_011_276, w_009_482, w_001_011);
  not1 I011_278(w_011_278, w_010_285);
  or2  I011_279(w_011_279, w_003_049, w_002_551);
  nand2 I011_280(w_011_280, w_001_006, w_006_216);
  or2  I011_281(w_011_281, w_006_222, w_001_019);
  and2 I011_284(w_011_284, w_010_217, w_004_046);
  and2 I011_286(w_011_286, w_010_767, w_000_564);
  nand2 I011_288(w_011_288, w_010_414, w_008_615);
  not1 I011_289(w_011_289, w_006_098);
  or2  I011_290(w_011_290, w_002_063, w_008_108);
  or2  I011_291(w_011_291, w_000_664, w_002_365);
  or2  I011_295(w_011_295, w_009_168, w_010_377);
  not1 I011_298(w_011_298, w_005_154);
  or2  I011_300(w_011_300, w_007_227, w_010_487);
  and2 I011_301(w_011_301, w_003_002, w_001_023);
  not1 I011_302(w_011_302, w_008_669);
  not1 I011_303(w_011_303, w_010_317);
  not1 I011_306(w_011_306, w_010_530);
  and2 I011_308(w_011_308, w_006_241, w_009_628);
  or2  I011_309(w_011_309, w_004_503, w_010_165);
  or2  I011_310(w_011_310, w_007_035, w_009_258);
  or2  I011_312(w_011_312, w_001_022, w_009_016);
  nand2 I011_315(w_011_315, w_003_071, w_006_101);
  and2 I011_317(w_011_317, w_009_336, w_006_190);
  or2  I011_319(w_011_319, w_000_119, w_001_011);
  and2 I011_320(w_011_320, w_005_020, w_010_754);
  not1 I011_321(w_011_321, w_000_701);
  not1 I011_322(w_011_322, w_001_014);
  and2 I011_324(w_011_324, w_000_566, w_005_092);
  not1 I011_325(w_011_325, w_008_202);
  or2  I011_328(w_011_328, w_001_032, w_000_702);
  or2  I011_329(w_011_329, w_003_082, w_006_221);
  nand2 I011_330(w_011_330, w_005_092, w_001_033);
  or2  I011_332(w_011_332, w_003_031, w_001_027);
  or2  I011_333(w_011_333, w_004_199, w_004_200);
  or2  I011_334(w_011_334, w_004_297, w_003_031);
  or2  I011_336(w_011_336, w_005_043, w_006_084);
  nand2 I011_337(w_011_337, w_006_076, w_007_205);
  not1 I011_338(w_011_338, w_001_029);
  or2  I011_339(w_011_339, w_002_047, w_006_049);
  not1 I011_341(w_011_341, w_009_354);
  not1 I011_342(w_011_342, w_010_735);
  nand2 I011_343(w_011_343, w_004_108, w_007_206);
  or2  I011_344(w_011_344, w_006_246, w_001_006);
  and2 I011_345(w_011_345, w_004_197, w_003_082);
  or2  I011_347(w_011_347, w_010_432, w_001_026);
  nand2 I011_350(w_011_350, w_000_063, w_008_191);
  not1 I011_351(w_011_351, w_009_531);
  not1 I011_352(w_011_352, w_001_025);
  and2 I011_353(w_011_353, w_008_247, w_002_471);
  or2  I011_356(w_011_356, w_006_084, w_008_376);
  nand2 I011_357(w_011_357, w_008_439, w_009_047);
  not1 I011_359(w_011_359, w_010_382);
  or2  I011_360(w_011_360, w_010_054, w_001_005);
  not1 I011_361(w_011_361, w_004_482);
  not1 I011_364(w_011_364, w_000_430);
  not1 I011_365(w_011_365, w_000_535);
  not1 I011_366(w_011_366, w_002_643);
  nand2 I011_367(w_011_367, w_004_261, w_000_486);
  or2  I011_368(w_011_368, w_006_070, w_007_453);
  and2 I011_371(w_011_371, w_005_280, w_002_175);
  not1 I011_372(w_011_372, w_002_263);
  or2  I011_373(w_011_373, w_004_106, w_010_659);
  or2  I011_374(w_011_374, w_008_345, w_008_205);
  or2  I011_378(w_011_378, w_004_468, w_007_278);
  nand2 I011_379(w_011_379, w_007_309, w_007_193);
  or2  I011_383(w_011_383, w_003_045, w_008_594);
  and2 I011_384(w_011_384, w_007_163, w_005_108);
  or2  I011_385(w_011_385, w_008_696, w_008_036);
  nand2 I011_387(w_011_387, w_008_183, w_004_123);
  nand2 I011_390(w_011_390, w_001_016, w_007_178);
  and2 I011_391(w_011_391, w_009_126, w_005_098);
  and2 I011_392(w_011_392, w_009_344, w_006_023);
  and2 I011_393(w_011_393, w_000_193, w_007_451);
  or2  I011_396(w_011_396, w_009_040, w_010_507);
  or2  I011_397(w_011_397, w_005_304, w_004_322);
  and2 I011_398(w_011_398, w_010_656, w_009_408);
  not1 I011_401(w_011_401, w_000_106);
  and2 I011_405(w_011_405, w_006_078, w_003_027);
  not1 I011_406(w_011_406, w_010_396);
  not1 I011_407(w_011_407, w_006_168);
  not1 I011_409(w_011_409, w_007_393);
  and2 I011_410(w_011_410, w_010_130, w_006_011);
  and2 I011_411(w_011_411, w_006_048, w_002_229);
  not1 I011_414(w_011_414, w_004_077);
  nand2 I011_416(w_011_416, w_008_210, w_003_029);
  or2  I011_419(w_011_419, w_002_405, w_009_331);
  not1 I011_420(w_011_420, w_008_266);
  nand2 I011_421(w_011_421, w_005_059, w_001_017);
  not1 I011_424(w_011_424, w_003_026);
  nand2 I011_426(w_011_426, w_010_220, w_004_121);
  nand2 I011_427(w_011_427, w_004_302, w_008_054);
  or2  I011_428(w_011_428, w_002_303, w_006_244);
  not1 I011_430(w_011_430, w_005_137);
  and2 I011_431(w_011_431, w_007_204, w_003_040);
  or2  I011_433(w_011_433, w_001_023, w_009_186);
  and2 I011_435(w_011_435, w_001_005, w_008_584);
  nand2 I011_437(w_011_437, w_000_505, w_008_703);
  or2  I011_438(w_011_438, w_002_459, w_000_266);
  or2  I011_439(w_011_439, w_003_025, w_004_293);
  and2 I011_440(w_011_440, w_000_032, w_002_374);
  and2 I011_441(w_011_441, w_008_207, w_008_441);
  not1 I011_443(w_011_443, w_003_038);
  nand2 I011_444(w_011_444, w_009_004, w_000_696);
  nand2 I011_446(w_011_446, w_003_056, w_000_578);
  not1 I011_450(w_011_450, w_003_022);
  and2 I011_455(w_011_455, w_009_038, w_004_089);
  and2 I011_457(w_011_457, w_008_290, w_006_029);
  and2 I011_458(w_011_458, w_005_072, w_004_253);
  and2 I011_459(w_011_459, w_003_064, w_006_110);
  and2 I011_460(w_011_460, w_000_222, w_008_023);
  or2  I011_461(w_011_461, w_001_033, w_004_040);
  or2  I011_462(w_011_462, w_005_099, w_002_134);
  not1 I011_463(w_011_463, w_005_067);
  and2 I011_465(w_011_465, w_002_683, w_010_056);
  nand2 I011_466(w_011_466, w_005_199, w_003_025);
  or2  I011_467(w_011_467, w_000_185, w_001_019);
  not1 I011_468(w_011_468, w_004_486);
  nand2 I011_469(w_011_469, w_007_103, w_007_135);
  or2  I011_471(w_011_471, w_007_033, w_000_342);
  and2 I011_472(w_011_472, w_010_399, w_000_540);
  or2  I011_473(w_011_473, w_003_033, w_000_056);
  or2  I011_474(w_011_474, w_002_502, w_007_153);
  and2 I011_477(w_011_477, w_006_165, w_003_035);
  or2  I011_480(w_011_480, w_009_281, w_000_231);
  and2 I011_481(w_011_481, w_006_096, w_001_008);
  not1 I011_486(w_011_486, w_010_609);
  nand2 I011_489(w_011_489, w_004_022, w_007_177);
  nand2 I011_490(w_011_490, w_004_063, w_005_272);
  not1 I011_491(w_011_491, w_005_220);
  or2  I011_492(w_011_492, w_005_155, w_006_245);
  and2 I011_494(w_011_494, w_002_504, w_004_343);
  and2 I011_500(w_011_500, w_003_043, w_007_237);
  not1 I011_502(w_011_502, w_005_026);
  or2  I011_503(w_011_503, w_010_447, w_006_053);
  not1 I011_504(w_011_504, w_003_029);
  not1 I011_508(w_011_508, w_006_161);
  or2  I011_510(w_011_510, w_008_526, w_000_320);
  and2 I011_511(w_011_511, w_003_009, w_009_119);
  or2  I011_512(w_011_512, w_000_624, w_007_426);
  nand2 I011_514(w_011_514, w_003_013, w_001_003);
  or2  I011_515(w_011_515, w_005_205, w_009_060);
  or2  I011_517(w_011_517, w_007_208, w_003_035);
  or2  I011_519(w_011_519, w_009_194, w_005_193);
  or2  I011_520(w_011_520, w_009_159, w_005_044);
  nand2 I011_521(w_011_521, w_008_724, w_004_232);
  or2  I011_523(w_011_523, w_010_357, w_001_026);
  nand2 I011_525(w_011_525, w_000_422, w_000_659);
  nand2 I011_527(w_011_527, w_009_147, w_007_060);
  nand2 I011_529(w_011_529, w_010_444, w_007_101);
  or2  I011_530(w_011_530, w_006_101, w_007_184);
  or2  I011_531(w_011_531, w_007_105, w_004_017);
  nand2 I011_532(w_011_532, w_002_677, w_004_269);
  nand2 I011_533(w_011_533, w_004_048, w_000_366);
  not1 I011_538(w_011_538, w_005_071);
  or2  I011_539(w_011_539, w_007_300, w_005_112);
  nand2 I011_540(w_011_540, w_007_350, w_004_148);
  or2  I011_541(w_011_541, w_004_015, w_007_472);
  or2  I011_542(w_011_542, w_005_072, w_000_305);
  and2 I011_543(w_011_543, w_006_188, w_005_023);
  and2 I011_544(w_011_544, w_006_014, w_002_541);
  not1 I011_545(w_011_545, w_001_031);
  not1 I011_546(w_011_546, w_006_014);
  or2  I011_548(w_011_548, w_004_354, w_002_415);
  nand2 I011_549(w_011_549, w_008_488, w_008_525);
  and2 I011_550(w_011_550, w_002_265, w_009_418);
  not1 I011_551(w_011_551, w_004_175);
  nand2 I011_554(w_011_554, w_003_007, w_006_200);
  and2 I011_555(w_011_555, w_008_421, w_006_024);
  or2  I011_556(w_011_556, w_004_256, w_004_272);
  or2  I011_557(w_011_557, w_002_690, w_005_230);
  and2 I011_558(w_011_558, w_003_037, w_008_656);
  and2 I011_559(w_011_559, w_002_212, w_001_030);
  not1 I011_560(w_011_560, w_009_462);
  and2 I011_561(w_011_561, w_002_468, w_010_614);
  or2  I011_562(w_011_562, w_003_016, w_007_391);
  and2 I011_563(w_011_563, w_009_033, w_003_077);
  not1 I011_564(w_011_564, w_006_187);
  not1 I011_565(w_011_565, w_009_116);
  or2  I011_566(w_011_566, w_009_194, w_000_006);
  or2  I011_567(w_011_567, w_004_096, w_010_613);
  and2 I011_568(w_011_568, w_002_633, w_010_089);
  not1 I011_569(w_011_569, w_003_020);
  and2 I011_570(w_011_570, w_006_237, w_009_073);
  and2 I011_571(w_011_571, w_007_179, w_005_131);
  or2  I011_572(w_011_572, w_002_077, w_002_309);
  or2  I011_575(w_011_575, w_002_655, w_007_415);
  or2  I011_576(w_011_576, w_007_142, w_007_126);
  and2 I011_579(w_011_579, w_006_227, w_000_421);
  not1 I011_582(w_011_582, w_003_052);
  not1 I011_583(w_011_583, w_008_264);
  not1 I011_586(w_011_586, w_007_149);
  not1 I011_587(w_011_587, w_003_079);
  nand2 I011_589(w_011_589, w_007_113, w_006_022);
  not1 I011_591(w_011_591, w_009_361);
  not1 I011_592(w_011_592, w_006_097);
  nand2 I011_594(w_011_594, w_000_055, w_007_179);
  and2 I011_596(w_011_596, w_008_114, w_005_028);
  nand2 I011_597(w_011_597, w_003_009, w_009_150);
  and2 I011_599(w_011_599, w_001_034, w_000_416);
  and2 I011_603(w_011_603, w_005_080, w_010_775);
  not1 I011_605(w_011_605, w_007_380);
  nand2 I011_606(w_011_606, w_007_314, w_007_232);
  not1 I011_607(w_011_607, w_006_156);
  not1 I011_611(w_011_611, w_002_230);
  and2 I011_615(w_011_615, w_005_031, w_008_078);
  nand2 I011_616(w_011_616, w_006_078, w_003_074);
  nand2 I011_617(w_011_617, w_010_358, w_007_100);
  and2 I011_618(w_011_618, w_004_265, w_002_219);
  or2  I011_620(w_011_620, w_004_418, w_009_019);
  not1 I011_622(w_011_622, w_005_160);
  not1 I011_624(w_011_624, w_009_403);
  not1 I011_626(w_011_626, w_002_106);
  and2 I011_629(w_011_629, w_005_288, w_001_035);
  or2  I011_630(w_011_630, w_006_032, w_008_084);
  and2 I011_631(w_011_631, w_004_346, w_007_088);
  or2  I011_632(w_011_632, w_002_488, w_006_235);
  not1 I011_633(w_011_633, w_001_020);
  nand2 I011_634(w_011_634, w_004_281, w_006_227);
  not1 I011_635(w_011_635, w_010_207);
  or2  I011_637(w_011_637, w_003_077, w_004_212);
  and2 I011_639(w_011_639, w_001_002, w_008_419);
  and2 I011_641(w_011_641, w_000_704, w_003_081);
  nand2 I011_642(w_011_642, w_000_181, w_006_081);
  or2  I012_000(w_012_000, w_000_297, w_011_337);
  nand2 I012_001(w_012_001, w_010_343, w_002_231);
  nand2 I012_002(w_012_002, w_005_058, w_001_004);
  not1 I012_003(w_012_003, w_008_061);
  nand2 I012_004(w_012_004, w_000_106, w_000_073);
  nand2 I012_005(w_012_005, w_010_308, w_004_145);
  nand2 I012_006(w_012_006, w_010_083, w_008_254);
  or2  I012_007(w_012_007, w_007_144, w_004_265);
  nand2 I012_008(w_012_008, w_011_048, w_011_017);
  or2  I012_009(w_012_009, w_000_157, w_004_436);
  not1 I012_010(w_012_010, w_007_114);
  and2 I012_011(w_012_011, w_007_221, w_007_259);
  or2  I012_012(w_012_012, w_011_596, w_000_542);
  and2 I012_013(w_012_013, w_008_348, w_009_584);
  not1 I012_015(w_012_015, w_011_205);
  nand2 I012_016(w_012_016, w_011_071, w_011_035);
  and2 I012_017(w_012_017, w_010_183, w_001_033);
  and2 I012_018(w_012_018, w_000_155, w_005_009);
  and2 I012_019(w_012_019, w_006_070, w_008_622);
  not1 I012_020(w_012_020, w_009_128);
  nand2 I012_021(w_012_021, w_002_360, w_003_000);
  not1 I012_022(w_012_022, w_002_012);
  or2  I012_023(w_012_023, w_005_088, w_009_416);
  not1 I012_024(w_012_024, w_007_117);
  nand2 I012_025(w_012_025, w_005_236, w_008_389);
  and2 I012_026(w_012_026, w_000_693, w_006_045);
  or2  I012_027(w_012_027, w_001_009, w_010_619);
  nand2 I012_028(w_012_028, w_000_179, w_002_655);
  or2  I012_029(w_012_029, w_004_219, w_003_041);
  or2  I012_030(w_012_030, w_004_009, w_008_431);
  and2 I012_031(w_012_031, w_003_047, w_011_043);
  not1 I012_032(w_012_032, w_000_271);
  nand2 I012_033(w_012_033, w_006_121, w_000_311);
  not1 I012_034(w_012_034, w_010_131);
  or2  I012_035(w_012_035, w_002_662, w_004_268);
  and2 I012_036(w_012_036, w_000_197, w_011_502);
  nand2 I012_037(w_012_037, w_007_029, w_011_143);
  and2 I012_038(w_012_038, w_006_203, w_003_009);
  or2  I012_039(w_012_039, w_007_365, w_004_202);
  nand2 I012_040(w_012_040, w_004_003, w_001_033);
  and2 I012_041(w_012_041, w_002_193, w_007_172);
  nand2 I012_042(w_012_042, w_003_060, w_008_214);
  or2  I012_043(w_012_043, w_011_121, w_008_074);
  nand2 I012_044(w_012_044, w_000_125, w_007_348);
  nand2 I012_045(w_012_045, w_004_099, w_000_093);
  or2  I012_046(w_012_046, w_011_150, w_011_508);
  and2 I012_047(w_012_047, w_007_233, w_009_078);
  or2  I012_048(w_012_048, w_008_349, w_000_252);
  nand2 I012_049(w_012_049, w_005_068, w_004_280);
  not1 I012_050(w_012_050, w_000_646);
  nand2 I012_051(w_012_051, w_011_194, w_006_085);
  not1 I012_052(w_012_052, w_011_041);
  nand2 I012_053(w_012_053, w_002_230, w_010_667);
  not1 I012_054(w_012_054, w_006_076);
  nand2 I012_055(w_012_055, w_000_703, w_003_005);
  and2 I012_056(w_012_056, w_011_437, w_001_026);
  not1 I012_057(w_012_057, w_003_003);
  not1 I012_058(w_012_058, w_010_077);
  or2  I012_059(w_012_059, w_008_020, w_000_030);
  nand2 I012_060(w_012_060, w_001_008, w_005_076);
  and2 I012_061(w_012_061, w_000_593, w_002_162);
  and2 I012_062(w_012_062, w_003_066, w_011_433);
  not1 I012_063(w_012_063, w_010_070);
  not1 I012_065(w_012_065, w_005_285);
  nand2 I012_066(w_012_066, w_005_305, w_000_652);
  and2 I012_067(w_012_067, w_005_096, w_006_052);
  not1 I012_068(w_012_068, w_010_645);
  or2  I012_069(w_012_069, w_001_020, w_004_217);
  and2 I012_070(w_012_070, w_001_015, w_006_041);
  and2 I012_071(w_012_071, w_000_396, w_003_066);
  not1 I012_072(w_012_072, w_000_062);
  not1 I012_073(w_012_073, w_010_719);
  not1 I012_074(w_012_074, w_002_228);
  nand2 I012_075(w_012_075, w_004_188, w_011_087);
  and2 I012_076(w_012_076, w_004_153, w_005_158);
  nand2 I012_077(w_012_077, w_004_165, w_004_325);
  nand2 I012_078(w_012_078, w_008_322, w_004_274);
  or2  I012_079(w_012_079, w_004_192, w_002_502);
  and2 I012_080(w_012_080, w_000_705, w_002_046);
  not1 I012_081(w_012_081, w_009_350);
  and2 I012_082(w_012_082, w_000_632, w_004_344);
  and2 I012_083(w_012_083, w_010_021, w_011_007);
  not1 I012_084(w_012_084, w_008_528);
  not1 I012_086(w_012_086, w_008_719);
  not1 I012_087(w_012_087, w_002_669);
  or2  I012_088(w_012_088, w_007_073, w_011_213);
  nand2 I012_089(w_012_089, w_005_147, w_009_221);
  nand2 I012_090(w_012_090, w_006_173, w_008_614);
  nand2 I012_091(w_012_091, w_009_121, w_006_218);
  or2  I012_092(w_012_092, w_006_054, w_001_009);
  and2 I012_093(w_012_093, w_001_021, w_002_596);
  or2  I012_094(w_012_094, w_003_063, w_002_026);
  and2 I012_095(w_012_095, w_010_243, w_007_221);
  and2 I012_096(w_012_096, w_011_021, w_010_491);
  and2 I012_098(w_012_098, w_010_481, w_010_680);
  or2  I012_099(w_012_099, w_010_053, w_009_481);
  nand2 I012_101(w_012_101, w_009_006, w_002_288);
  not1 I012_102(w_012_102, w_011_519);
  nand2 I012_103(w_012_103, w_001_007, w_003_040);
  nand2 I012_104(w_012_104, w_004_208, w_003_048);
  nand2 I012_105(w_012_105, w_006_031, w_001_034);
  and2 I012_106(w_012_106, w_010_381, w_009_200);
  not1 I012_107(w_012_107, w_010_140);
  or2  I012_108(w_012_108, w_007_017, w_003_056);
  or2  I012_109(w_012_109, w_006_130, w_004_287);
  or2  I012_110(w_012_110, w_007_390, w_004_089);
  and2 I012_111(w_012_111, w_008_710, w_011_278);
  and2 I012_112(w_012_112, w_004_020, w_008_262);
  and2 I012_113(w_012_113, w_006_014, w_010_592);
  nand2 I012_114(w_012_114, w_011_167, w_010_726);
  not1 I012_115(w_012_115, w_007_107);
  or2  I012_116(w_012_116, w_003_003, w_003_061);
  not1 I012_118(w_012_118, w_007_292);
  not1 I012_119(w_012_119, w_009_545);
  not1 I012_120(w_012_120, w_000_041);
  or2  I012_121(w_012_121, w_008_135, w_011_450);
  nand2 I012_122(w_012_122, w_010_301, w_006_043);
  nand2 I012_123(w_012_123, w_001_019, w_008_090);
  nand2 I012_124(w_012_124, w_001_016, w_002_271);
  or2  I012_125(w_012_125, w_000_502, w_000_437);
  and2 I012_126(w_012_126, w_002_534, w_010_238);
  nand2 I012_127(w_012_127, w_011_051, w_011_411);
  not1 I012_129(w_012_129, w_000_314);
  or2  I012_130(w_012_130, w_009_404, w_008_694);
  not1 I012_131(w_012_131, w_002_165);
  nand2 I012_132(w_012_132, w_003_072, w_011_045);
  or2  I012_134(w_012_134, w_005_202, w_008_604);
  or2  I012_135(w_012_135, w_003_063, w_006_238);
  and2 I012_136(w_012_136, w_007_258, w_005_042);
  not1 I012_137(w_012_137, w_006_126);
  and2 I012_138(w_012_138, w_008_291, w_003_050);
  or2  I012_140(w_012_140, w_008_444, w_007_386);
  or2  I012_141(w_012_141, w_007_190, w_007_076);
  and2 I012_142(w_012_142, w_001_017, w_008_284);
  and2 I012_143(w_012_143, w_002_516, w_007_212);
  not1 I012_145(w_012_145, w_003_028);
  or2  I012_147(w_012_147, w_000_318, w_000_354);
  or2  I012_149(w_012_149, w_008_332, w_005_086);
  or2  I012_150(w_012_150, w_007_473, w_000_515);
  and2 I012_151(w_012_151, w_011_056, w_002_302);
  and2 I012_152(w_012_152, w_007_360, w_003_071);
  nand2 I012_153(w_012_153, w_000_294, w_001_000);
  and2 I012_154(w_012_154, w_001_020, w_001_035);
  not1 I012_155(w_012_155, w_010_004);
  nand2 I012_157(w_012_157, w_003_075, w_011_126);
  nand2 I012_158(w_012_158, w_003_024, w_001_014);
  nand2 I012_162(w_012_162, w_006_168, w_007_129);
  and2 I012_163(w_012_163, w_001_009, w_009_243);
  and2 I012_164(w_012_164, w_011_567, w_007_279);
  not1 I012_165(w_012_165, w_006_056);
  and2 I012_167(w_012_167, w_009_473, w_011_079);
  nand2 I012_168(w_012_168, w_009_118, w_010_235);
  and2 I012_169(w_012_169, w_005_046, w_009_074);
  nand2 I012_170(w_012_170, w_006_065, w_011_286);
  or2  I012_171(w_012_171, w_007_117, w_007_023);
  nand2 I012_172(w_012_172, w_005_145, w_003_060);
  nand2 I012_174(w_012_174, w_009_508, w_003_021);
  nand2 I012_175(w_012_175, w_008_149, w_001_006);
  nand2 I012_176(w_012_176, w_000_683, w_009_020);
  or2  I012_177(w_012_177, w_002_619, w_002_078);
  and2 I012_178(w_012_178, w_006_087, w_001_035);
  nand2 I012_179(w_012_179, w_010_777, w_008_543);
  and2 I012_181(w_012_181, w_009_394, w_001_036);
  nand2 I012_182(w_012_182, w_008_559, w_003_062);
  nand2 I012_183(w_012_183, w_008_048, w_002_099);
  or2  I012_185(w_012_185, w_007_422, w_000_517);
  or2  I012_187(w_012_187, w_002_018, w_005_207);
  and2 I012_188(w_012_188, w_006_164, w_004_159);
  or2  I012_189(w_012_189, w_007_091, w_008_083);
  or2  I012_190(w_012_190, w_002_182, w_008_688);
  nand2 I012_191(w_012_191, w_005_087, w_010_418);
  or2  I012_192(w_012_192, w_006_005, w_002_083);
  not1 I012_193(w_012_193, w_003_020);
  and2 I012_194(w_012_194, w_001_027, w_008_271);
  or2  I012_198(w_012_198, w_007_000, w_010_745);
  nand2 I012_199(w_012_199, w_000_292, w_001_019);
  or2  I012_200(w_012_200, w_005_262, w_002_705);
  and2 I012_201(w_012_201, w_009_598, w_003_057);
  or2  I012_202(w_012_202, w_006_192, w_008_615);
  nand2 I012_203(w_012_203, w_006_250, w_001_035);
  nand2 I012_204(w_012_204, w_011_446, w_011_481);
  nand2 I012_205(w_012_205, w_006_200, w_007_281);
  not1 I012_206(w_012_206, w_004_060);
  nand2 I012_207(w_012_207, w_011_123, w_003_077);
  and2 I012_208(w_012_208, w_010_622, w_009_417);
  nand2 I012_209(w_012_209, w_010_232, w_007_284);
  or2  I012_210(w_012_210, w_000_167, w_000_295);
  or2  I012_211(w_012_211, w_011_329, w_004_122);
  nand2 I012_212(w_012_212, w_011_437, w_001_019);
  not1 I012_213(w_012_213, w_008_302);
  and2 I012_214(w_012_214, w_003_040, w_004_192);
  or2  I012_215(w_012_215, w_001_023, w_004_241);
  nand2 I012_216(w_012_216, w_011_235, w_008_636);
  not1 I012_217(w_012_217, w_000_483);
  nand2 I012_219(w_012_219, w_006_007, w_008_434);
  nand2 I012_221(w_012_221, w_005_254, w_008_319);
  not1 I012_223(w_012_223, w_001_009);
  and2 I012_224(w_012_224, w_001_008, w_008_149);
  and2 I012_225(w_012_225, w_011_071, w_008_482);
  nand2 I012_226(w_012_226, w_008_468, w_008_033);
  and2 I012_227(w_012_227, w_010_385, w_000_671);
  nand2 I012_228(w_012_228, w_000_190, w_000_525);
  or2  I012_229(w_012_229, w_000_510, w_011_617);
  not1 I012_230(w_012_230, w_007_071);
  not1 I012_231(w_012_231, w_003_062);
  nand2 I012_232(w_012_232, w_003_049, w_007_127);
  nand2 I012_233(w_012_233, w_007_277, w_003_057);
  or2  I012_234(w_012_234, w_001_027, w_009_119);
  and2 I012_235(w_012_235, w_010_491, w_004_093);
  and2 I012_236(w_012_236, w_009_313, w_007_284);
  and2 I012_237(w_012_237, w_003_049, w_006_074);
  not1 I012_238(w_012_238, w_005_201);
  not1 I012_239(w_012_239, w_004_362);
  or2  I012_240(w_012_240, w_000_191, w_008_496);
  or2  I012_241(w_012_241, w_010_298, w_006_117);
  not1 I012_242(w_012_242, w_008_314);
  nand2 I012_243(w_012_243, w_004_019, w_000_485);
  not1 I012_244(w_012_244, w_002_329);
  or2  I012_245(w_012_245, w_004_360, w_004_210);
  or2  I012_246(w_012_246, w_009_216, w_010_548);
  or2  I012_247(w_012_247, w_002_291, w_005_230);
  nand2 I012_249(w_012_249, w_007_209, w_002_035);
  and2 I012_250(w_012_250, w_002_433, w_002_256);
  not1 I012_252(w_012_252, w_004_004);
  and2 I012_253(w_012_253, w_001_023, w_010_649);
  nand2 I012_254(w_012_254, w_000_141, w_005_282);
  or2  I012_255(w_012_255, w_004_011, w_004_239);
  not1 I012_256(w_012_256, w_000_448);
  and2 I012_257(w_012_257, w_007_228, w_006_228);
  not1 I012_258(w_012_258, w_006_037);
  not1 I012_259(w_012_259, w_011_321);
  not1 I012_260(w_012_260, w_009_193);
  and2 I012_261(w_012_261, w_008_063, w_005_312);
  nand2 I012_262(w_012_262, w_002_008, w_010_760);
  or2  I012_263(w_012_263, w_009_480, w_008_343);
  and2 I012_264(w_012_264, w_000_031, w_008_724);
  not1 I012_267(w_012_267, w_007_232);
  not1 I012_268(w_012_268, w_005_096);
  or2  I012_269(w_012_269, w_011_424, w_003_077);
  or2  I012_270(w_012_270, w_000_706, w_009_499);
  and2 I012_271(w_012_271, w_001_012, w_000_349);
  nand2 I012_272(w_012_272, w_009_149, w_011_220);
  and2 I012_273(w_012_273, w_001_026, w_000_465);
  and2 I012_274(w_012_274, w_011_249, w_010_136);
  or2  I012_275(w_012_275, w_003_084, w_009_251);
  nand2 I012_276(w_012_276, w_010_407, w_003_003);
  nand2 I012_277(w_012_277, w_008_428, w_009_532);
  or2  I012_278(w_012_278, w_009_209, w_000_056);
  not1 I012_279(w_012_279, w_001_034);
  and2 I012_281(w_012_281, w_005_046, w_005_103);
  or2  I012_282(w_012_282, w_002_192, w_008_188);
  not1 I012_285(w_012_285, w_005_007);
  and2 I012_286(w_012_286, w_010_005, w_007_043);
  or2  I012_287(w_012_287, w_003_016, w_002_412);
  and2 I012_288(w_012_288, w_011_353, w_001_031);
  or2  I012_289(w_012_289, w_002_682, w_001_032);
  not1 I012_290(w_012_290, w_011_374);
  or2  I012_291(w_012_291, w_011_078, w_006_238);
  and2 I012_292(w_012_292, w_003_079, w_004_225);
  and2 I012_293(w_012_293, w_004_110, w_005_068);
  nand2 I012_294(w_012_294, w_011_156, w_008_055);
  or2  I012_295(w_012_295, w_009_549, w_002_039);
  nand2 I012_296(w_012_296, w_007_223, w_005_025);
  nand2 I012_297(w_012_297, w_011_018, w_010_057);
  nand2 I012_298(w_012_298, w_010_716, w_000_495);
  or2  I012_299(w_012_299, w_004_003, w_009_058);
  not1 I012_300(w_012_300, w_008_085);
  or2  I012_301(w_012_301, w_004_492, w_006_092);
  or2  I012_302(w_012_302, w_001_031, w_005_037);
  nand2 I012_303(w_012_303, w_002_219, w_006_236);
  not1 I012_304(w_012_304, w_004_036);
  or2  I012_305(w_012_305, w_007_462, w_005_275);
  nand2 I012_306(w_012_306, w_010_149, w_000_707);
  not1 I012_308(w_012_308, w_011_459);
  nand2 I012_309(w_012_309, w_000_561, w_000_596);
  and2 I012_310(w_012_310, w_003_028, w_002_524);
  not1 I012_311(w_012_311, w_011_271);
  nand2 I012_312(w_012_312, w_006_227, w_000_144);
  or2  I012_313(w_012_313, w_002_645, w_005_263);
  and2 I012_314(w_012_314, w_006_176, w_000_396);
  not1 I012_315(w_012_315, w_011_407);
  or2  I012_316(w_012_316, w_003_083, w_006_044);
  and2 I012_317(w_012_317, w_009_412, w_011_549);
  or2  I012_319(w_012_319, w_004_148, w_005_002);
  nand2 I012_320(w_012_320, w_008_485, w_008_178);
  or2  I012_321(w_012_321, w_007_354, w_001_021);
  and2 I012_322(w_012_322, w_001_035, w_010_452);
  nand2 I012_323(w_012_323, w_004_048, w_003_070);
  and2 I012_324(w_012_324, w_002_426, w_006_138);
  nand2 I012_325(w_012_325, w_007_340, w_001_027);
  nand2 I012_327(w_012_327, w_006_105, w_002_028);
  not1 I012_328(w_012_328, w_002_497);
  not1 I012_330(w_012_330, w_011_529);
  not1 I012_331(w_012_331, w_006_156);
  or2  I012_332(w_012_332, w_010_507, w_000_307);
  and2 I012_333(w_012_333, w_005_039, w_004_366);
  and2 I012_335(w_012_335, w_007_124, w_006_029);
  nand2 I012_336(w_012_336, w_011_490, w_003_082);
  and2 I012_337(w_012_337, w_003_079, w_002_669);
  or2  I012_338(w_012_338, w_007_153, w_004_222);
  not1 I012_340(w_012_340, w_000_524);
  not1 I012_342(w_012_342, w_006_008);
  not1 I012_344(w_012_344, w_011_069);
  or2  I012_345(w_012_345, w_000_619, w_006_085);
  not1 I012_346(w_012_346, w_009_549);
  not1 I012_347(w_012_347, w_000_481);
  and2 I012_348(w_012_348, w_002_037, w_004_067);
  or2  I012_350(w_012_350, w_001_036, w_008_339);
  and2 I013_000(w_013_000, w_007_219, w_002_586);
  nand2 I013_001(w_013_001, w_003_075, w_004_116);
  not1 I013_002(w_013_002, w_001_011);
  not1 I013_003(w_013_003, w_002_501);
  and2 I013_004(w_013_004, w_004_193, w_006_192);
  nand2 I013_005(w_013_005, w_011_099, w_000_354);
  nand2 I013_006(w_013_006, w_003_002, w_004_255);
  nand2 I013_008(w_013_008, w_005_054, w_011_379);
  or2  I013_009(w_013_009, w_002_085, w_008_015);
  nand2 I013_010(w_013_010, w_012_165, w_012_107);
  or2  I013_011(w_013_011, w_007_300, w_006_072);
  not1 I013_012(w_013_012, w_006_231);
  not1 I013_013(w_013_013, w_011_233);
  nand2 I013_015(w_013_015, w_009_414, w_006_002);
  nand2 I013_016(w_013_016, w_010_593, w_005_303);
  or2  I013_017(w_013_017, w_004_371, w_004_474);
  not1 I013_020(w_013_020, w_004_198);
  or2  I013_021(w_013_021, w_011_300, w_010_109);
  not1 I013_022(w_013_022, w_004_107);
  not1 I013_023(w_013_023, w_001_023);
  and2 I013_024(w_013_024, w_012_145, w_007_422);
  and2 I013_025(w_013_025, w_004_255, w_007_088);
  nand2 I013_026(w_013_026, w_001_021, w_008_320);
  or2  I013_027(w_013_027, w_004_506, w_012_134);
  and2 I013_028(w_013_028, w_010_004, w_005_024);
  and2 I013_029(w_013_029, w_009_513, w_004_093);
  and2 I013_030(w_013_030, w_007_206, w_001_020);
  and2 I013_031(w_013_031, w_009_079, w_007_144);
  nand2 I013_032(w_013_032, w_007_063, w_006_162);
  and2 I013_034(w_013_034, w_000_424, w_008_035);
  or2  I013_035(w_013_035, w_001_008, w_012_129);
  nand2 I013_036(w_013_036, w_005_316, w_004_501);
  or2  I013_037(w_013_037, w_005_199, w_002_176);
  or2  I013_040(w_013_040, w_002_434, w_006_060);
  or2  I013_041(w_013_041, w_000_191, w_008_292);
  and2 I013_042(w_013_042, w_003_015, w_003_066);
  or2  I013_043(w_013_043, w_006_009, w_000_323);
  not1 I013_044(w_013_044, w_002_180);
  nand2 I013_046(w_013_046, w_009_053, w_008_003);
  or2  I013_047(w_013_047, w_001_014, w_001_005);
  or2  I013_048(w_013_048, w_011_446, w_011_236);
  not1 I013_049(w_013_049, w_003_048);
  nand2 I013_050(w_013_050, w_009_117, w_008_220);
  or2  I013_053(w_013_053, w_012_119, w_007_128);
  and2 I013_054(w_013_054, w_011_089, w_007_334);
  or2  I013_055(w_013_055, w_006_079, w_006_055);
  not1 I013_059(w_013_059, w_000_023);
  or2  I013_060(w_013_060, w_012_015, w_004_267);
  nand2 I013_061(w_013_061, w_004_317, w_001_017);
  and2 I013_062(w_013_062, w_003_037, w_002_071);
  not1 I013_063(w_013_063, w_009_054);
  and2 I013_064(w_013_064, w_002_024, w_004_220);
  or2  I013_065(w_013_065, w_008_608, w_002_326);
  not1 I013_066(w_013_066, w_002_702);
  nand2 I013_067(w_013_067, w_002_619, w_000_079);
  not1 I013_068(w_013_068, w_004_238);
  nand2 I013_069(w_013_069, w_005_177, w_005_306);
  and2 I013_070(w_013_070, w_001_028, w_010_263);
  and2 I013_071(w_013_071, w_012_200, w_004_061);
  and2 I013_072(w_013_072, w_012_221, w_012_041);
  and2 I013_073(w_013_073, w_003_039, w_001_023);
  or2  I013_074(w_013_074, w_003_017, w_009_118);
  not1 I013_075(w_013_075, w_011_592);
  not1 I013_076(w_013_076, w_005_098);
  nand2 I013_077(w_013_077, w_006_122, w_003_008);
  nand2 I013_078(w_013_078, w_004_269, w_003_037);
  not1 I013_079(w_013_079, w_004_186);
  not1 I013_080(w_013_080, w_007_186);
  not1 I013_081(w_013_081, w_012_172);
  or2  I013_083(w_013_083, w_011_473, w_000_663);
  nand2 I013_086(w_013_086, w_003_012, w_001_034);
  and2 I013_087(w_013_087, w_003_010, w_008_605);
  nand2 I013_088(w_013_088, w_009_051, w_011_170);
  and2 I013_089(w_013_089, w_002_288, w_003_048);
  not1 I013_090(w_013_090, w_005_058);
  and2 I013_091(w_013_091, w_010_144, w_006_014);
  not1 I013_092(w_013_092, w_000_405);
  or2  I013_093(w_013_093, w_006_226, w_011_379);
  nand2 I013_095(w_013_095, w_000_034, w_005_244);
  not1 I013_096(w_013_096, w_007_051);
  and2 I013_097(w_013_097, w_010_365, w_008_010);
  not1 I013_098(w_013_098, w_007_154);
  nand2 I013_099(w_013_099, w_010_156, w_006_085);
  or2  I013_100(w_013_100, w_012_270, w_012_328);
  nand2 I013_102(w_013_102, w_007_094, w_002_047);
  not1 I013_103(w_013_103, w_012_010);
  not1 I013_104(w_013_104, w_011_085);
  not1 I013_105(w_013_105, w_005_007);
  or2  I013_106(w_013_106, w_004_377, w_001_034);
  or2  I013_107(w_013_107, w_008_555, w_009_126);
  nand2 I013_108(w_013_108, w_004_503, w_001_035);
  not1 I013_109(w_013_109, w_009_351);
  not1 I013_110(w_013_110, w_009_445);
  or2  I013_111(w_013_111, w_006_044, w_009_462);
  not1 I013_112(w_013_112, w_009_068);
  or2  I013_114(w_013_114, w_004_429, w_007_120);
  nand2 I013_115(w_013_115, w_000_363, w_008_494);
  nand2 I013_116(w_013_116, w_003_013, w_006_233);
  nand2 I013_117(w_013_117, w_004_230, w_004_216);
  and2 I013_118(w_013_118, w_002_230, w_007_267);
  nand2 I013_121(w_013_121, w_012_119, w_001_013);
  or2  I013_122(w_013_122, w_009_060, w_003_044);
  or2  I013_123(w_013_123, w_009_084, w_008_105);
  nand2 I013_124(w_013_124, w_012_323, w_010_342);
  and2 I013_125(w_013_125, w_004_133, w_005_134);
  not1 I013_126(w_013_126, w_001_035);
  or2  I013_127(w_013_127, w_008_755, w_011_088);
  or2  I013_128(w_013_128, w_012_296, w_001_002);
  and2 I013_129(w_013_129, w_006_005, w_012_236);
  or2  I013_130(w_013_130, w_008_341, w_004_495);
  nand2 I013_131(w_013_131, w_001_001, w_003_003);
  or2  I013_132(w_013_132, w_010_412, w_011_634);
  or2  I013_133(w_013_133, w_000_094, w_008_449);
  or2  I013_134(w_013_134, w_002_145, w_004_155);
  not1 I013_135(w_013_135, w_006_009);
  not1 I013_136(w_013_136, w_006_245);
  nand2 I013_137(w_013_137, w_003_053, w_002_653);
  not1 I013_138(w_013_138, w_005_243);
  not1 I013_139(w_013_139, w_001_033);
  or2  I013_140(w_013_140, w_011_237, w_008_376);
  not1 I013_141(w_013_141, w_003_083);
  nand2 I013_142(w_013_142, w_009_107, w_012_298);
  nand2 I013_144(w_013_144, w_008_664, w_004_207);
  and2 I013_145(w_013_145, w_006_175, w_001_002);
  or2  I013_146(w_013_146, w_003_009, w_002_047);
  and2 I013_147(w_013_147, w_012_335, w_012_164);
  and2 I013_148(w_013_148, w_012_138, w_004_280);
  not1 I013_150(w_013_150, w_000_334);
  not1 I013_151(w_013_151, w_006_251);
  or2  I013_153(w_013_153, w_007_154, w_005_060);
  nand2 I013_154(w_013_154, w_008_029, w_001_000);
  nand2 I013_155(w_013_155, w_006_010, w_001_022);
  or2  I013_156(w_013_156, w_002_472, w_001_015);
  nand2 I013_157(w_013_157, w_008_387, w_011_527);
  or2  I013_158(w_013_158, w_006_078, w_005_248);
  not1 I013_159(w_013_159, w_007_448);
  not1 I013_160(w_013_160, w_012_060);
  or2  I013_161(w_013_161, w_009_441, w_005_290);
  or2  I013_162(w_013_162, w_000_579, w_011_015);
  and2 I013_163(w_013_163, w_002_487, w_004_415);
  not1 I013_164(w_013_164, w_012_002);
  nand2 I013_165(w_013_165, w_012_201, w_001_036);
  and2 I013_166(w_013_166, w_007_453, w_001_011);
  or2  I013_168(w_013_168, w_003_084, w_007_098);
  or2  I013_169(w_013_169, w_007_113, w_011_427);
  nand2 I013_170(w_013_170, w_004_394, w_006_089);
  or2  I013_171(w_013_171, w_001_016, w_010_561);
  and2 I013_172(w_013_172, w_004_420, w_009_342);
  not1 I013_174(w_013_174, w_008_560);
  and2 I013_175(w_013_175, w_004_183, w_006_074);
  and2 I013_176(w_013_176, w_007_053, w_007_039);
  or2  I013_178(w_013_178, w_010_327, w_007_218);
  nand2 I013_179(w_013_179, w_005_112, w_002_067);
  not1 I013_180(w_013_180, w_000_280);
  or2  I013_181(w_013_181, w_011_393, w_000_061);
  not1 I013_183(w_013_183, w_003_030);
  not1 I013_184(w_013_184, w_003_018);
  nand2 I013_185(w_013_185, w_010_584, w_009_363);
  not1 I013_186(w_013_186, w_002_085);
  not1 I013_188(w_013_188, w_001_019);
  nand2 I013_189(w_013_189, w_004_023, w_001_006);
  nand2 I013_190(w_013_190, w_000_393, w_009_130);
  nand2 I013_191(w_013_191, w_000_162, w_009_563);
  not1 I013_194(w_013_194, w_010_414);
  or2  I013_195(w_013_195, w_011_060, w_008_051);
  not1 I013_197(w_013_197, w_005_022);
  not1 I013_199(w_013_199, w_011_260);
  or2  I013_200(w_013_200, w_010_042, w_001_020);
  and2 I013_201(w_013_201, w_002_563, w_010_006);
  and2 I013_202(w_013_202, w_008_047, w_003_027);
  or2  I013_203(w_013_203, w_012_062, w_002_258);
  nand2 I013_204(w_013_204, w_007_151, w_003_070);
  not1 I013_205(w_013_205, w_006_070);
  and2 I013_206(w_013_206, w_006_078, w_003_027);
  not1 I013_207(w_013_207, w_005_061);
  not1 I013_208(w_013_208, w_007_142);
  or2  I013_209(w_013_209, w_012_114, w_006_209);
  or2  I013_210(w_013_210, w_007_272, w_008_300);
  nand2 I013_211(w_013_211, w_007_234, w_001_000);
  and2 I013_214(w_013_214, w_000_625, w_010_264);
  not1 I013_215(w_013_215, w_008_426);
  or2  I013_217(w_013_217, w_002_313, w_006_030);
  or2  I013_218(w_013_218, w_009_612, w_012_152);
  and2 I013_219(w_013_219, w_006_087, w_001_019);
  nand2 I013_220(w_013_220, w_009_321, w_005_114);
  and2 I013_222(w_013_222, w_012_291, w_012_305);
  nand2 I013_224(w_013_224, w_004_297, w_007_013);
  not1 I013_229(w_013_229, w_008_718);
  not1 I013_230(w_013_230, w_012_087);
  and2 I013_232(w_013_232, w_009_003, w_006_079);
  nand2 I013_235(w_013_235, w_012_036, w_006_140);
  or2  I013_236(w_013_236, w_003_031, w_011_078);
  not1 I013_237(w_013_237, w_003_030);
  or2  I013_239(w_013_239, w_007_096, w_010_060);
  and2 I013_242(w_013_242, w_006_230, w_008_361);
  nand2 I013_243(w_013_243, w_002_478, w_010_756);
  and2 I013_246(w_013_246, w_010_685, w_003_071);
  and2 I013_249(w_013_249, w_007_137, w_007_107);
  not1 I013_251(w_013_251, w_012_024);
  and2 I013_256(w_013_256, w_011_391, w_002_554);
  not1 I013_257(w_013_257, w_004_066);
  or2  I013_258(w_013_258, w_002_511, w_009_382);
  and2 I013_259(w_013_259, w_010_757, w_004_276);
  nand2 I013_260(w_013_260, w_012_091, w_007_088);
  not1 I013_263(w_013_263, w_010_405);
  and2 I013_265(w_013_265, w_010_076, w_011_063);
  or2  I013_266(w_013_266, w_010_020, w_009_478);
  or2  I013_269(w_013_269, w_005_162, w_006_110);
  and2 I013_270(w_013_270, w_003_005, w_007_120);
  not1 I013_272(w_013_272, w_000_210);
  and2 I013_274(w_013_274, w_000_709, w_012_010);
  or2  I013_275(w_013_275, w_000_251, w_009_222);
  not1 I013_278(w_013_278, w_003_020);
  and2 I013_279(w_013_279, w_003_037, w_000_133);
  nand2 I013_284(w_013_284, w_000_135, w_008_045);
  or2  I013_286(w_013_286, w_007_054, w_007_394);
  not1 I013_288(w_013_288, w_010_777);
  not1 I013_290(w_013_290, w_005_009);
  and2 I013_292(w_013_292, w_011_158, w_008_533);
  nand2 I013_293(w_013_293, w_006_007, w_000_487);
  and2 I013_295(w_013_295, w_006_088, w_008_502);
  not1 I013_296(w_013_296, w_004_034);
  and2 I013_297(w_013_297, w_009_553, w_006_024);
  or2  I013_301(w_013_301, w_012_303, w_003_068);
  and2 I013_302(w_013_302, w_000_462, w_008_084);
  not1 I013_303(w_013_303, w_005_113);
  and2 I013_305(w_013_305, w_002_597, w_005_128);
  not1 I013_306(w_013_306, w_012_223);
  or2  I013_307(w_013_307, w_005_006, w_001_017);
  not1 I013_309(w_013_309, w_001_004);
  nand2 I013_311(w_013_311, w_001_013, w_012_235);
  nand2 I013_313(w_013_313, w_008_428, w_004_161);
  or2  I013_316(w_013_316, w_011_062, w_008_533);
  or2  I013_317(w_013_317, w_009_433, w_005_252);
  nand2 I013_318(w_013_318, w_006_105, w_012_060);
  or2  I013_320(w_013_320, w_004_088, w_008_142);
  or2  I013_321(w_013_321, w_003_016, w_004_256);
  or2  I013_322(w_013_322, w_012_281, w_002_065);
  nand2 I013_323(w_013_323, w_012_247, w_009_486);
  nand2 I013_326(w_013_326, w_003_016, w_007_207);
  nand2 I013_327(w_013_327, w_003_058, w_002_094);
  not1 I013_329(w_013_329, w_004_242);
  and2 I013_330(w_013_330, w_000_438, w_012_049);
  nand2 I013_331(w_013_331, w_000_357, w_005_066);
  nand2 I013_332(w_013_332, w_005_155, w_005_099);
  or2  I013_334(w_013_334, w_005_164, w_004_156);
  or2  I013_339(w_013_339, w_005_209, w_012_338);
  not1 I013_340(w_013_340, w_012_229);
  not1 I013_344(w_013_344, w_012_141);
  or2  I013_346(w_013_346, w_006_251, w_009_016);
  or2  I013_348(w_013_348, w_008_071, w_002_067);
  not1 I013_349(w_013_349, w_001_025);
  nand2 I013_352(w_013_352, w_005_005, w_000_343);
  or2  I013_353(w_013_353, w_008_399, w_008_027);
  nand2 I013_357(w_013_357, w_000_285, w_000_604);
  and2 I013_358(w_013_358, w_005_135, w_008_241);
  not1 I013_359(w_013_359, w_000_565);
  not1 I013_361(w_013_361, w_005_077);
  and2 I013_363(w_013_363, w_005_074, w_008_760);
  nand2 I013_367(w_013_367, w_009_581, w_011_491);
  and2 I013_369(w_013_369, w_000_044, w_004_094);
  and2 I013_370(w_013_370, w_007_268, w_004_229);
  and2 I013_371(w_013_371, w_005_225, w_001_025);
  nand2 I013_372(w_013_372, w_009_411, w_012_058);
  and2 I013_373(w_013_373, w_007_471, w_011_124);
  not1 I013_374(w_013_374, w_009_222);
  not1 I013_376(w_013_376, w_007_419);
  and2 I013_379(w_013_379, w_006_251, w_011_463);
  and2 I013_380(w_013_380, w_001_009, w_009_096);
  not1 I013_382(w_013_382, w_005_267);
  not1 I013_385(w_013_385, w_011_397);
  or2  I013_386(w_013_386, w_000_205, w_010_000);
  or2  I013_391(w_013_391, w_007_295, w_006_221);
  not1 I013_392(w_013_392, w_001_008);
  nand2 I013_394(w_013_394, w_012_151, w_012_011);
  or2  I013_396(w_013_396, w_003_040, w_006_047);
  and2 I013_397(w_013_397, w_011_387, w_009_138);
  or2  I013_399(w_013_399, w_005_141, w_012_230);
  nand2 I013_400(w_013_400, w_011_136, w_005_135);
  not1 I013_401(w_013_401, w_006_017);
  or2  I013_403(w_013_403, w_007_464, w_006_054);
  and2 I013_404(w_013_404, w_003_035, w_001_003);
  nand2 I013_407(w_013_407, w_005_277, w_010_042);
  nand2 I013_408(w_013_408, w_004_059, w_007_076);
  not1 I013_409(w_013_409, w_012_315);
  nand2 I013_411(w_013_411, w_010_550, w_004_365);
  nand2 I013_412(w_013_412, w_002_039, w_004_061);
  not1 I013_413(w_013_413, w_002_069);
  not1 I013_414(w_013_414, w_004_198);
  not1 I013_415(w_013_415, w_006_213);
  and2 I013_416(w_013_416, w_002_304, w_008_168);
  not1 I013_418(w_013_418, w_010_611);
  and2 I013_419(w_013_419, w_000_025, w_000_238);
  not1 I013_422(w_013_422, w_004_161);
  and2 I013_426(w_013_426, w_007_040, w_011_503);
  nand2 I013_428(w_013_428, w_003_066, w_006_228);
  not1 I013_429(w_013_429, w_004_089);
  and2 I013_431(w_013_431, w_005_294, w_011_525);
  and2 I013_432(w_013_432, w_009_010, w_006_205);
  or2  I013_436(w_013_436, w_003_027, w_001_002);
  nand2 I013_437(w_013_437, w_001_032, w_010_429);
  nand2 I013_439(w_013_439, w_004_346, w_010_240);
  or2  I013_442(w_013_442, w_003_010, w_000_169);
  not1 I013_443(w_013_443, w_011_310);
  and2 I013_444(w_013_444, w_004_423, w_006_235);
  and2 I013_445(w_013_445, w_006_035, w_010_010);
  and2 I013_446(w_013_446, w_004_287, w_011_023);
  or2  I013_447(w_013_447, w_008_601, w_003_049);
  and2 I013_448(w_013_448, w_002_007, w_004_451);
  or2  I013_452(w_013_452, w_010_447, w_012_190);
  or2  I013_453(w_013_453, w_010_213, w_000_466);
  not1 I013_455(w_013_455, w_008_338);
  not1 I013_458(w_013_458, w_011_066);
  and2 I013_461(w_013_461, w_007_158, w_006_198);
  or2  I013_462(w_013_462, w_003_054, w_008_012);
  not1 I013_463(w_013_463, w_008_257);
  or2  I013_464(w_013_464, w_001_004, w_010_009);
  and2 I013_466(w_013_466, w_012_017, w_004_346);
  or2  I013_467(w_013_467, w_007_101, w_004_434);
  or2  I013_468(w_013_468, w_011_339, w_011_562);
  not1 I013_469(w_013_469, w_006_068);
  and2 I013_470(w_013_470, w_004_383, w_002_107);
  or2  I013_471(w_013_471, w_012_116, w_003_039);
  nand2 I013_478(w_013_478, w_008_215, w_002_251);
  not1 I013_479(w_013_479, w_007_160);
  not1 I013_484(w_013_484, w_008_062);
  not1 I013_489(w_013_489, w_006_115);
  not1 I013_494(w_013_494, w_004_172);
  and2 I013_496(w_013_496, w_003_031, w_004_046);
  nand2 I013_501(w_013_501, w_012_279, w_008_743);
  not1 I013_506(w_013_506, w_006_015);
  or2  I013_507(w_013_507, w_008_724, w_009_173);
  nand2 I013_509(w_013_509, w_006_219, w_007_211);
  not1 I013_510(w_013_510, w_006_101);
  nand2 I013_511(w_013_511, w_011_044, w_000_593);
  nand2 I013_514(w_013_514, w_008_019, w_010_002);
  and2 I013_515(w_013_515, w_010_614, w_001_026);
  not1 I013_517(w_013_517, w_009_016);
  not1 I013_518(w_013_518, w_011_439);
  or2  I013_519(w_013_519, w_010_519, w_006_227);
  not1 I013_520(w_013_520, w_009_406);
  or2  I013_521(w_013_521, w_000_149, w_008_331);
  not1 I013_522(w_013_522, w_011_235);
  or2  I013_523(w_013_523, w_012_132, w_002_210);
  or2  I013_524(w_013_524, w_002_417, w_008_333);
  nand2 I013_526(w_013_526, w_011_196, w_000_091);
  or2  I013_527(w_013_527, w_002_302, w_011_199);
  nand2 I013_528(w_013_528, w_000_348, w_001_007);
  not1 I013_529(w_013_529, w_001_020);
  nand2 I013_530(w_013_530, w_000_573, w_011_206);
  nand2 I013_534(w_013_534, w_011_037, w_010_117);
  nand2 I013_536(w_013_536, w_001_008, w_000_100);
  or2  I013_538(w_013_538, w_002_315, w_008_589);
  or2  I013_539(w_013_539, w_001_001, w_005_108);
  or2  I013_540(w_013_540, w_004_026, w_011_500);
  nand2 I013_541(w_013_541, w_012_078, w_002_416);
  and2 I013_542(w_013_542, w_009_169, w_005_004);
  not1 I013_543(w_013_543, w_003_048);
  and2 I013_544(w_013_544, w_011_010, w_009_110);
  and2 I013_545(w_013_545, w_006_193, w_012_309);
  nand2 I013_546(w_013_546, w_006_010, w_000_175);
  and2 I013_548(w_013_548, w_009_471, w_010_275);
  or2  I013_551(w_013_551, w_004_024, w_000_237);
  not1 I013_552(w_013_552, w_008_574);
  and2 I013_555(w_013_555, w_005_145, w_011_092);
  nand2 I013_556(w_013_556, w_000_494, w_008_414);
  or2  I013_558(w_013_558, w_002_265, w_004_484);
  nand2 I013_559(w_013_559, w_007_348, w_008_482);
  nand2 I013_560(w_013_560, w_009_062, w_011_615);
  or2  I013_561(w_013_561, w_003_004, w_004_280);
  nand2 I013_562(w_013_562, w_000_199, w_001_019);
  or2  I013_563(w_013_563, w_002_152, w_010_598);
  and2 I013_564(w_013_564, w_008_750, w_006_140);
  not1 I013_565(w_013_565, w_004_260);
  and2 I013_570(w_013_570, w_010_211, w_003_009);
  nand2 I013_571(w_013_571, w_009_082, w_008_033);
  and2 I013_572(w_013_572, w_008_433, w_000_494);
  nand2 I013_573(w_013_573, w_002_340, w_010_656);
  not1 I013_574(w_013_574, w_001_003);
  or2  I013_575(w_013_575, w_009_491, w_001_005);
  not1 I013_576(w_013_576, w_001_009);
  or2  I013_578(w_013_578, w_008_494, w_010_276);
  or2  I013_582(w_013_582, w_009_258, w_005_063);
  not1 I013_583(w_013_583, w_010_423);
  nand2 I013_584(w_013_586, w_013_585, w_003_044);
  not1 I013_585(w_013_587, w_013_586);
  and2 I013_586(w_013_588, w_013_587, w_010_181);
  and2 I013_587(w_013_589, w_013_588, w_009_168);
  and2 I013_588(w_013_590, w_013_589, w_012_002);
  nand2 I013_589(w_013_591, w_013_590, w_012_285);
  and2 I013_590(w_013_592, w_013_591, w_005_104);
  not1 I013_591(w_013_593, w_013_592);
  nand2 I013_592(w_013_594, w_013_593, w_005_242);
  nand2 I013_593(w_013_595, w_001_000, w_013_594);
  and2 I013_594(w_013_596, w_011_345, w_013_595);
  nand2 I013_595(w_013_585, w_013_596, w_003_067);
  not1 I014_000(w_014_000, w_007_300);
  or2  I014_001(w_014_001, w_002_176, w_007_276);
  and2 I014_002(w_014_002, w_000_193, w_010_291);
  nand2 I014_003(w_014_003, w_001_032, w_009_021);
  or2  I014_004(w_014_004, w_005_262, w_006_106);
  nand2 I014_005(w_014_005, w_008_337, w_010_013);
  not1 I014_007(w_014_007, w_000_172);
  not1 I014_008(w_014_008, w_005_000);
  not1 I014_009(w_014_009, w_005_194);
  not1 I014_010(w_014_010, w_010_289);
  nand2 I014_011(w_014_011, w_004_158, w_000_207);
  not1 I014_012(w_014_012, w_005_063);
  not1 I014_013(w_014_013, w_012_301);
  and2 I014_014(w_014_014, w_007_166, w_010_135);
  and2 I014_015(w_014_015, w_005_110, w_004_117);
  and2 I014_016(w_014_016, w_006_201, w_011_099);
  nand2 I014_017(w_014_017, w_001_000, w_007_060);
  nand2 I014_018(w_014_018, w_009_219, w_008_700);
  or2  I014_019(w_014_019, w_013_017, w_011_372);
  not1 I014_021(w_014_021, w_011_227);
  not1 I014_022(w_014_022, w_013_055);
  nand2 I014_023(w_014_023, w_003_061, w_002_223);
  or2  I014_024(w_014_024, w_003_043, w_008_029);
  not1 I014_025(w_014_025, w_004_056);
  and2 I014_026(w_014_026, w_012_072, w_006_206);
  nand2 I014_027(w_014_027, w_002_007, w_002_357);
  not1 I014_028(w_014_028, w_002_067);
  or2  I014_029(w_014_029, w_010_349, w_002_109);
  and2 I014_030(w_014_030, w_005_170, w_004_044);
  nand2 I014_031(w_014_031, w_005_158, w_004_391);
  nand2 I014_032(w_014_032, w_006_157, w_008_016);
  nand2 I014_034(w_014_034, w_002_261, w_001_018);
  and2 I014_035(w_014_035, w_004_269, w_005_146);
  and2 I014_036(w_014_036, w_008_315, w_010_194);
  or2  I014_037(w_014_037, w_006_084, w_012_350);
  and2 I014_039(w_014_039, w_007_152, w_005_176);
  and2 I014_040(w_014_040, w_000_498, w_013_046);
  nand2 I014_041(w_014_041, w_007_082, w_010_154);
  or2  I014_042(w_014_042, w_012_240, w_000_556);
  nand2 I014_043(w_014_043, w_000_154, w_013_232);
  and2 I014_044(w_014_044, w_010_670, w_004_104);
  and2 I014_045(w_014_045, w_007_032, w_012_147);
  nand2 I014_046(w_014_046, w_010_354, w_007_073);
  and2 I014_047(w_014_047, w_004_086, w_011_058);
  or2  I014_048(w_014_048, w_004_004, w_009_370);
  or2  I014_049(w_014_049, w_008_056, w_011_597);
  or2  I014_050(w_014_050, w_002_459, w_005_221);
  nand2 I014_052(w_014_052, w_005_286, w_000_357);
  not1 I014_053(w_014_053, w_008_461);
  or2  I014_054(w_014_054, w_003_010, w_006_119);
  and2 I014_055(w_014_055, w_001_030, w_009_164);
  and2 I014_056(w_014_056, w_005_123, w_007_429);
  or2  I014_057(w_014_057, w_013_169, w_011_569);
  nand2 I014_058(w_014_058, w_001_003, w_012_272);
  not1 I014_059(w_014_059, w_012_181);
  or2  I014_060(w_014_060, w_005_195, w_002_466);
  nand2 I014_061(w_014_061, w_008_644, w_011_583);
  and2 I014_062(w_014_062, w_005_109, w_002_022);
  and2 I014_064(w_014_064, w_007_280, w_001_017);
  not1 I014_066(w_014_066, w_011_189);
  or2  I014_067(w_014_067, w_013_208, w_006_154);
  and2 I014_068(w_014_068, w_001_005, w_000_208);
  not1 I014_069(w_014_069, w_002_142);
  nand2 I014_070(w_014_070, w_010_057, w_007_223);
  not1 I014_071(w_014_071, w_012_185);
  or2  I014_072(w_014_072, w_004_029, w_007_332);
  nand2 I014_073(w_014_073, w_004_100, w_004_195);
  nand2 I014_074(w_014_074, w_001_033, w_009_056);
  nand2 I014_075(w_014_075, w_009_428, w_003_035);
  not1 I014_076(w_014_076, w_004_410);
  or2  I014_077(w_014_077, w_012_116, w_002_200);
  or2  I014_080(w_014_080, w_001_019, w_007_204);
  nand2 I014_081(w_014_081, w_000_572, w_001_002);
  or2  I014_082(w_014_082, w_004_185, w_007_474);
  or2  I014_083(w_014_083, w_003_004, w_002_003);
  or2  I014_084(w_014_084, w_000_382, w_004_123);
  and2 I014_085(w_014_085, w_007_039, w_003_071);
  not1 I014_088(w_014_088, w_002_265);
  or2  I014_089(w_014_089, w_007_257, w_008_566);
  and2 I014_090(w_014_090, w_008_122, w_009_524);
  or2  I014_092(w_014_092, w_000_293, w_003_014);
  nand2 I014_093(w_014_093, w_013_183, w_000_028);
  or2  I014_094(w_014_094, w_007_237, w_009_117);
  and2 I014_095(w_014_095, w_004_158, w_007_378);
  nand2 I014_096(w_014_096, w_000_417, w_003_024);
  or2  I014_097(w_014_097, w_013_293, w_007_065);
  not1 I014_099(w_014_099, w_013_030);
  or2  I014_100(w_014_100, w_011_642, w_009_182);
  or2  I014_101(w_014_101, w_002_481, w_001_030);
  not1 I014_102(w_014_102, w_007_445);
  or2  I014_103(w_014_103, w_007_414, w_004_466);
  and2 I014_104(w_014_104, w_003_057, w_007_228);
  and2 I014_105(w_014_105, w_003_029, w_004_424);
  and2 I014_106(w_014_106, w_002_238, w_010_049);
  or2  I014_108(w_014_108, w_007_278, w_003_016);
  and2 I014_109(w_014_109, w_004_373, w_012_056);
  and2 I014_110(w_014_110, w_012_121, w_010_413);
  not1 I014_111(w_014_111, w_010_732);
  and2 I014_112(w_014_112, w_001_005, w_012_023);
  not1 I014_113(w_014_113, w_008_424);
  nand2 I014_114(w_014_114, w_011_208, w_009_555);
  not1 I014_115(w_014_115, w_002_033);
  or2  I014_116(w_014_116, w_001_013, w_002_310);
  and2 I014_117(w_014_117, w_008_702, w_000_586);
  nand2 I014_119(w_014_119, w_010_384, w_002_709);
  and2 I014_120(w_014_120, w_001_018, w_003_008);
  not1 I014_121(w_014_121, w_012_303);
  nand2 I014_122(w_014_122, w_013_096, w_008_475);
  or2  I014_123(w_014_123, w_009_154, w_005_231);
  and2 I014_124(w_014_124, w_012_134, w_011_190);
  and2 I014_125(w_014_125, w_001_012, w_001_022);
  not1 I014_126(w_014_126, w_001_005);
  not1 I014_127(w_014_127, w_002_320);
  not1 I014_129(w_014_129, w_005_136);
  not1 I014_130(w_014_130, w_012_303);
  nand2 I014_131(w_014_131, w_009_061, w_004_019);
  nand2 I014_132(w_014_132, w_012_017, w_007_333);
  nand2 I014_133(w_014_133, w_009_012, w_009_177);
  not1 I014_134(w_014_134, w_009_095);
  and2 I014_135(w_014_135, w_007_005, w_000_122);
  or2  I014_136(w_014_136, w_012_340, w_006_144);
  not1 I014_137(w_014_137, w_003_023);
  or2  I014_138(w_014_138, w_012_340, w_009_035);
  nand2 I014_140(w_014_140, w_003_084, w_006_099);
  and2 I014_141(w_014_141, w_011_295, w_004_410);
  and2 I014_142(w_014_142, w_009_415, w_008_269);
  and2 I014_143(w_014_143, w_007_161, w_007_171);
  nand2 I014_144(w_014_144, w_008_171, w_006_121);
  not1 I014_145(w_014_145, w_002_239);
  and2 I014_146(w_014_146, w_008_025, w_013_489);
  nand2 I014_147(w_014_147, w_003_039, w_013_220);
  not1 I014_148(w_014_148, w_001_002);
  not1 I014_149(w_014_149, w_009_598);
  not1 I014_150(w_014_150, w_004_111);
  or2  I014_151(w_014_151, w_004_048, w_007_097);
  and2 I014_152(w_014_152, w_012_219, w_012_020);
  not1 I014_153(w_014_153, w_003_001);
  nand2 I014_155(w_014_155, w_012_101, w_005_030);
  or2  I014_156(w_014_156, w_009_509, w_008_757);
  and2 I014_157(w_014_157, w_002_080, w_008_317);
  or2  I014_158(w_014_158, w_010_427, w_006_183);
  nand2 I014_159(w_014_159, w_003_048, w_003_082);
  and2 I014_160(w_014_160, w_005_145, w_008_150);
  and2 I014_161(w_014_161, w_005_138, w_007_166);
  or2  I014_162(w_014_162, w_006_144, w_010_626);
  nand2 I014_163(w_014_163, w_000_480, w_011_099);
  not1 I014_164(w_014_164, w_011_437);
  or2  I014_165(w_014_165, w_001_018, w_011_350);
  nand2 I014_166(w_014_166, w_012_324, w_003_080);
  not1 I014_167(w_014_167, w_011_024);
  not1 I014_168(w_014_168, w_000_643);
  nand2 I014_169(w_014_169, w_009_521, w_013_023);
  not1 I014_171(w_014_171, w_011_334);
  nand2 I014_172(w_014_172, w_012_311, w_002_128);
  and2 I014_173(w_014_173, w_007_181, w_005_106);
  nand2 I014_174(w_014_174, w_008_095, w_010_308);
  not1 I014_175(w_014_175, w_009_151);
  or2  I014_176(w_014_176, w_002_672, w_007_169);
  and2 I014_177(w_014_177, w_002_033, w_004_074);
  nand2 I014_178(w_014_178, w_013_408, w_012_003);
  and2 I014_179(w_014_179, w_001_033, w_002_118);
  or2  I014_180(w_014_180, w_007_061, w_006_004);
  nand2 I014_181(w_014_181, w_002_664, w_013_523);
  nand2 I014_182(w_014_182, w_006_098, w_010_705);
  not1 I014_183(w_014_183, w_010_348);
  and2 I014_184(w_014_184, w_012_071, w_013_369);
  nand2 I014_185(w_014_185, w_010_626, w_003_004);
  and2 I014_186(w_014_186, w_005_079, w_009_211);
  and2 I014_187(w_014_187, w_001_012, w_005_278);
  nand2 I014_188(w_014_188, w_002_321, w_000_523);
  and2 I014_189(w_014_189, w_010_428, w_003_010);
  and2 I014_190(w_014_190, w_005_305, w_009_626);
  or2  I014_191(w_014_191, w_002_056, w_004_031);
  nand2 I014_192(w_014_192, w_006_036, w_006_091);
  nand2 I014_193(w_014_193, w_001_012, w_010_596);
  nand2 I014_194(w_014_194, w_007_071, w_008_700);
  and2 I014_195(w_014_195, w_001_009, w_002_552);
  or2  I014_196(w_014_196, w_003_002, w_009_088);
  or2  I014_197(w_014_197, w_005_136, w_006_036);
  nand2 I014_198(w_014_198, w_011_131, w_005_215);
  nand2 I014_201(w_014_201, w_012_211, w_003_051);
  nand2 I014_202(w_014_202, w_010_698, w_006_242);
  not1 I014_203(w_014_203, w_013_371);
  or2  I014_205(w_014_205, w_004_325, w_009_011);
  and2 I014_206(w_014_206, w_003_027, w_011_576);
  and2 I014_209(w_014_209, w_003_027, w_004_165);
  or2  I014_210(w_014_210, w_002_088, w_011_575);
  not1 I014_211(w_014_211, w_010_014);
  nand2 I014_212(w_014_212, w_013_107, w_008_728);
  or2  I014_214(w_014_214, w_003_052, w_000_712);
  nand2 I014_215(w_014_215, w_009_445, w_002_078);
  and2 I014_216(w_014_216, w_004_085, w_004_052);
  nand2 I014_217(w_014_217, w_001_036, w_003_007);
  not1 I014_218(w_014_218, w_000_179);
  not1 I014_219(w_014_219, w_006_107);
  or2  I014_220(w_014_220, w_013_403, w_000_086);
  and2 I014_221(w_014_221, w_001_031, w_003_052);
  and2 I014_222(w_014_222, w_012_292, w_004_092);
  and2 I014_224(w_014_224, w_000_635, w_001_018);
  or2  I014_225(w_014_225, w_001_012, w_005_121);
  and2 I014_226(w_014_226, w_011_005, w_013_349);
  nand2 I014_228(w_014_228, w_005_068, w_005_139);
  and2 I014_229(w_014_229, w_007_259, w_012_106);
  not1 I014_231(w_014_231, w_009_021);
  and2 I014_233(w_014_233, w_011_020, w_007_067);
  and2 I014_234(w_014_234, w_003_047, w_012_026);
  not1 I014_235(w_014_235, w_003_008);
  or2  I014_236(w_014_236, w_004_102, w_002_671);
  and2 I014_237(w_014_237, w_002_113, w_009_374);
  nand2 I014_238(w_014_238, w_004_068, w_002_335);
  and2 I014_240(w_014_240, w_013_468, w_008_384);
  nand2 I014_241(w_014_241, w_006_158, w_000_319);
  and2 I014_242(w_014_242, w_007_249, w_002_688);
  and2 I014_243(w_014_243, w_000_598, w_013_200);
  and2 I014_245(w_014_245, w_011_228, w_005_289);
  nand2 I014_246(w_014_246, w_003_081, w_001_020);
  not1 I014_247(w_014_247, w_008_211);
  not1 I014_248(w_014_248, w_006_082);
  not1 I014_249(w_014_249, w_000_683);
  not1 I014_250(w_014_250, w_008_355);
  not1 I014_252(w_014_252, w_006_211);
  nand2 I014_253(w_014_253, w_005_036, w_013_538);
  not1 I014_254(w_014_254, w_004_027);
  nand2 I014_256(w_014_256, w_009_301, w_003_056);
  nand2 I014_257(w_014_257, w_001_018, w_005_065);
  nand2 I014_258(w_014_258, w_004_034, w_005_315);
  not1 I014_259(w_014_259, w_010_779);
  or2  I014_260(w_014_260, w_001_021, w_010_559);
  and2 I014_261(w_014_261, w_013_139, w_004_469);
  and2 I014_264(w_014_264, w_004_274, w_012_086);
  not1 I014_265(w_014_265, w_001_026);
  or2  I014_266(w_014_266, w_011_187, w_004_268);
  or2  I014_267(w_014_267, w_013_538, w_001_010);
  or2  I014_268(w_014_268, w_005_031, w_005_060);
  or2  I014_269(w_014_269, w_013_263, w_011_607);
  not1 I014_271(w_014_271, w_003_010);
  or2  I014_272(w_014_272, w_004_206, w_008_284);
  or2  I014_273(w_014_273, w_012_262, w_000_663);
  and2 I014_274(w_014_274, w_001_007, w_013_219);
  and2 I014_276(w_014_276, w_001_026, w_013_443);
  nand2 I014_277(w_014_277, w_004_453, w_012_039);
  or2  I014_279(w_014_279, w_010_157, w_010_748);
  or2  I014_280(w_014_280, w_008_348, w_004_150);
  nand2 I014_281(w_014_281, w_011_301, w_008_453);
  or2  I014_282(w_014_282, w_008_700, w_005_166);
  not1 I014_284(w_014_284, w_011_033);
  and2 I014_285(w_014_285, w_005_274, w_003_075);
  and2 I014_286(w_014_286, w_013_024, w_003_062);
  and2 I014_287(w_014_287, w_005_125, w_011_210);
  or2  I014_288(w_014_288, w_005_025, w_010_351);
  nand2 I014_289(w_014_289, w_001_019, w_000_296);
  and2 I014_290(w_014_290, w_000_550, w_007_132);
  and2 I014_291(w_014_291, w_013_047, w_006_156);
  not1 I014_292(w_014_292, w_012_082);
  not1 I014_294(w_014_294, w_005_149);
  or2  I014_295(w_014_295, w_007_283, w_008_085);
  nand2 I015_001(w_015_001, w_011_112, w_006_123);
  not1 I015_003(w_015_003, w_007_032);
  or2  I015_004(w_015_004, w_012_315, w_012_107);
  and2 I015_005(w_015_005, w_012_122, w_002_600);
  or2  I015_006(w_015_006, w_012_012, w_000_626);
  and2 I015_007(w_015_007, w_001_002, w_002_707);
  not1 I015_008(w_015_008, w_000_283);
  and2 I015_010(w_015_010, w_010_688, w_013_041);
  or2  I015_011(w_015_011, w_010_356, w_011_036);
  nand2 I015_013(w_015_013, w_013_506, w_000_272);
  not1 I015_014(w_015_014, w_001_015);
  not1 I015_015(w_015_015, w_005_130);
  or2  I015_016(w_015_016, w_011_308, w_002_471);
  and2 I015_017(w_015_017, w_004_359, w_008_192);
  or2  I015_019(w_015_019, w_007_349, w_012_162);
  and2 I015_020(w_015_020, w_002_571, w_005_240);
  and2 I015_022(w_015_022, w_011_368, w_002_677);
  and2 I015_023(w_015_023, w_012_348, w_004_161);
  nand2 I015_024(w_015_024, w_012_003, w_002_055);
  nand2 I015_026(w_015_026, w_009_166, w_011_542);
  not1 I015_027(w_015_027, w_009_301);
  and2 I015_029(w_015_029, w_009_259, w_003_041);
  nand2 I015_033(w_015_033, w_005_033, w_007_139);
  and2 I015_036(w_015_036, w_000_321, w_001_008);
  nand2 I015_038(w_015_038, w_007_224, w_005_123);
  and2 I015_040(w_015_040, w_009_031, w_012_281);
  or2  I015_041(w_015_041, w_006_212, w_007_007);
  nand2 I015_042(w_015_042, w_001_003, w_014_185);
  and2 I015_043(w_015_043, w_006_097, w_007_111);
  nand2 I015_044(w_015_044, w_006_054, w_011_164);
  not1 I015_045(w_015_045, w_014_130);
  nand2 I015_046(w_015_046, w_014_093, w_002_013);
  and2 I015_047(w_015_047, w_007_207, w_009_553);
  or2  I015_048(w_015_048, w_008_112, w_012_288);
  not1 I015_049(w_015_049, w_011_031);
  and2 I015_051(w_015_051, w_005_156, w_008_434);
  not1 I015_052(w_015_052, w_007_228);
  and2 I015_054(w_015_054, w_002_513, w_002_147);
  not1 I015_055(w_015_055, w_010_259);
  nand2 I015_056(w_015_056, w_005_186, w_005_036);
  or2  I015_057(w_015_057, w_000_351, w_008_637);
  and2 I015_058(w_015_058, w_005_026, w_011_605);
  nand2 I015_059(w_015_059, w_003_067, w_011_642);
  nand2 I015_060(w_015_060, w_000_148, w_004_099);
  or2  I015_061(w_015_061, w_006_247, w_008_658);
  not1 I015_062(w_015_062, w_003_063);
  or2  I015_065(w_015_065, w_012_273, w_013_095);
  or2  I015_067(w_015_067, w_010_526, w_005_118);
  or2  I015_068(w_015_068, w_006_017, w_013_025);
  nand2 I015_069(w_015_069, w_008_121, w_006_225);
  and2 I015_070(w_015_070, w_012_172, w_013_463);
  nand2 I015_071(w_015_071, w_000_297, w_006_212);
  or2  I015_072(w_015_072, w_008_640, w_004_224);
  not1 I015_073(w_015_073, w_014_196);
  nand2 I015_079(w_015_079, w_006_079, w_005_177);
  or2  I015_080(w_015_080, w_011_374, w_006_008);
  and2 I015_081(w_015_081, w_007_110, w_003_014);
  not1 I015_082(w_015_082, w_005_061);
  or2  I015_083(w_015_083, w_007_142, w_000_080);
  or2  I015_084(w_015_084, w_003_061, w_001_002);
  or2  I015_086(w_015_086, w_003_076, w_014_167);
  nand2 I015_087(w_015_087, w_010_335, w_002_400);
  nand2 I015_088(w_015_088, w_001_027, w_011_541);
  nand2 I015_089(w_015_089, w_001_006, w_005_005);
  not1 I015_090(w_015_090, w_012_275);
  and2 I015_091(w_015_091, w_000_484, w_011_138);
  not1 I015_092(w_015_092, w_001_024);
  and2 I015_093(w_015_093, w_012_262, w_014_153);
  nand2 I015_095(w_015_095, w_014_072, w_001_013);
  and2 I015_096(w_015_096, w_003_041, w_001_024);
  or2  I015_097(w_015_097, w_013_142, w_010_595);
  and2 I015_099(w_015_099, w_014_046, w_013_571);
  or2  I015_100(w_015_100, w_004_276, w_012_252);
  and2 I015_102(w_015_102, w_005_236, w_007_413);
  not1 I015_103(w_015_103, w_008_064);
  nand2 I015_104(w_015_104, w_013_206, w_009_383);
  and2 I015_105(w_015_105, w_000_220, w_010_467);
  nand2 I015_106(w_015_106, w_001_035, w_001_027);
  nand2 I015_107(w_015_107, w_005_196, w_003_065);
  not1 I015_108(w_015_108, w_000_051);
  not1 I015_110(w_015_110, w_006_202);
  not1 I015_111(w_015_111, w_002_221);
  not1 I015_112(w_015_112, w_007_304);
  or2  I015_113(w_015_113, w_011_073, w_014_188);
  and2 I015_114(w_015_114, w_013_179, w_013_081);
  nand2 I015_115(w_015_115, w_010_731, w_001_000);
  nand2 I015_116(w_015_116, w_013_049, w_005_224);
  nand2 I015_117(w_015_117, w_000_018, w_003_017);
  or2  I015_118(w_015_118, w_006_132, w_004_265);
  nand2 I015_119(w_015_119, w_005_077, w_002_491);
  nand2 I015_120(w_015_120, w_004_444, w_009_142);
  or2  I015_121(w_015_121, w_006_216, w_003_022);
  not1 I015_123(w_015_123, w_006_007);
  and2 I015_124(w_015_124, w_001_017, w_008_232);
  or2  I015_126(w_015_126, w_002_421, w_000_714);
  or2  I015_127(w_015_127, w_009_248, w_014_181);
  not1 I015_128(w_015_128, w_002_520);
  not1 I015_129(w_015_129, w_010_017);
  and2 I015_131(w_015_131, w_002_668, w_005_128);
  or2  I015_132(w_015_132, w_010_078, w_004_165);
  nand2 I015_133(w_015_133, w_013_002, w_012_273);
  nand2 I015_134(w_015_134, w_013_072, w_009_121);
  not1 I015_135(w_015_135, w_011_641);
  or2  I015_136(w_015_136, w_013_191, w_003_080);
  nand2 I015_137(w_015_137, w_004_409, w_008_078);
  nand2 I015_139(w_015_139, w_005_085, w_002_474);
  and2 I015_142(w_015_142, w_009_469, w_000_712);
  and2 I015_143(w_015_143, w_011_430, w_009_210);
  nand2 I015_144(w_015_144, w_003_045, w_004_158);
  not1 I015_146(w_015_146, w_003_006);
  and2 I015_149(w_015_149, w_002_125, w_001_022);
  or2  I015_151(w_015_151, w_004_163, w_007_189);
  not1 I015_152(w_015_152, w_008_012);
  nand2 I015_155(w_015_155, w_006_145, w_011_352);
  and2 I015_158(w_015_158, w_006_103, w_003_073);
  and2 I015_160(w_015_160, w_005_132, w_012_177);
  nand2 I015_161(w_015_161, w_012_048, w_008_371);
  or2  I015_162(w_015_162, w_004_213, w_012_088);
  nand2 I015_163(w_015_163, w_010_073, w_012_060);
  nand2 I015_164(w_015_164, w_014_246, w_011_028);
  nand2 I015_165(w_015_165, w_000_356, w_009_141);
  not1 I015_166(w_015_166, w_005_130);
  or2  I015_167(w_015_167, w_009_177, w_012_256);
  nand2 I015_168(w_015_168, w_013_530, w_006_031);
  not1 I015_170(w_015_170, w_013_316);
  not1 I015_172(w_015_172, w_010_286);
  or2  I015_174(w_015_174, w_005_068, w_009_479);
  not1 I015_177(w_015_177, w_002_040);
  nand2 I015_178(w_015_178, w_010_698, w_010_161);
  not1 I015_180(w_015_180, w_005_053);
  or2  I015_183(w_015_183, w_004_029, w_009_020);
  or2  I015_186(w_015_186, w_004_213, w_007_054);
  nand2 I015_187(w_015_187, w_013_218, w_002_566);
  or2  I015_188(w_015_188, w_014_143, w_002_078);
  and2 I015_190(w_015_190, w_002_193, w_010_283);
  not1 I015_191(w_015_191, w_000_715);
  not1 I015_192(w_015_192, w_000_716);
  nand2 I015_194(w_015_194, w_006_136, w_005_084);
  nand2 I015_196(w_015_196, w_003_042, w_009_510);
  not1 I015_197(w_015_197, w_003_023);
  and2 I015_198(w_015_198, w_006_172, w_002_163);
  and2 I015_200(w_015_200, w_012_000, w_014_039);
  or2  I015_201(w_015_201, w_005_107, w_013_108);
  not1 I015_202(w_015_202, w_010_114);
  nand2 I015_204(w_015_204, w_006_061, w_002_609);
  nand2 I015_205(w_015_205, w_004_263, w_012_219);
  nand2 I015_208(w_015_208, w_009_208, w_003_061);
  not1 I015_209(w_015_209, w_013_067);
  nand2 I015_210(w_015_210, w_003_019, w_008_304);
  or2  I015_212(w_015_212, w_013_416, w_003_072);
  and2 I015_214(w_015_214, w_009_579, w_010_757);
  not1 I015_215(w_015_215, w_005_165);
  nand2 I015_220(w_015_220, w_014_186, w_001_036);
  nand2 I015_222(w_015_222, w_004_128, w_006_004);
  not1 I015_223(w_015_223, w_000_108);
  nand2 I015_224(w_015_224, w_006_137, w_000_403);
  not1 I015_229(w_015_229, w_006_017);
  and2 I015_230(w_015_230, w_013_184, w_006_028);
  not1 I015_232(w_015_232, w_013_078);
  nand2 I015_234(w_015_234, w_012_264, w_001_027);
  and2 I015_235(w_015_235, w_011_416, w_005_139);
  not1 I015_236(w_015_236, w_003_053);
  and2 I015_240(w_015_240, w_001_025, w_010_136);
  not1 I015_246(w_015_246, w_008_314);
  nand2 I015_248(w_015_248, w_007_261, w_012_038);
  nand2 I015_249(w_015_249, w_014_039, w_014_101);
  and2 I015_252(w_015_252, w_003_081, w_008_526);
  nand2 I015_253(w_015_253, w_001_022, w_005_062);
  not1 I015_254(w_015_254, w_008_093);
  or2  I015_256(w_015_256, w_011_020, w_000_717);
  nand2 I015_257(w_015_257, w_000_706, w_005_307);
  nand2 I015_258(w_015_258, w_009_000, w_010_472);
  and2 I015_259(w_015_259, w_005_127, w_010_691);
  or2  I015_260(w_015_260, w_003_018, w_000_718);
  and2 I015_261(w_015_261, w_008_420, w_001_014);
  or2  I015_263(w_015_263, w_013_180, w_010_705);
  nand2 I015_265(w_015_265, w_013_496, w_002_011);
  and2 I015_266(w_015_266, w_012_054, w_005_313);
  nand2 I015_267(w_015_267, w_006_024, w_006_107);
  or2  I015_269(w_015_269, w_014_134, w_010_487);
  or2  I015_271(w_015_271, w_004_457, w_008_243);
  and2 I015_272(w_015_272, w_005_238, w_012_084);
  or2  I015_275(w_015_275, w_011_289, w_008_039);
  and2 I015_276(w_015_276, w_000_420, w_002_645);
  or2  I015_277(w_015_277, w_007_250, w_013_332);
  nand2 I015_278(w_015_278, w_006_118, w_000_088);
  nand2 I015_280(w_015_280, w_011_591, w_001_016);
  or2  I015_281(w_015_281, w_012_317, w_000_115);
  nand2 I015_283(w_015_283, w_000_120, w_007_016);
  nand2 I015_286(w_015_286, w_002_046, w_001_001);
  and2 I015_287(w_015_287, w_007_146, w_007_010);
  nand2 I015_288(w_015_288, w_011_201, w_003_002);
  not1 I015_290(w_015_290, w_010_353);
  nand2 I015_295(w_015_295, w_007_255, w_011_155);
  and2 I015_296(w_015_296, w_008_184, w_013_008);
  nand2 I015_299(w_015_299, w_003_059, w_003_039);
  or2  I015_301(w_015_301, w_005_186, w_011_322);
  or2  I015_302(w_015_302, w_007_321, w_008_093);
  and2 I015_308(w_015_308, w_000_117, w_009_143);
  not1 I015_309(w_015_309, w_008_646);
  not1 I015_314(w_015_314, w_014_158);
  nand2 I015_315(w_015_315, w_010_031, w_004_085);
  or2  I015_317(w_015_317, w_001_015, w_012_140);
  and2 I015_318(w_015_318, w_002_193, w_007_103);
  nand2 I015_319(w_015_319, w_010_482, w_009_357);
  or2  I015_322(w_015_322, w_007_057, w_003_041);
  and2 I015_323(w_015_323, w_009_472, w_009_581);
  not1 I015_325(w_015_325, w_007_131);
  or2  I015_328(w_015_328, w_013_046, w_003_082);
  and2 I015_332(w_015_332, w_007_356, w_003_002);
  not1 I015_333(w_015_333, w_014_142);
  and2 I015_335(w_015_335, w_005_162, w_002_363);
  not1 I015_336(w_015_336, w_005_214);
  and2 I015_339(w_015_339, w_002_690, w_009_336);
  and2 I015_340(w_015_340, w_000_272, w_000_240);
  nand2 I015_343(w_015_343, w_011_103, w_010_682);
  not1 I015_344(w_015_344, w_011_271);
  and2 I015_346(w_015_346, w_009_021, w_012_273);
  not1 I015_347(w_015_347, w_008_416);
  not1 I015_348(w_015_348, w_012_210);
  nand2 I015_351(w_015_351, w_011_490, w_004_226);
  nand2 I015_353(w_015_353, w_013_175, w_013_558);
  or2  I015_354(w_015_354, w_004_283, w_005_186);
  nand2 I015_355(w_015_355, w_011_197, w_011_014);
  and2 I015_357(w_015_357, w_002_518, w_008_018);
  or2  I015_360(w_015_360, w_008_117, w_012_088);
  or2  I015_363(w_015_363, w_008_338, w_010_358);
  not1 I015_366(w_015_366, w_004_008);
  and2 I015_369(w_015_369, w_001_000, w_010_013);
  nand2 I015_370(w_015_370, w_005_033, w_002_369);
  and2 I015_371(w_015_371, w_013_008, w_005_159);
  not1 I015_372(w_015_372, w_002_524);
  and2 I015_373(w_015_373, w_013_010, w_014_032);
  nand2 I015_374(w_015_374, w_014_106, w_002_386);
  nand2 I015_376(w_015_376, w_010_218, w_001_024);
  not1 I015_377(w_015_377, w_003_074);
  nand2 I015_379(w_015_379, w_010_080, w_000_720);
  not1 I015_382(w_015_382, w_012_200);
  or2  I015_384(w_015_384, w_011_020, w_013_305);
  or2  I015_385(w_015_385, w_014_226, w_004_209);
  nand2 I015_386(w_015_386, w_004_160, w_001_022);
  not1 I015_387(w_015_387, w_002_505);
  or2  I015_389(w_015_389, w_014_156, w_012_202);
  and2 I015_390(w_015_390, w_008_391, w_012_027);
  nand2 I015_392(w_015_392, w_002_309, w_006_019);
  and2 I015_393(w_015_393, w_010_003, w_010_249);
  not1 I015_394(w_015_394, w_004_307);
  nand2 I015_396(w_015_396, w_012_034, w_006_221);
  not1 I015_399(w_015_399, w_003_025);
  or2  I015_400(w_015_400, w_007_041, w_003_079);
  and2 I015_401(w_015_401, w_000_553, w_003_012);
  nand2 I015_402(w_015_402, w_008_603, w_009_111);
  and2 I015_405(w_015_405, w_011_196, w_006_026);
  not1 I015_407(w_015_407, w_011_520);
  not1 I015_408(w_015_408, w_011_273);
  and2 I015_413(w_015_413, w_012_092, w_011_406);
  and2 I015_416(w_015_416, w_009_272, w_006_143);
  or2  I015_417(w_015_417, w_009_038, w_005_146);
  and2 I015_418(w_015_418, w_010_219, w_007_059);
  not1 I015_421(w_015_421, w_014_291);
  and2 I015_423(w_015_423, w_006_048, w_002_013);
  and2 I015_426(w_015_426, w_003_009, w_012_255);
  or2  I015_428(w_015_428, w_014_122, w_013_307);
  or2  I015_429(w_015_429, w_013_176, w_004_362);
  or2  I015_430(w_015_430, w_011_391, w_000_688);
  not1 I015_431(w_015_431, w_012_252);
  or2  I015_432(w_015_432, w_005_004, w_005_290);
  not1 I015_433(w_015_433, w_003_012);
  nand2 I015_434(w_015_434, w_002_319, w_002_389);
  and2 I015_435(w_015_435, w_008_360, w_009_017);
  or2  I015_436(w_015_436, w_000_608, w_014_037);
  and2 I015_439(w_015_439, w_000_657, w_009_158);
  nand2 I015_440(w_015_440, w_004_255, w_008_738);
  not1 I015_441(w_015_441, w_002_328);
  nand2 I015_442(w_015_442, w_010_688, w_007_092);
  not1 I015_443(w_015_443, w_014_252);
  or2  I015_445(w_015_445, w_004_419, w_011_047);
  nand2 I015_447(w_015_447, w_008_292, w_005_106);
  nand2 I015_448(w_015_448, w_003_041, w_014_256);
  not1 I015_449(w_015_449, w_001_017);
  and2 I015_458(w_015_458, w_004_121, w_014_147);
  nand2 I015_459(w_015_459, w_013_016, w_008_662);
  nand2 I015_461(w_015_461, w_003_002, w_013_545);
  or2  I015_463(w_015_463, w_002_123, w_012_057);
  nand2 I015_464(w_015_464, w_008_244, w_011_489);
  or2  I015_467(w_015_467, w_001_026, w_003_081);
  nand2 I015_468(w_015_468, w_001_031, w_008_124);
  nand2 I015_469(w_015_469, w_005_146, w_003_042);
  nand2 I015_471(w_015_471, w_003_057, w_014_025);
  or2  I015_474(w_015_474, w_004_269, w_008_708);
  nand2 I015_476(w_015_476, w_003_007, w_012_088);
  or2  I015_477(w_015_477, w_014_209, w_002_201);
  nand2 I015_478(w_015_478, w_005_291, w_001_035);
  and2 I015_479(w_015_479, w_004_341, w_005_087);
  not1 I015_480(w_015_480, w_005_134);
  and2 I015_481(w_015_481, w_013_394, w_004_374);
  nand2 I015_484(w_015_484, w_001_010, w_005_133);
  nand2 I015_490(w_015_490, w_002_045, w_013_028);
  not1 I015_491(w_015_491, w_011_352);
  and2 I015_497(w_015_497, w_002_624, w_009_072);
  not1 I015_498(w_015_498, w_012_073);
  or2  I015_499(w_015_499, w_007_038, w_013_088);
  and2 I015_501(w_015_501, w_012_080, w_001_028);
  nand2 I015_502(w_015_502, w_002_510, w_009_293);
  or2  I015_504(w_015_504, w_005_018, w_007_437);
  not1 I015_506(w_015_506, w_012_247);
  nand2 I015_511(w_015_511, w_003_024, w_004_205);
  and2 I015_513(w_015_513, w_011_279, w_014_238);
  and2 I015_516(w_015_516, w_007_201, w_000_722);
  or2  I015_517(w_015_517, w_013_087, w_004_051);
  or2  I015_521(w_015_521, w_004_401, w_001_004);
  or2  I015_523(w_015_523, w_013_078, w_012_029);
  or2  I015_524(w_015_524, w_001_005, w_012_193);
  nand2 I015_526(w_015_526, w_007_079, w_004_070);
  not1 I015_527(w_015_527, w_009_026);
  not1 I015_529(w_015_529, w_005_066);
  nand2 I015_530(w_015_530, w_003_025, w_007_132);
  and2 I015_534(w_015_534, w_006_036, w_009_301);
  or2  I015_538(w_015_538, w_003_051, w_011_141);
  nand2 I015_543(w_015_543, w_010_265, w_002_436);
  and2 I015_544(w_015_544, w_011_538, w_002_056);
  not1 I015_546(w_015_546, w_002_116);
  or2  I015_547(w_015_547, w_009_100, w_010_450);
  and2 I015_548(w_015_548, w_001_006, w_005_129);
  not1 I015_550(w_015_550, w_014_101);
  and2 I015_552(w_015_552, w_008_499, w_012_001);
  or2  I015_555(w_015_555, w_011_343, w_011_205);
  not1 I015_556(w_015_556, w_005_019);
  or2  I015_557(w_015_557, w_010_288, w_011_155);
  nand2 I015_558(w_015_558, w_013_190, w_011_244);
  or2  I015_559(w_015_559, w_000_148, w_004_123);
  and2 I015_561(w_015_561, w_010_644, w_012_016);
  nand2 I015_562(w_015_562, w_000_124, w_011_170);
  and2 I015_565(w_015_565, w_001_009, w_007_321);
  not1 I015_566(w_015_566, w_003_031);
  and2 I015_568(w_015_568, w_005_317, w_012_138);
  or2  I015_570(w_015_570, w_004_437, w_002_083);
  nand2 I015_577(w_015_577, w_002_163, w_014_102);
  not1 I015_579(w_015_579, w_011_364);
  not1 I015_580(w_015_580, w_008_541);
  not1 I015_582(w_015_582, w_011_103);
  nand2 I015_584(w_015_584, w_010_193, w_014_245);
  and2 I015_585(w_015_585, w_001_021, w_011_133);
  or2  I015_589(w_015_589, w_007_184, w_012_008);
  or2  I015_590(w_015_590, w_009_441, w_002_368);
  not1 I015_591(w_015_591, w_007_036);
  nand2 I015_596(w_015_596, w_013_374, w_011_229);
  or2  I015_598(w_015_598, w_012_338, w_005_183);
  and2 I015_600(w_015_600, w_004_364, w_012_350);
  or2  I015_603(w_015_603, w_011_155, w_004_034);
  or2  I015_604(w_015_604, w_001_026, w_013_209);
  or2  I015_605(w_015_605, w_003_031, w_011_455);
  or2  I015_606(w_015_606, w_014_224, w_007_070);
  and2 I015_607(w_015_607, w_011_420, w_004_360);
  and2 I015_608(w_015_608, w_012_162, w_013_042);
  and2 I015_612(w_015_612, w_011_102, w_002_127);
  not1 I015_613(w_015_613, w_008_351);
  and2 I015_614(w_015_614, w_003_043, w_013_080);
  nand2 I015_615(w_015_615, w_005_058, w_007_166);
  and2 I015_616(w_015_616, w_011_131, w_000_505);
  not1 I015_618(w_015_618, w_014_235);
  not1 I015_619(w_015_619, w_011_180);
  or2  I015_620(w_015_620, w_008_032, w_009_021);
  and2 I015_624(w_015_624, w_002_511, w_011_419);
  nand2 I015_625(w_015_625, w_000_325, w_004_290);
  not1 I015_629(w_015_629, w_001_021);
  and2 I015_632(w_015_632, w_007_252, w_014_205);
  and2 I015_633(w_015_633, w_003_001, w_011_515);
  not1 I015_636(w_015_636, w_001_009);
  or2  I015_637(w_015_637, w_014_125, w_008_509);
  nand2 I015_641(w_015_641, w_001_013, w_010_596);
  or2  I015_642(w_015_642, w_010_362, w_008_619);
  nand2 I015_644(w_015_644, w_009_240, w_004_150);
  not1 I015_647(w_015_647, w_008_386);
  not1 I015_648(w_015_648, w_001_006);
  nand2 I015_649(w_015_649, w_003_017, w_009_507);
  or2  I015_650(w_015_650, w_014_168, w_004_410);
  nand2 I015_651(w_015_651, w_007_438, w_010_580);
  not1 I015_652(w_015_652, w_007_169);
  not1 I015_653(w_015_653, w_000_378);
  nand2 I015_654(w_015_654, w_002_041, w_012_327);
  not1 I015_658(w_015_658, w_005_303);
  not1 I015_660(w_015_660, w_014_076);
  and2 I015_662(w_015_662, w_010_482, w_008_030);
  not1 I015_663(w_015_663, w_005_213);
  and2 I015_664(w_015_664, w_007_240, w_007_389);
  and2 I015_665(w_015_665, w_012_045, w_011_087);
  nand2 I015_668(w_015_668, w_013_211, w_013_159);
  and2 I015_669(w_015_669, w_001_008, w_003_007);
  or2  I015_671(w_015_671, w_002_346, w_004_107);
  or2  I015_673(w_015_673, w_000_084, w_012_059);
  not1 I015_675(w_015_675, w_008_650);
  and2 I015_676(w_015_676, w_014_285, w_002_080);
  or2  I015_677(w_015_677, w_010_263, w_002_106);
  nand2 I016_000(w_016_000, w_003_075, w_014_175);
  and2 I016_001(w_016_001, w_004_335, w_005_153);
  nand2 I016_002(w_016_002, w_009_095, w_014_026);
  nand2 I016_003(w_016_003, w_013_518, w_010_343);
  not1 I016_004(w_016_004, w_009_125);
  and2 I016_005(w_016_005, w_009_442, w_007_064);
  and2 I016_006(w_016_006, w_001_000, w_012_260);
  nand2 I016_007(w_016_007, w_010_732, w_011_078);
  and2 I016_008(w_016_008, w_000_231, w_015_266);
  nand2 I017_001(w_017_001, w_016_000, w_008_382);
  nand2 I017_002(w_017_002, w_015_146, w_012_137);
  or2  I017_003(w_017_003, w_004_225, w_003_082);
  or2  I017_004(w_017_004, w_010_327, w_010_107);
  not1 I017_005(w_017_005, w_002_279);
  nand2 I017_006(w_017_006, w_004_326, w_001_035);
  and2 I017_007(w_017_007, w_009_032, w_005_047);
  not1 I017_008(w_017_008, w_013_429);
  or2  I017_009(w_017_009, w_011_576, w_002_081);
  or2  I017_010(w_017_010, w_006_219, w_008_005);
  nand2 I017_012(w_017_012, w_003_047, w_011_514);
  nand2 I017_013(w_017_013, w_012_027, w_010_514);
  not1 I017_014(w_017_014, w_007_079);
  and2 I017_015(w_017_015, w_003_032, w_007_129);
  not1 I017_016(w_017_016, w_000_122);
  and2 I017_017(w_017_017, w_007_211, w_002_693);
  not1 I017_018(w_017_018, w_003_056);
  not1 I017_019(w_017_019, w_009_065);
  nand2 I017_020(w_017_020, w_013_339, w_012_091);
  and2 I017_022(w_017_022, w_009_052, w_004_201);
  not1 I017_023(w_017_023, w_010_560);
  nand2 I017_024(w_017_024, w_000_235, w_010_186);
  nand2 I017_025(w_017_025, w_011_182, w_016_006);
  and2 I017_026(w_017_026, w_004_439, w_007_177);
  nand2 I017_027(w_017_027, w_012_199, w_004_044);
  and2 I017_028(w_017_028, w_015_033, w_007_121);
  or2  I017_029(w_017_029, w_011_066, w_010_533);
  not1 I017_030(w_017_030, w_007_261);
  or2  I017_031(w_017_031, w_008_129, w_013_129);
  nand2 I017_032(w_017_032, w_004_146, w_008_699);
  not1 I017_033(w_017_033, w_007_111);
  or2  I017_034(w_017_034, w_010_661, w_014_160);
  not1 I017_035(w_017_035, w_004_211);
  not1 I017_036(w_017_036, w_003_066);
  and2 I017_037(w_017_037, w_011_270, w_000_053);
  not1 I017_038(w_017_038, w_013_467);
  and2 I017_040(w_017_040, w_016_005, w_008_217);
  nand2 I017_042(w_017_042, w_003_041, w_003_070);
  or2  I017_043(w_017_043, w_006_055, w_007_269);
  not1 I017_045(w_017_045, w_009_539);
  not1 I017_047(w_017_047, w_002_206);
  not1 I017_048(w_017_048, w_006_063);
  and2 I017_050(w_017_050, w_000_724, w_015_649);
  nand2 I017_051(w_017_051, w_008_178, w_012_019);
  and2 I017_052(w_017_052, w_004_071, w_002_050);
  and2 I017_053(w_017_053, w_006_158, w_014_004);
  or2  I017_054(w_017_054, w_007_138, w_011_054);
  and2 I017_055(w_017_055, w_000_213, w_000_022);
  or2  I017_056(w_017_056, w_006_069, w_004_331);
  nand2 I017_057(w_017_057, w_007_186, w_001_014);
  and2 I017_059(w_017_059, w_001_005, w_008_059);
  and2 I017_060(w_017_060, w_000_550, w_007_469);
  and2 I017_063(w_017_063, w_015_026, w_001_007);
  and2 I017_064(w_017_064, w_014_161, w_009_629);
  or2  I017_065(w_017_065, w_001_001, w_009_543);
  or2  I017_066(w_017_066, w_003_062, w_000_692);
  nand2 I017_068(w_017_068, w_007_189, w_016_007);
  not1 I017_069(w_017_069, w_005_100);
  nand2 I017_070(w_017_070, w_004_126, w_001_028);
  not1 I017_071(w_017_071, w_007_227);
  or2  I017_072(w_017_072, w_002_566, w_013_096);
  and2 I017_073(w_017_073, w_004_477, w_016_008);
  nand2 I017_075(w_017_075, w_015_051, w_013_089);
  nand2 I017_078(w_017_078, w_007_166, w_013_444);
  and2 I017_080(w_017_080, w_000_378, w_009_504);
  not1 I017_082(w_017_082, w_002_384);
  or2  I017_085(w_017_085, w_010_012, w_016_005);
  nand2 I017_086(w_017_086, w_010_036, w_005_234);
  and2 I017_087(w_017_087, w_005_131, w_016_007);
  and2 I017_088(w_017_088, w_016_002, w_011_010);
  nand2 I017_089(w_017_089, w_013_237, w_006_246);
  not1 I017_091(w_017_091, w_009_215);
  and2 I017_092(w_017_092, w_011_561, w_010_368);
  and2 I017_093(w_017_093, w_004_246, w_016_001);
  and2 I017_094(w_017_094, w_005_089, w_007_158);
  or2  I017_095(w_017_095, w_015_121, w_004_181);
  and2 I017_096(w_017_096, w_001_031, w_001_011);
  or2  I017_097(w_017_097, w_011_603, w_010_633);
  nand2 I017_098(w_017_098, w_004_054, w_012_321);
  or2  I017_099(w_017_099, w_014_228, w_015_240);
  nand2 I017_100(w_017_100, w_007_396, w_011_599);
  and2 I017_101(w_017_101, w_005_127, w_002_624);
  or2  I017_102(w_017_102, w_006_037, w_003_023);
  or2  I017_103(w_017_103, w_011_270, w_009_189);
  and2 I017_104(w_017_104, w_015_413, w_009_215);
  and2 I017_107(w_017_107, w_005_208, w_015_301);
  and2 I017_108(w_017_108, w_008_126, w_002_012);
  or2  I017_111(w_017_111, w_010_145, w_008_161);
  and2 I017_112(w_017_112, w_006_002, w_006_193);
  nand2 I017_114(w_017_114, w_001_031, w_001_019);
  or2  I017_115(w_017_115, w_005_248, w_000_091);
  not1 I017_116(w_017_116, w_005_066);
  and2 I017_118(w_017_118, w_007_459, w_012_230);
  and2 I017_119(w_017_119, w_001_036, w_012_193);
  and2 I017_120(w_017_120, w_013_010, w_013_015);
  or2  I017_121(w_017_121, w_005_094, w_006_210);
  or2  I017_122(w_017_122, w_002_263, w_014_084);
  not1 I017_123(w_017_123, w_010_263);
  and2 I017_124(w_017_124, w_007_130, w_001_028);
  or2  I017_125(w_017_125, w_014_036, w_009_004);
  and2 I017_126(w_017_126, w_013_147, w_001_011);
  or2  I017_127(w_017_127, w_006_066, w_002_051);
  nand2 I017_128(w_017_128, w_016_004, w_002_679);
  and2 I017_130(w_017_130, w_009_095, w_002_073);
  nand2 I017_131(w_017_131, w_011_527, w_014_292);
  and2 I017_132(w_017_132, w_006_171, w_011_204);
  nand2 I017_133(w_017_133, w_013_156, w_012_030);
  nand2 I017_134(w_017_134, w_005_057, w_011_071);
  not1 I017_135(w_017_135, w_013_145);
  or2  I017_138(w_017_138, w_002_061, w_008_664);
  and2 I017_140(w_017_140, w_005_139, w_001_030);
  not1 I017_141(w_017_141, w_012_241);
  or2  I017_142(w_017_142, w_016_002, w_008_520);
  not1 I017_144(w_017_144, w_002_358);
  or2  I017_146(w_017_146, w_004_083, w_007_296);
  not1 I017_151(w_017_151, w_006_208);
  and2 I017_154(w_017_154, w_010_494, w_003_059);
  or2  I017_156(w_017_156, w_005_158, w_016_005);
  or2  I017_157(w_017_157, w_004_456, w_015_010);
  or2  I017_159(w_017_159, w_001_021, w_001_000);
  or2  I017_162(w_017_162, w_011_492, w_016_003);
  not1 I017_164(w_017_164, w_012_016);
  or2  I017_165(w_017_165, w_008_694, w_009_134);
  nand2 I017_166(w_017_166, w_002_575, w_008_659);
  nand2 I017_168(w_017_168, w_006_200, w_010_032);
  not1 I017_171(w_017_171, w_001_000);
  nand2 I017_174(w_017_174, w_002_209, w_016_006);
  and2 I017_176(w_017_176, w_002_683, w_008_043);
  nand2 I017_177(w_017_177, w_008_134, w_010_471);
  and2 I017_178(w_017_178, w_011_189, w_000_505);
  and2 I017_179(w_017_179, w_006_214, w_015_402);
  not1 I017_184(w_017_184, w_005_150);
  nand2 I017_186(w_017_186, w_002_042, w_008_473);
  or2  I017_187(w_017_187, w_010_313, w_001_007);
  not1 I017_189(w_017_189, w_016_004);
  nand2 I017_190(w_017_190, w_008_486, w_016_004);
  not1 I017_191(w_017_191, w_001_006);
  and2 I017_193(w_017_193, w_012_245, w_012_208);
  nand2 I017_194(w_017_194, w_014_224, w_011_347);
  or2  I017_197(w_017_197, w_003_073, w_003_036);
  not1 I017_200(w_017_200, w_004_279);
  or2  I017_201(w_017_201, w_001_025, w_016_004);
  nand2 I017_206(w_017_206, w_007_289, w_003_069);
  nand2 I017_207(w_017_207, w_008_580, w_005_044);
  or2  I017_211(w_017_211, w_000_252, w_009_492);
  or2  I017_214(w_017_214, w_014_237, w_000_447);
  and2 I017_215(w_017_215, w_012_290, w_008_334);
  and2 I017_218(w_017_218, w_014_085, w_014_072);
  and2 I017_222(w_017_222, w_009_214, w_014_289);
  not1 I017_224(w_017_224, w_011_633);
  not1 I017_226(w_017_226, w_012_061);
  or2  I017_227(w_017_227, w_013_028, w_006_125);
  nand2 I017_228(w_017_228, w_002_115, w_007_063);
  nand2 I017_229(w_017_229, w_004_011, w_011_557);
  or2  I017_232(w_017_232, w_004_022, w_013_288);
  and2 I017_234(w_017_234, w_004_063, w_009_366);
  not1 I017_235(w_017_235, w_002_033);
  or2  I017_236(w_017_236, w_006_162, w_008_709);
  nand2 I017_238(w_017_238, w_010_491, w_012_350);
  and2 I017_240(w_017_240, w_003_027, w_003_033);
  and2 I017_242(w_017_242, w_005_283, w_009_159);
  not1 I017_243(w_017_243, w_009_068);
  nand2 I017_245(w_017_245, w_005_076, w_005_218);
  not1 I017_246(w_017_246, w_003_079);
  or2  I017_247(w_017_247, w_016_007, w_007_004);
  not1 I017_248(w_017_248, w_016_006);
  or2  I017_249(w_017_249, w_008_085, w_003_077);
  and2 I017_251(w_017_251, w_013_561, w_011_096);
  and2 I017_252(w_017_252, w_016_005, w_012_295);
  not1 I017_256(w_017_256, w_014_185);
  not1 I017_257(w_017_257, w_011_082);
  not1 I017_258(w_017_258, w_012_007);
  or2  I017_260(w_017_260, w_011_480, w_012_096);
  or2  I017_262(w_017_262, w_010_686, w_012_000);
  and2 I017_263(w_017_263, w_006_089, w_011_491);
  and2 I017_264(w_017_264, w_013_573, w_008_674);
  or2  I017_267(w_017_267, w_009_084, w_007_420);
  not1 I017_269(w_017_269, w_015_080);
  nand2 I017_270(w_017_270, w_000_571, w_008_182);
  and2 I017_271(w_017_271, w_008_056, w_010_695);
  nand2 I017_272(w_017_272, w_000_636, w_002_157);
  and2 I017_274(w_017_274, w_013_442, w_009_274);
  nand2 I017_279(w_017_279, w_007_324, w_015_471);
  and2 I017_280(w_017_280, w_002_137, w_013_453);
  and2 I017_283(w_017_283, w_002_327, w_011_606);
  not1 I017_286(w_017_286, w_000_044);
  not1 I017_288(w_017_288, w_015_615);
  not1 I017_291(w_017_291, w_001_000);
  not1 I017_292(w_017_292, w_007_147);
  not1 I017_293(w_017_293, w_011_042);
  and2 I017_294(w_017_294, w_013_258, w_005_028);
  not1 I017_295(w_017_295, w_007_241);
  nand2 I017_297(w_017_297, w_015_618, w_012_346);
  not1 I017_298(w_017_298, w_003_063);
  nand2 I017_305(w_017_305, w_007_282, w_014_153);
  not1 I017_306(w_017_306, w_010_196);
  not1 I017_309(w_017_309, w_012_157);
  and2 I017_312(w_017_312, w_000_693, w_008_442);
  or2  I017_314(w_017_314, w_008_068, w_008_179);
  not1 I017_315(w_017_315, w_008_220);
  nand2 I017_318(w_017_318, w_015_498, w_013_202);
  nand2 I017_319(w_017_319, w_012_078, w_007_150);
  and2 I017_321(w_017_321, w_007_293, w_010_172);
  and2 I017_322(w_017_322, w_006_201, w_013_128);
  or2  I017_323(w_017_323, w_010_550, w_006_196);
  and2 I017_325(w_017_325, w_014_193, w_012_183);
  or2  I017_329(w_017_329, w_010_232, w_010_268);
  or2  I017_333(w_017_333, w_002_225, w_011_512);
  nand2 I017_336(w_017_336, w_011_156, w_014_276);
  and2 I017_337(w_017_337, w_008_143, w_010_278);
  and2 I017_338(w_017_338, w_001_022, w_003_063);
  nand2 I017_341(w_017_341, w_007_109, w_005_126);
  nand2 I017_343(w_017_343, w_013_164, w_000_068);
  not1 I017_344(w_017_344, w_016_008);
  and2 I017_345(w_017_345, w_002_159, w_014_040);
  nand2 I017_347(w_017_347, w_004_398, w_014_152);
  or2  I017_349(w_017_349, w_008_543, w_005_018);
  nand2 I017_352(w_017_352, w_012_027, w_011_365);
  nand2 I017_356(w_017_356, w_009_180, w_002_627);
  nand2 I017_357(w_017_357, w_016_005, w_000_057);
  nand2 I017_359(w_017_359, w_000_383, w_005_234);
  and2 I017_360(w_017_360, w_008_721, w_000_096);
  or2  I017_364(w_017_364, w_000_685, w_010_229);
  not1 I017_365(w_017_365, w_004_418);
  not1 I017_366(w_017_366, w_001_005);
  not1 I017_367(w_017_367, w_009_445);
  or2  I017_368(w_017_368, w_007_033, w_007_273);
  nand2 I017_370(w_017_370, w_009_080, w_000_727);
  and2 I017_371(w_017_371, w_008_180, w_014_105);
  or2  I017_372(w_017_372, w_011_142, w_005_305);
  and2 I017_373(w_017_373, w_006_094, w_014_032);
  and2 I017_374(w_017_374, w_009_536, w_011_050);
  or2  I017_375(w_017_375, w_015_022, w_007_037);
  or2  I017_376(w_017_376, w_000_239, w_001_036);
  not1 I017_379(w_017_379, w_000_728);
  or2  I017_380(w_017_380, w_005_296, w_006_066);
  and2 I017_381(w_017_381, w_000_017, w_012_324);
  nand2 I017_385(w_017_385, w_000_611, w_011_368);
  not1 I017_386(w_017_386, w_010_681);
  nand2 I017_390(w_017_390, w_010_133, w_013_524);
  and2 I017_392(w_017_392, w_015_471, w_016_004);
  nand2 I017_394(w_017_394, w_008_121, w_016_008);
  or2  I017_399(w_017_399, w_000_250, w_010_232);
  and2 I017_402(w_017_402, w_010_558, w_005_046);
  or2  I017_403(w_017_403, w_001_009, w_014_069);
  or2  I017_404(w_017_404, w_003_003, w_008_032);
  and2 I017_406(w_017_406, w_008_152, w_000_469);
  or2  I017_407(w_017_407, w_016_008, w_006_056);
  and2 I017_408(w_017_408, w_001_001, w_011_045);
  nand2 I017_409(w_017_409, w_006_229, w_008_107);
  not1 I017_410(w_017_410, w_004_308);
  or2  I017_412(w_017_412, w_016_001, w_003_008);
  and2 I017_415(w_017_415, w_006_144, w_009_054);
  or2  I017_416(w_017_416, w_000_514, w_013_284);
  and2 I017_419(w_017_419, w_002_150, w_012_082);
  or2  I017_421(w_017_421, w_008_510, w_014_177);
  nand2 I017_422(w_017_422, w_006_026, w_000_555);
  and2 I017_424(w_017_424, w_014_069, w_009_102);
  or2  I017_425(w_017_425, w_012_154, w_009_625);
  and2 I017_426(w_017_426, w_007_057, w_010_431);
  nand2 I017_428(w_017_428, w_012_108, w_002_491);
  not1 I017_429(w_017_429, w_002_047);
  not1 I017_430(w_017_430, w_015_479);
  nand2 I017_433(w_017_433, w_014_104, w_014_196);
  nand2 I017_434(w_017_434, w_008_072, w_013_205);
  or2  I017_435(w_017_435, w_000_612, w_008_186);
  nand2 I017_436(w_017_436, w_002_080, w_009_185);
  or2  I017_437(w_017_437, w_001_014, w_003_049);
  or2  I017_438(w_017_438, w_014_242, w_004_460);
  nand2 I017_439(w_017_439, w_003_024, w_011_332);
  or2  I017_443(w_017_443, w_008_471, w_009_614);
  or2  I017_447(w_017_447, w_008_038, w_006_015);
  or2  I017_449(w_017_449, w_015_132, w_000_175);
  or2  I017_451(w_017_451, w_008_053, w_001_005);
  not1 I017_453(w_017_453, w_001_008);
  or2  I017_458(w_017_458, w_005_114, w_006_238);
  nand2 I017_460(w_017_460, w_011_336, w_005_089);
  or2  I017_461(w_017_461, w_007_001, w_016_003);
  not1 I017_462(w_017_462, w_011_147);
  nand2 I017_463(w_017_463, w_005_255, w_008_721);
  not1 I017_464(w_017_464, w_004_316);
  or2  I017_467(w_017_467, w_015_222, w_002_710);
  not1 I017_468(w_017_468, w_014_243);
  or2  I017_470(w_017_470, w_016_006, w_003_031);
  or2  I017_471(w_017_471, w_014_023, w_007_213);
  or2  I017_475(w_017_475, w_007_165, w_010_080);
  and2 I017_477(w_017_477, w_008_299, w_012_226);
  not1 I017_479(w_017_479, w_012_001);
  and2 I017_480(w_017_480, w_007_186, w_005_115);
  or2  I017_482(w_017_482, w_006_252, w_001_022);
  nand2 I017_483(w_017_483, w_010_354, w_004_260);
  or2  I017_484(w_017_484, w_007_065, w_011_157);
  nand2 I017_485(w_017_485, w_015_197, w_014_047);
  nand2 I017_487(w_017_487, w_015_504, w_015_663);
  nand2 I017_492(w_017_492, w_001_026, w_009_133);
  or2  I017_495(w_017_495, w_015_167, w_000_421);
  and2 I017_496(w_017_496, w_015_089, w_005_160);
  nand2 I017_497(w_017_497, w_012_036, w_011_032);
  or2  I017_498(w_017_498, w_016_001, w_016_005);
  and2 I017_499(w_017_499, w_008_140, w_012_042);
  not1 I017_501(w_017_501, w_010_403);
  or2  I017_502(w_017_502, w_001_006, w_001_029);
  nand2 I017_506(w_017_506, w_000_401, w_001_026);
  not1 I017_508(w_017_508, w_000_162);
  not1 I017_512(w_017_512, w_004_029);
  not1 I017_513(w_017_513, w_012_080);
  nand2 I017_515(w_017_515, w_004_340, w_000_541);
  or2  I017_517(w_017_517, w_016_008, w_008_514);
  nand2 I017_518(w_017_518, w_011_566, w_013_409);
  nand2 I017_522(w_017_522, w_006_015, w_016_003);
  and2 I017_523(w_017_523, w_003_059, w_002_082);
  nand2 I017_524(w_017_524, w_010_149, w_008_099);
  nand2 I017_525(w_017_525, w_004_060, w_008_569);
  and2 I017_529(w_017_529, w_004_077, w_010_163);
  and2 I017_531(w_017_531, w_014_174, w_003_075);
  or2  I017_532(w_017_532, w_015_223, w_014_183);
  not1 I017_536(w_017_536, w_011_154);
  and2 I017_538(w_017_538, w_006_031, w_003_047);
  and2 I017_540(w_017_540, w_016_004, w_016_005);
  and2 I017_541(w_017_541, w_002_578, w_009_443);
  nand2 I017_543(w_017_543, w_016_001, w_009_120);
  not1 I017_546(w_017_546, w_001_007);
  nand2 I017_549(w_017_549, w_001_032, w_009_051);
  nand2 I017_552(w_017_552, w_005_233, w_015_196);
  nand2 I017_553(w_017_553, w_012_135, w_002_442);
  nand2 I017_555(w_017_555, w_000_731, w_013_382);
  and2 I017_559(w_017_559, w_016_002, w_003_057);
  nand2 I017_560(w_017_560, w_010_032, w_007_403);
  nand2 I017_561(w_017_561, w_010_529, w_011_148);
  nand2 I017_562(w_017_562, w_015_413, w_007_045);
  and2 I017_564(w_017_564, w_015_480, w_008_377);
  and2 I017_565(w_017_565, w_012_102, w_007_180);
  not1 I017_567(w_017_567, w_009_611);
  nand2 I017_569(w_017_569, w_009_019, w_013_302);
  nand2 I017_572(w_017_572, w_004_345, w_000_511);
  not1 I017_575(w_017_575, w_014_119);
  or2  I017_576(w_017_576, w_006_028, w_007_269);
  or2  I017_578(w_017_578, w_007_470, w_009_100);
  or2  I017_579(w_017_579, w_004_446, w_013_102);
  and2 I017_581(w_017_581, w_000_687, w_010_426);
  nand2 I017_587(w_017_587, w_010_365, w_001_017);
  and2 I017_589(w_017_589, w_014_177, w_005_049);
  not1 I017_590(w_017_590, w_002_664);
  or2  I017_591(w_017_591, w_009_091, w_010_403);
  not1 I017_592(w_017_592, w_000_186);
  not1 I017_594(w_017_594, w_016_006);
  not1 I017_596(w_017_596, w_005_311);
  or2  I017_597(w_017_597, w_015_071, w_004_308);
  nand2 I017_598(w_017_598, w_014_133, w_004_223);
  and2 I017_599(w_017_599, w_012_301, w_015_160);
  and2 I017_601(w_017_601, w_014_201, w_008_351);
  nand2 I017_603(w_017_603, w_011_134, w_007_342);
  and2 I017_606(w_017_606, w_016_002, w_015_550);
  or2  I017_607(w_017_607, w_016_008, w_011_001);
  or2  I017_609(w_017_609, w_003_083, w_012_061);
  and2 I017_611(w_017_611, w_012_059, w_000_537);
  not1 I017_612(w_017_612, w_005_108);
  not1 I017_613(w_017_613, w_004_171);
  nand2 I017_616(w_017_616, w_005_137, w_008_076);
  nand2 I017_620(w_017_620, w_008_017, w_003_003);
  or2  I017_623(w_017_623, w_009_564, w_015_530);
  not1 I017_625(w_017_625, w_005_227);
  nand2 I017_626(w_017_626, w_009_025, w_007_432);
  nand2 I017_629(w_017_629, w_016_006, w_015_065);
  and2 I017_631(w_017_631, w_005_263, w_016_004);
  or2  I017_636(w_017_636, w_013_066, w_007_289);
  and2 I017_639(w_017_639, w_007_234, w_005_223);
  or2  I017_640(w_017_640, w_004_013, w_003_064);
  not1 I017_648(w_017_648, w_009_176);
  or2  I017_649(w_017_649, w_012_063, w_014_100);
  nand2 I017_650(w_017_650, w_005_117, w_007_211);
  not1 I017_651(w_017_651, w_001_023);
  nand2 I017_653(w_017_653, w_014_093, w_014_104);
  or2  I017_655(w_017_655, w_003_024, w_016_004);
  and2 I017_657(w_017_657, w_003_034, w_014_121);
  and2 I017_659(w_017_659, w_008_198, w_000_035);
  not1 I017_660(w_017_660, w_012_078);
  or2  I017_662(w_017_662, w_014_076, w_014_171);
  not1 I017_663(w_017_663, w_002_673);
  not1 I017_664(w_017_664, w_013_003);
  nand2 I017_667(w_017_667, w_010_429, w_008_644);
  and2 I017_669(w_017_669, w_014_175, w_016_003);
  nand2 I017_670(w_017_670, w_000_691, w_014_041);
  nand2 I018_000(w_018_000, w_002_486, w_004_368);
  not1 I018_001(w_018_001, w_017_092);
  nand2 I018_002(w_018_002, w_005_270, w_004_213);
  not1 I018_003(w_018_003, w_007_434);
  not1 I018_004(w_018_004, w_006_090);
  not1 I018_005(w_018_005, w_016_003);
  and2 I018_006(w_018_006, w_003_002, w_001_002);
  not1 I018_007(w_018_007, w_009_191);
  and2 I018_008(w_018_008, w_004_020, w_006_249);
  and2 I018_009(w_018_009, w_013_049, w_015_636);
  nand2 I018_010(w_018_010, w_014_265, w_002_398);
  or2  I018_011(w_018_011, w_014_003, w_003_040);
  nand2 I018_012(w_018_012, w_000_188, w_003_042);
  not1 I018_013(w_018_013, w_003_022);
  and2 I018_014(w_018_014, w_010_179, w_014_012);
  nand2 I018_015(w_018_015, w_001_029, w_007_336);
  nand2 I018_016(w_018_016, w_002_172, w_002_086);
  not1 I018_017(w_018_017, w_004_484);
  nand2 I018_018(w_018_018, w_016_003, w_005_048);
  or2  I018_019(w_018_019, w_005_236, w_000_506);
  or2  I018_020(w_018_020, w_001_012, w_000_732);
  and2 I018_021(w_018_021, w_012_319, w_013_005);
  or2  I018_022(w_018_022, w_000_341, w_017_060);
  or2  I018_023(w_018_023, w_017_498, w_013_494);
  nand2 I018_024(w_018_024, w_017_650, w_002_058);
  or2  I018_025(w_018_025, w_017_639, w_014_053);
  or2  I018_026(w_018_026, w_006_215, w_006_079);
  or2  I018_027(w_018_027, w_011_390, w_016_008);
  and2 I018_028(w_018_028, w_004_161, w_015_093);
  or2  I018_029(w_018_029, w_001_019, w_004_002);
  and2 I018_030(w_018_030, w_015_405, w_003_035);
  nand2 I018_031(w_018_031, w_006_213, w_016_005);
  nand2 I018_032(w_018_032, w_009_223, w_012_055);
  nand2 I018_033(w_018_033, w_005_125, w_009_462);
  nand2 I018_034(w_018_034, w_017_596, w_016_008);
  nand2 I018_035(w_018_035, w_004_290, w_005_026);
  and2 I018_036(w_018_036, w_008_033, w_016_001);
  and2 I018_037(w_018_037, w_009_473, w_017_392);
  not1 I018_038(w_018_038, w_012_055);
  or2  I018_039(w_018_039, w_007_013, w_000_590);
  not1 I018_040(w_018_040, w_010_604);
  not1 I018_041(w_018_041, w_009_122);
  not1 I018_042(w_018_042, w_004_071);
  and2 I018_043(w_018_043, w_000_465, w_016_004);
  nand2 I018_044(w_018_044, w_001_036, w_006_166);
  or2  I019_000(w_019_000, w_005_212, w_015_590);
  and2 I019_001(w_019_001, w_012_116, w_008_666);
  or2  I019_002(w_019_002, w_016_008, w_008_538);
  nand2 I019_003(w_019_003, w_001_029, w_008_342);
  or2  I019_004(w_019_004, w_017_007, w_002_003);
  not1 I019_005(w_019_005, w_008_710);
  not1 I019_006(w_019_006, w_010_531);
  nand2 I019_007(w_019_007, w_015_295, w_005_148);
  nand2 I019_008(w_019_008, w_018_003, w_015_463);
  nand2 I019_009(w_019_009, w_009_455, w_009_267);
  not1 I019_010(w_019_010, w_010_199);
  and2 I019_011(w_019_011, w_010_432, w_018_003);
  and2 I019_012(w_019_012, w_000_082, w_013_293);
  and2 I019_013(w_019_013, w_004_024, w_010_210);
  nand2 I019_014(w_019_014, w_012_198, w_017_156);
  not1 I019_015(w_019_015, w_013_035);
  or2  I019_016(w_019_016, w_000_274, w_005_317);
  or2  I019_017(w_019_017, w_016_000, w_004_243);
  and2 I019_018(w_019_018, w_003_049, w_013_135);
  not1 I019_019(w_019_019, w_007_428);
  nand2 I019_020(w_019_020, w_011_004, w_012_108);
  not1 I020_000(w_020_000, w_008_662);
  nand2 I020_001(w_020_001, w_015_502, w_018_009);
  nand2 I020_002(w_020_002, w_013_035, w_019_002);
  or2  I020_003(w_020_003, w_007_125, w_012_219);
  and2 I020_004(w_020_004, w_016_002, w_015_155);
  not1 I020_005(w_020_005, w_015_662);
  nand2 I020_006(w_020_006, w_019_000, w_018_031);
  nand2 I020_007(w_020_007, w_019_002, w_014_257);
  nand2 I020_008(w_020_008, w_013_206, w_015_020);
  or2  I020_009(w_020_009, w_006_068, w_006_100);
  nand2 I020_010(w_020_010, w_019_019, w_007_427);
  nand2 I020_011(w_020_011, w_002_134, w_001_013);
  and2 I020_012(w_020_012, w_000_733, w_001_002);
  nand2 I020_013(w_020_013, w_009_422, w_016_000);
  not1 I020_015(w_020_015, w_016_008);
  not1 I020_016(w_020_016, w_014_201);
  or2  I020_018(w_020_018, w_013_050, w_016_001);
  and2 I020_019(w_020_019, w_005_157, w_008_386);
  or2  I020_020(w_020_020, w_019_003, w_018_021);
  or2  I020_021(w_020_021, w_002_101, w_000_734);
  and2 I020_022(w_020_022, w_019_018, w_008_624);
  nand2 I020_023(w_020_023, w_002_322, w_001_004);
  or2  I020_024(w_020_024, w_003_028, w_012_240);
  and2 I020_025(w_020_025, w_000_636, w_008_068);
  nand2 I020_027(w_020_027, w_016_006, w_008_230);
  nand2 I020_028(w_020_028, w_009_213, w_007_198);
  not1 I020_029(w_020_029, w_007_022);
  or2  I020_030(w_020_030, w_009_378, w_003_059);
  and2 I020_031(w_020_031, w_018_024, w_012_150);
  nand2 I020_032(w_020_032, w_012_338, w_015_232);
  and2 I020_033(w_020_033, w_005_252, w_011_102);
  not1 I020_034(w_020_034, w_000_332);
  or2  I020_035(w_020_035, w_001_023, w_012_313);
  nand2 I020_036(w_020_036, w_019_012, w_013_136);
  nand2 I020_037(w_020_037, w_008_042, w_007_378);
  and2 I020_038(w_020_038, w_019_016, w_015_051);
  and2 I020_039(w_020_039, w_003_041, w_012_068);
  not1 I020_042(w_020_042, w_016_004);
  nand2 I020_043(w_020_043, w_009_267, w_002_097);
  or2  I020_044(w_020_044, w_010_027, w_017_269);
  not1 I020_045(w_020_045, w_005_035);
  not1 I020_049(w_020_049, w_011_462);
  not1 I020_050(w_020_050, w_009_265);
  nand2 I020_051(w_020_051, w_008_367, w_004_039);
  nand2 I020_054(w_020_054, w_000_735, w_018_019);
  not1 I020_055(w_020_055, w_005_137);
  or2  I020_057(w_020_057, w_015_654, w_018_000);
  not1 I020_058(w_020_058, w_007_237);
  not1 I020_059(w_020_059, w_008_669);
  or2  I020_062(w_020_062, w_002_188, w_011_372);
  nand2 I020_063(w_020_063, w_014_217, w_017_040);
  not1 I020_064(w_020_064, w_017_029);
  or2  I020_065(w_020_065, w_003_014, w_009_065);
  nand2 I020_067(w_020_067, w_010_638, w_006_158);
  or2  I020_068(w_020_068, w_010_338, w_005_059);
  nand2 I020_069(w_020_069, w_019_017, w_010_312);
  and2 I020_071(w_020_071, w_003_020, w_013_206);
  or2  I020_072(w_020_072, w_015_272, w_015_010);
  and2 I020_074(w_020_074, w_011_631, w_006_170);
  and2 I020_075(w_020_075, w_005_168, w_006_069);
  and2 I020_076(w_020_076, w_015_152, w_013_121);
  and2 I020_077(w_020_077, w_009_264, w_006_243);
  not1 I020_078(w_020_078, w_003_050);
  not1 I020_080(w_020_080, w_013_128);
  nand2 I020_083(w_020_083, w_012_192, w_014_164);
  not1 I020_084(w_020_084, w_006_025);
  not1 I020_086(w_020_086, w_018_003);
  and2 I020_087(w_020_087, w_004_178, w_014_222);
  nand2 I020_088(w_020_088, w_002_283, w_005_038);
  nand2 I020_090(w_020_090, w_008_499, w_006_127);
  not1 I020_091(w_020_091, w_012_111);
  or2  I020_092(w_020_092, w_011_330, w_005_137);
  nand2 I020_094(w_020_094, w_004_238, w_006_198);
  not1 I020_095(w_020_095, w_012_237);
  or2  I020_096(w_020_096, w_002_069, w_001_034);
  and2 I020_098(w_020_098, w_003_066, w_009_045);
  and2 I020_099(w_020_099, w_006_177, w_013_121);
  and2 I020_100(w_020_100, w_003_046, w_015_067);
  not1 I020_102(w_020_102, w_015_070);
  and2 I020_103(w_020_103, w_016_008, w_001_001);
  nand2 I020_105(w_020_105, w_010_510, w_008_248);
  not1 I020_107(w_020_107, w_016_005);
  or2  I020_108(w_020_108, w_003_036, w_014_224);
  and2 I020_109(w_020_109, w_000_575, w_011_120);
  nand2 I020_110(w_020_110, w_007_398, w_016_007);
  nand2 I020_114(w_020_114, w_011_244, w_005_247);
  or2  I020_115(w_020_115, w_001_016, w_005_192);
  not1 I020_116(w_020_116, w_000_440);
  or2  I020_118(w_020_118, w_011_209, w_000_544);
  and2 I020_119(w_020_119, w_011_586, w_008_356);
  nand2 I020_122(w_020_122, w_008_394, w_016_001);
  and2 I020_123(w_020_123, w_016_002, w_009_103);
  nand2 I020_124(w_020_124, w_008_131, w_012_328);
  and2 I020_125(w_020_125, w_005_105, w_016_003);
  not1 I020_126(w_020_126, w_005_105);
  or2  I020_129(w_020_129, w_018_035, w_010_554);
  and2 I020_130(w_020_130, w_019_019, w_015_387);
  nand2 I020_131(w_020_131, w_007_137, w_003_002);
  nand2 I020_132(w_020_132, w_000_581, w_017_625);
  nand2 I020_134(w_020_134, w_010_322, w_010_280);
  and2 I020_135(w_020_135, w_008_218, w_003_008);
  and2 I020_136(w_020_136, w_003_019, w_016_000);
  not1 I020_138(w_020_138, w_002_031);
  nand2 I020_139(w_020_139, w_000_120, w_001_026);
  or2  I020_140(w_020_140, w_012_143, w_000_736);
  not1 I020_142(w_020_142, w_011_384);
  or2  I020_144(w_020_144, w_010_177, w_004_038);
  and2 I020_146(w_020_146, w_006_222, w_000_638);
  or2  I020_147(w_020_147, w_015_091, w_005_198);
  and2 I020_148(w_020_148, w_007_086, w_015_413);
  nand2 I020_149(w_020_149, w_006_038, w_005_009);
  nand2 I020_151(w_020_151, w_003_001, w_005_026);
  or2  I020_152(w_020_152, w_006_039, w_001_006);
  nand2 I020_153(w_020_153, w_014_001, w_007_319);
  and2 I020_154(w_020_154, w_011_566, w_000_486);
  nand2 I020_155(w_020_155, w_015_164, w_008_312);
  or2  I020_157(w_020_157, w_011_127, w_014_209);
  or2  I020_158(w_020_158, w_007_293, w_010_680);
  or2  I020_160(w_020_160, w_019_018, w_011_251);
  not1 I020_161(w_020_161, w_002_179);
  not1 I020_162(w_020_162, w_010_491);
  or2  I020_163(w_020_163, w_007_132, w_001_028);
  and2 I020_164(w_020_164, w_004_266, w_018_013);
  and2 I020_165(w_020_165, w_017_037, w_014_083);
  not1 I020_166(w_020_166, w_000_163);
  or2  I020_167(w_020_167, w_005_097, w_000_289);
  or2  I020_169(w_020_169, w_011_414, w_018_025);
  and2 I020_170(w_020_170, w_019_004, w_012_016);
  and2 I020_171(w_020_171, w_010_749, w_012_288);
  not1 I020_172(w_020_172, w_007_034);
  and2 I020_173(w_020_173, w_019_007, w_005_085);
  not1 I020_175(w_020_175, w_007_359);
  or2  I020_177(w_020_177, w_017_123, w_006_225);
  or2  I020_179(w_020_179, w_015_256, w_009_024);
  and2 I020_180(w_020_180, w_014_291, w_015_431);
  not1 I020_181(w_020_181, w_002_419);
  nand2 I020_183(w_020_183, w_005_026, w_017_024);
  and2 I020_184(w_020_184, w_015_120, w_003_038);
  and2 I020_186(w_020_186, w_001_004, w_008_747);
  not1 I020_188(w_020_188, w_002_011);
  and2 I020_189(w_020_189, w_002_003, w_004_047);
  nand2 I020_192(w_020_192, w_015_001, w_007_126);
  not1 I020_193(w_020_193, w_015_108);
  not1 I020_196(w_020_196, w_009_489);
  not1 I020_198(w_020_198, w_010_751);
  or2  I020_199(w_020_199, w_013_565, w_012_301);
  or2  I020_203(w_020_203, w_008_521, w_007_074);
  and2 I020_205(w_020_205, w_004_184, w_018_027);
  not1 I020_208(w_020_208, w_019_001);
  nand2 I020_209(w_020_209, w_019_011, w_012_115);
  and2 I020_210(w_020_210, w_012_188, w_007_438);
  and2 I020_216(w_020_216, w_003_012, w_008_518);
  or2  I020_217(w_020_217, w_012_004, w_016_003);
  and2 I020_221(w_020_221, w_006_248, w_013_290);
  nand2 I020_225(w_020_225, w_011_092, w_003_075);
  not1 I020_226(w_020_226, w_006_169);
  and2 I020_230(w_020_230, w_018_017, w_017_063);
  or2  I020_232(w_020_232, w_004_425, w_012_261);
  not1 I020_236(w_020_236, w_010_283);
  nand2 I020_240(w_020_240, w_010_091, w_002_598);
  not1 I020_244(w_020_244, w_006_021);
  and2 I020_246(w_020_246, w_017_197, w_019_002);
  and2 I020_247(w_020_247, w_014_157, w_001_027);
  nand2 I020_248(w_020_248, w_002_102, w_007_140);
  or2  I020_250(w_020_250, w_008_153, w_007_047);
  and2 I020_251(w_020_251, w_004_136, w_009_163);
  and2 I020_252(w_020_252, w_017_343, w_014_132);
  not1 I020_255(w_020_255, w_006_059);
  not1 I020_257(w_020_257, w_005_031);
  or2  I020_259(w_020_259, w_015_379, w_003_005);
  or2  I020_260(w_020_260, w_012_333, w_000_067);
  not1 I020_264(w_020_264, w_018_009);
  and2 I020_266(w_020_266, w_008_020, w_003_053);
  and2 I020_267(w_020_267, w_015_363, w_016_001);
  not1 I020_269(w_020_269, w_011_411);
  nand2 I020_271(w_020_271, w_005_123, w_001_021);
  nand2 I020_272(w_020_272, w_002_368, w_007_168);
  nand2 I020_277(w_020_277, w_007_046, w_014_082);
  nand2 I020_278(w_020_278, w_016_005, w_002_027);
  not1 I020_280(w_020_280, w_006_070);
  and2 I020_281(w_020_281, w_004_242, w_005_247);
  or2  I020_283(w_020_283, w_017_467, w_018_014);
  and2 I020_285(w_020_285, w_019_004, w_000_339);
  not1 I020_287(w_020_287, w_005_254);
  and2 I020_288(w_020_288, w_007_039, w_005_201);
  nand2 I020_290(w_020_290, w_006_076, w_001_000);
  nand2 I020_291(w_020_291, w_018_022, w_016_008);
  nand2 I020_296(w_020_296, w_002_291, w_007_009);
  and2 I020_297(w_020_297, w_008_694, w_004_167);
  and2 I020_300(w_020_300, w_009_480, w_013_519);
  nand2 I020_301(w_020_301, w_014_044, w_004_400);
  not1 I020_305(w_020_305, w_004_321);
  not1 I020_306(w_020_306, w_013_132);
  not1 I020_307(w_020_307, w_011_128);
  and2 I020_309(w_020_309, w_002_343, w_005_100);
  or2  I020_311(w_020_311, w_006_192, w_019_000);
  nand2 I020_314(w_020_314, w_003_066, w_002_004);
  not1 I020_315(w_020_315, w_018_003);
  or2  I020_319(w_020_319, w_015_248, w_009_549);
  nand2 I020_320(w_020_320, w_012_244, w_010_216);
  or2  I020_322(w_020_322, w_010_633, w_011_635);
  or2  I020_327(w_020_327, w_009_412, w_004_495);
  or2  I020_329(w_020_329, w_004_299, w_006_202);
  nand2 I020_331(w_020_331, w_013_098, w_019_014);
  nand2 I020_334(w_020_334, w_004_099, w_004_152);
  and2 I020_335(w_020_335, w_001_030, w_019_019);
  not1 I020_339(w_020_339, w_007_207);
  not1 I020_340(w_020_340, w_005_047);
  not1 I020_341(w_020_341, w_008_573);
  nand2 I020_342(w_020_342, w_007_088, w_017_007);
  and2 I020_347(w_020_347, w_000_404, w_010_568);
  not1 I020_348(w_020_348, w_005_168);
  not1 I020_350(w_020_350, w_007_407);
  not1 I020_355(w_020_355, w_000_092);
  not1 I020_356(w_020_356, w_010_610);
  and2 I020_359(w_020_359, w_012_076, w_018_036);
  nand2 I020_361(w_020_361, w_008_493, w_009_080);
  and2 I020_363(w_020_363, w_015_258, w_005_309);
  and2 I020_364(w_020_364, w_015_212, w_010_587);
  or2  I020_370(w_020_370, w_001_014, w_002_411);
  or2  I020_372(w_020_372, w_018_027, w_015_080);
  not1 I020_374(w_020_374, w_015_052);
  nand2 I020_378(w_020_378, w_013_070, w_012_001);
  or2  I020_379(w_020_379, w_000_661, w_016_007);
  not1 I020_380(w_020_380, w_005_092);
  and2 I020_381(w_020_381, w_000_738, w_004_102);
  nand2 I020_383(w_020_383, w_013_307, w_010_565);
  nand2 I020_386(w_020_386, w_001_023, w_001_001);
  nand2 I020_387(w_020_387, w_006_118, w_009_022);
  not1 I020_389(w_020_389, w_015_668);
  not1 I020_391(w_020_391, w_019_001);
  and2 I020_393(w_020_393, w_001_002, w_009_598);
  nand2 I020_394(w_020_394, w_000_585, w_013_091);
  not1 I020_395(w_020_395, w_016_000);
  or2  I020_396(w_020_396, w_000_144, w_012_299);
  nand2 I020_398(w_020_398, w_008_009, w_012_214);
  or2  I020_399(w_020_399, w_002_236, w_009_383);
  not1 I020_400(w_020_400, w_011_181);
  not1 I020_403(w_020_403, w_008_079);
  not1 I020_404(w_020_404, w_019_007);
  and2 I020_406(w_020_406, w_011_407, w_006_242);
  or2  I020_407(w_020_407, w_007_337, w_013_128);
  or2  I020_408(w_020_408, w_004_231, w_014_290);
  not1 I020_409(w_020_409, w_013_009);
  and2 I020_410(w_020_410, w_006_124, w_015_568);
  or2  I020_411(w_020_411, w_014_234, w_016_007);
  and2 I020_412(w_020_412, w_012_025, w_017_523);
  and2 I020_416(w_020_416, w_008_621, w_001_036);
  not1 I020_417(w_020_417, w_008_526);
  not1 I020_420(w_020_420, w_017_501);
  or2  I020_423(w_020_423, w_018_007, w_018_032);
  not1 I020_425(w_020_425, w_019_016);
  or2  I020_426(w_020_426, w_001_016, w_009_360);
  not1 I020_427(w_020_427, w_011_466);
  nand2 I020_428(w_020_428, w_004_184, w_014_151);
  or2  I020_429(w_020_429, w_000_039, w_019_019);
  or2  I020_430(w_020_430, w_018_012, w_007_100);
  and2 I020_433(w_020_433, w_002_522, w_013_534);
  not1 I020_436(w_020_436, w_009_570);
  not1 I020_438(w_020_438, w_009_139);
  or2  I020_441(w_020_441, w_017_224, w_014_153);
  or2  I020_442(w_020_442, w_001_011, w_010_088);
  or2  I020_445(w_020_445, w_019_016, w_017_323);
  nand2 I020_446(w_020_446, w_005_262, w_008_678);
  not1 I020_447(w_020_447, w_001_029);
  nand2 I020_448(w_020_448, w_007_198, w_012_277);
  nand2 I020_450(w_020_450, w_000_404, w_011_540);
  and2 I020_451(w_020_451, w_006_121, w_009_037);
  nand2 I020_452(w_020_452, w_006_108, w_006_143);
  nand2 I020_453(w_020_453, w_014_021, w_001_033);
  and2 I020_455(w_020_455, w_009_451, w_012_275);
  nand2 I020_457(w_020_457, w_009_023, w_009_108);
  or2  I020_460(w_020_460, w_013_517, w_000_583);
  or2  I020_461(w_020_461, w_004_223, w_004_129);
  and2 I020_462(w_020_462, w_001_030, w_016_004);
  nand2 I020_463(w_020_463, w_011_032, w_005_201);
  nand2 I020_465(w_020_465, w_019_016, w_008_411);
  nand2 I020_466(w_020_466, w_013_092, w_008_273);
  and2 I020_472(w_020_472, w_014_096, w_009_435);
  nand2 I020_473(w_020_473, w_001_033, w_005_219);
  nand2 I020_474(w_020_474, w_016_001, w_003_005);
  or2  I020_475(w_020_475, w_006_081, w_014_077);
  nand2 I020_476(w_020_476, w_011_544, w_011_273);
  or2  I020_479(w_020_479, w_013_303, w_005_086);
  not1 I020_482(w_020_482, w_002_084);
  or2  I020_483(w_020_483, w_006_122, w_000_339);
  nand2 I020_484(w_020_484, w_019_013, w_014_156);
  nand2 I020_489(w_020_489, w_019_002, w_011_131);
  or2  I020_490(w_020_490, w_006_070, w_007_151);
  and2 I020_494(w_020_494, w_011_118, w_016_001);
  or2  I020_495(w_020_495, w_019_005, w_008_090);
  and2 I020_498(w_020_498, w_004_024, w_005_062);
  nand2 I020_500(w_020_500, w_008_535, w_011_431);
  or2  I020_501(w_020_501, w_007_127, w_002_586);
  and2 I020_502(w_020_502, w_010_677, w_018_042);
  not1 I020_506(w_020_506, w_002_329);
  nand2 I020_508(w_020_508, w_013_331, w_015_616);
  or2  I020_511(w_020_511, w_014_148, w_002_455);
  and2 I020_512(w_020_512, w_001_019, w_019_017);
  and2 I020_513(w_020_513, w_002_451, w_002_119);
  nand2 I020_514(w_020_514, w_013_080, w_003_038);
  and2 I020_515(w_020_515, w_018_026, w_000_324);
  and2 I020_516(w_020_516, w_004_027, w_006_035);
  nand2 I020_517(w_020_517, w_011_309, w_008_426);
  and2 I020_518(w_020_518, w_004_367, w_015_136);
  not1 I020_519(w_020_519, w_003_000);
  or2  I020_520(w_020_520, w_005_289, w_017_590);
  not1 I020_521(w_020_521, w_000_181);
  or2  I020_525(w_020_525, w_007_314, w_015_648);
  and2 I020_527(w_020_527, w_001_019, w_010_747);
  and2 I020_529(w_020_529, w_011_032, w_006_011);
  not1 I020_530(w_020_530, w_013_334);
  not1 I020_536(w_020_536, w_005_169);
  not1 I020_539(w_020_539, w_018_025);
  or2  I020_543(w_020_543, w_010_352, w_007_118);
  or2  I020_545(w_020_545, w_019_008, w_008_381);
  not1 I020_546(w_020_546, w_018_003);
  not1 I020_547(w_020_547, w_003_042);
  and2 I020_549(w_020_549, w_010_769, w_012_124);
  nand2 I020_550(w_020_550, w_014_082, w_010_452);
  and2 I020_551(w_020_551, w_000_498, w_019_005);
  and2 I020_554(w_020_554, w_016_008, w_003_074);
  nand2 I020_561(w_020_561, w_004_338, w_012_027);
  or2  I020_562(w_020_562, w_008_346, w_006_130);
  or2  I020_564(w_020_564, w_000_230, w_004_037);
  or2  I020_565(w_020_565, w_019_017, w_007_056);
  nand2 I020_568(w_020_568, w_016_007, w_001_023);
  and2 I020_569(w_020_569, w_018_014, w_009_155);
  and2 I020_571(w_020_571, w_010_444, w_014_075);
  and2 I020_576(w_020_576, w_007_224, w_010_321);
  nand2 I020_577(w_020_577, w_007_251, w_001_001);
  nand2 I020_584(w_020_584, w_004_097, w_011_227);
  nand2 I020_586(w_020_586, w_012_009, w_008_090);
  nand2 I020_588(w_020_588, w_006_017, w_007_139);
  not1 I020_590(w_020_590, w_010_506);
  or2  I020_591(w_020_591, w_016_004, w_005_015);
  and2 I020_592(w_020_592, w_012_059, w_005_232);
  not1 I020_595(w_020_595, w_017_055);
  not1 I020_598(w_020_598, w_005_220);
  nand2 I020_599(w_020_599, w_019_014, w_007_018);
  or2  I020_602(w_020_602, w_011_160, w_007_179);
  and2 I020_603(w_020_603, w_012_151, w_017_576);
  or2  I020_604(w_020_604, w_013_013, w_018_010);
  and2 I020_605(w_020_605, w_004_500, w_003_015);
  and2 I020_606(w_020_606, w_011_265, w_010_714);
  not1 I020_607(w_020_607, w_002_270);
  and2 I020_609(w_020_609, w_004_047, w_015_675);
  or2  I020_610(w_020_610, w_007_377, w_007_073);
  not1 I020_615(w_020_615, w_010_564);
  not1 I020_616(w_020_618, w_020_617);
  not1 I020_617(w_020_619, w_020_618);
  and2 I020_618(w_020_620, w_005_019, w_020_619);
  nand2 I020_619(w_020_617, w_020_631, w_020_620);
  or2  I020_620(w_020_625, w_012_158, w_020_624);
  not1 I020_621(w_020_626, w_020_625);
  and2 I020_622(w_020_627, w_019_006, w_020_626);
  or2  I020_623(w_020_628, w_004_319, w_020_627);
  and2 I020_624(w_020_629, w_018_007, w_020_628);
  not1 I020_625(w_020_624, w_020_617);
  and2 I020_626(w_020_631, w_009_270, w_020_629);
  nand2 I021_000(w_021_000, w_014_047, w_004_210);
  or2  I021_001(w_021_001, w_015_377, w_020_250);
  not1 I021_003(w_021_003, w_001_013);
  nand2 I021_004(w_021_004, w_003_066, w_020_494);
  not1 I021_005(w_021_005, w_009_392);
  not1 I021_006(w_021_006, w_011_559);
  and2 I021_007(w_021_007, w_015_323, w_015_258);
  or2  I021_009(w_021_009, w_019_020, w_019_016);
  nand2 I021_010(w_021_010, w_009_023, w_002_227);
  and2 I021_011(w_021_011, w_003_039, w_019_020);
  and2 I021_013(w_021_013, w_016_008, w_003_034);
  not1 I021_014(w_021_014, w_018_039);
  nand2 I021_015(w_021_015, w_008_179, w_003_078);
  and2 I021_016(w_021_016, w_020_115, w_009_125);
  nand2 I021_017(w_021_017, w_018_015, w_012_154);
  not1 I021_018(w_021_018, w_015_170);
  or2  I021_021(w_021_021, w_016_007, w_006_246);
  or2  I021_022(w_021_022, w_014_132, w_012_175);
  and2 I021_023(w_021_023, w_010_009, w_020_147);
  and2 I021_024(w_021_024, w_017_477, w_005_259);
  nand2 I021_025(w_021_025, w_020_132, w_006_213);
  or2  I021_026(w_021_026, w_019_017, w_018_028);
  not1 I021_027(w_021_027, w_006_100);
  and2 I021_028(w_021_028, w_013_559, w_019_000);
  nand2 I021_029(w_021_029, w_008_477, w_000_740);
  not1 I021_032(w_021_032, w_011_257);
  nand2 I021_033(w_021_033, w_008_435, w_004_438);
  or2  I021_034(w_021_034, w_009_245, w_008_426);
  and2 I021_035(w_021_035, w_004_377, w_014_115);
  nand2 I021_036(w_021_036, w_014_103, w_016_004);
  nand2 I021_037(w_021_037, w_005_140, w_003_014);
  and2 I021_039(w_021_039, w_011_112, w_004_493);
  or2  I021_040(w_021_040, w_002_264, w_007_151);
  not1 I021_041(w_021_041, w_011_543);
  nand2 I021_042(w_021_042, w_002_453, w_001_020);
  not1 I021_043(w_021_043, w_017_258);
  or2  I021_044(w_021_044, w_000_588, w_019_000);
  and2 I021_045(w_021_045, w_005_164, w_009_215);
  nand2 I021_047(w_021_047, w_013_115, w_006_012);
  or2  I021_048(w_021_048, w_015_360, w_017_462);
  and2 I021_050(w_021_050, w_013_125, w_009_393);
  not1 I021_051(w_021_051, w_014_083);
  not1 I021_054(w_021_054, w_003_060);
  nand2 I021_055(w_021_055, w_016_003, w_013_380);
  not1 I021_056(w_021_056, w_009_136);
  nand2 I021_059(w_021_059, w_000_214, w_017_492);
  not1 I021_060(w_021_060, w_011_383);
  not1 I021_061(w_021_061, w_019_012);
  and2 I021_062(w_021_062, w_005_305, w_016_002);
  or2  I021_064(w_021_064, w_007_217, w_008_327);
  and2 I021_066(w_021_066, w_014_109, w_001_015);
  and2 I021_067(w_021_067, w_011_469, w_015_041);
  nand2 I021_068(w_021_068, w_015_355, w_004_274);
  or2  I021_069(w_021_069, w_005_042, w_014_022);
  and2 I021_071(w_021_071, w_019_016, w_003_077);
  not1 I021_072(w_021_072, w_009_629);
  nand2 I021_073(w_021_073, w_008_362, w_004_123);
  nand2 I021_074(w_021_074, w_020_517, w_013_397);
  or2  I021_077(w_021_077, w_015_267, w_019_007);
  or2  I021_078(w_021_078, w_002_081, w_020_285);
  not1 I021_079(w_021_079, w_006_135);
  or2  I021_080(w_021_080, w_010_064, w_019_010);
  or2  I021_081(w_021_081, w_010_673, w_016_006);
  and2 I021_082(w_021_082, w_003_000, w_005_154);
  not1 I021_083(w_021_083, w_015_096);
  nand2 I021_084(w_021_084, w_009_363, w_017_119);
  or2  I021_085(w_021_085, w_017_201, w_008_301);
  nand2 I021_086(w_021_086, w_014_241, w_011_566);
  and2 I021_088(w_021_088, w_003_038, w_018_005);
  or2  I021_089(w_021_089, w_002_537, w_012_327);
  not1 I021_090(w_021_090, w_010_056);
  or2  I021_091(w_021_091, w_004_175, w_009_030);
  and2 I021_092(w_021_092, w_018_018, w_018_031);
  not1 I021_093(w_021_093, w_006_031);
  and2 I021_094(w_021_094, w_014_030, w_018_001);
  nand2 I021_095(w_021_095, w_020_451, w_020_183);
  and2 I021_096(w_021_096, w_000_089, w_002_019);
  nand2 I021_097(w_021_097, w_010_006, w_004_407);
  nand2 I021_098(w_021_098, w_014_025, w_007_050);
  and2 I021_099(w_021_099, w_004_058, w_013_132);
  or2  I021_100(w_021_100, w_002_645, w_005_127);
  nand2 I021_101(w_021_101, w_007_219, w_019_005);
  not1 I021_102(w_021_102, w_009_035);
  nand2 I021_103(w_021_103, w_009_137, w_010_646);
  not1 I021_104(w_021_104, w_015_605);
  or2  I021_105(w_021_105, w_006_171, w_002_468);
  and2 I021_106(w_021_106, w_004_236, w_004_416);
  or2  I021_108(w_021_108, w_006_240, w_001_024);
  or2  I021_110(w_021_110, w_013_507, w_002_576);
  and2 I021_111(w_021_111, w_017_194, w_001_001);
  not1 I021_112(w_021_112, w_013_331);
  nand2 I021_113(w_021_113, w_018_029, w_006_159);
  or2  I021_114(w_021_114, w_006_180, w_010_718);
  nand2 I021_115(w_021_115, w_012_202, w_018_032);
  and2 I021_116(w_021_116, w_019_006, w_018_017);
  or2  I021_117(w_021_117, w_020_063, w_012_124);
  not1 I021_118(w_021_118, w_013_073);
  and2 I021_119(w_021_119, w_006_188, w_011_151);
  and2 I021_121(w_021_121, w_003_038, w_003_033);
  not1 I021_122(w_021_122, w_019_016);
  not1 I021_123(w_021_123, w_018_008);
  nand2 I021_124(w_021_124, w_007_192, w_017_126);
  and2 I021_125(w_021_125, w_011_159, w_001_023);
  and2 I021_126(w_021_126, w_007_134, w_014_057);
  not1 I021_127(w_021_127, w_009_609);
  nand2 I021_128(w_021_128, w_010_453, w_013_326);
  not1 I021_130(w_021_130, w_006_192);
  or2  I021_131(w_021_131, w_013_418, w_004_384);
  or2  I021_136(w_021_136, w_013_154, w_002_652);
  and2 I021_137(w_021_137, w_006_144, w_017_088);
  nand2 I021_138(w_021_138, w_019_008, w_017_587);
  and2 I021_139(w_021_139, w_013_563, w_019_020);
  or2  I021_140(w_021_140, w_006_166, w_015_474);
  nand2 I021_141(w_021_141, w_007_463, w_017_631);
  or2  I021_142(w_021_142, w_008_480, w_014_088);
  and2 I021_143(w_021_143, w_020_309, w_011_582);
  or2  I021_144(w_021_144, w_013_107, w_000_059);
  not1 I021_145(w_021_145, w_002_070);
  or2  I021_146(w_021_146, w_019_018, w_020_584);
  nand2 I021_147(w_021_147, w_012_260, w_005_303);
  not1 I021_148(w_021_148, w_020_135);
  nand2 I021_149(w_021_149, w_005_167, w_006_244);
  nand2 I021_150(w_021_150, w_006_106, w_019_008);
  nand2 I021_152(w_021_152, w_017_319, w_003_049);
  not1 I021_153(w_021_153, w_000_718);
  or2  I021_154(w_021_154, w_012_081, w_002_505);
  nand2 I021_155(w_021_155, w_001_007, w_014_057);
  not1 I021_158(w_021_158, w_014_060);
  not1 I021_160(w_021_160, w_002_224);
  or2  I021_161(w_021_161, w_018_028, w_019_014);
  or2  I021_162(w_021_162, w_007_237, w_007_057);
  and2 I021_163(w_021_163, w_012_098, w_009_537);
  or2  I021_164(w_021_164, w_013_048, w_008_526);
  nand2 I021_165(w_021_165, w_010_588, w_003_017);
  not1 I021_166(w_021_166, w_012_350);
  or2  I021_167(w_021_167, w_014_126, w_004_302);
  nand2 I021_168(w_021_168, w_002_632, w_016_006);
  or2  I021_169(w_021_169, w_001_014, w_017_082);
  not1 I021_170(w_021_170, w_003_001);
  nand2 I021_171(w_021_171, w_016_004, w_011_530);
  nand2 I021_172(w_021_172, w_000_319, w_002_202);
  not1 I021_174(w_021_174, w_020_374);
  or2  I021_175(w_021_175, w_002_558, w_006_151);
  nand2 I021_176(w_021_176, w_007_260, w_002_443);
  not1 I021_177(w_021_177, w_006_167);
  not1 I021_179(w_021_179, w_004_214);
  not1 I021_180(w_021_180, w_011_148);
  and2 I021_181(w_021_181, w_002_250, w_002_054);
  not1 I021_182(w_021_182, w_017_036);
  nand2 I021_183(w_021_183, w_019_016, w_001_019);
  nand2 I021_184(w_021_184, w_006_249, w_015_511);
  and2 I021_187(w_021_187, w_009_127, w_014_025);
  or2  I021_188(w_021_188, w_016_007, w_001_032);
  not1 I021_189(w_021_189, w_018_015);
  not1 I021_190(w_021_190, w_014_266);
  not1 I021_191(w_021_191, w_019_004);
  nand2 I021_192(w_021_192, w_001_005, w_020_255);
  or2  I021_193(w_021_193, w_012_028, w_014_148);
  or2  I021_194(w_021_194, w_013_278, w_020_177);
  nand2 I021_195(w_021_195, w_005_250, w_020_473);
  nand2 I021_196(w_021_196, w_016_006, w_009_317);
  nand2 I021_199(w_021_199, w_015_059, w_001_019);
  or2  I021_200(w_021_200, w_016_007, w_016_000);
  nand2 I021_201(w_021_201, w_016_008, w_009_487);
  or2  I021_202(w_021_202, w_008_161, w_001_004);
  or2  I021_203(w_021_203, w_008_654, w_002_429);
  or2  I021_204(w_021_204, w_018_001, w_004_067);
  nand2 I021_205(w_021_205, w_006_066, w_014_177);
  or2  I021_207(w_021_207, w_010_450, w_000_573);
  not1 I021_208(w_021_208, w_008_565);
  nand2 I021_209(w_021_209, w_009_102, w_007_079);
  and2 I021_210(w_021_210, w_007_027, w_013_510);
  not1 I021_211(w_021_211, w_017_578);
  not1 I021_212(w_021_212, w_000_196);
  not1 I021_213(w_021_213, w_006_128);
  and2 I021_214(w_021_214, w_005_136, w_019_002);
  not1 I021_215(w_021_215, w_006_011);
  nand2 I021_216(w_021_216, w_013_204, w_009_130);
  or2  I021_217(w_021_217, w_010_656, w_018_029);
  nand2 I021_218(w_021_218, w_001_006, w_014_184);
  or2  I021_219(w_021_219, w_011_202, w_016_002);
  or2  I021_220(w_021_220, w_020_386, w_017_338);
  nand2 I021_221(w_021_221, w_015_317, w_006_188);
  or2  I021_222(w_021_222, w_014_003, w_011_042);
  and2 I021_223(w_021_223, w_014_012, w_012_249);
  not1 I021_224(w_021_224, w_001_029);
  not1 I021_225(w_021_225, w_013_098);
  nand2 I021_226(w_021_226, w_001_024, w_001_022);
  not1 I021_227(w_021_227, w_001_035);
  or2  I021_230(w_021_230, w_003_049, w_013_068);
  and2 I021_231(w_021_231, w_001_021, w_015_214);
  and2 I021_232(w_021_232, w_005_026, w_008_052);
  or2  I021_233(w_021_233, w_009_092, w_017_246);
  nand2 I021_234(w_021_234, w_005_260, w_016_001);
  not1 I021_235(w_021_235, w_007_299);
  or2  I021_236(w_021_236, w_009_224, w_008_495);
  and2 I021_237(w_021_237, w_019_006, w_015_044);
  not1 I021_238(w_021_238, w_009_488);
  not1 I021_239(w_021_239, w_014_111);
  not1 I021_240(w_021_240, w_018_009);
  not1 I021_241(w_021_241, w_019_013);
  and2 I021_242(w_021_242, w_010_453, w_019_003);
  not1 I021_243(w_021_243, w_018_044);
  nand2 I021_244(w_021_244, w_006_252, w_020_090);
  nand2 I021_246(w_021_246, w_017_003, w_015_183);
  or2  I021_247(w_021_247, w_002_474, w_010_611);
  and2 I021_248(w_021_248, w_007_035, w_006_240);
  not1 I021_249(w_021_249, w_002_383);
  and2 I021_250(w_021_250, w_020_164, w_016_006);
  and2 I021_251(w_021_251, w_015_044, w_014_001);
  nand2 I021_255(w_021_255, w_017_006, w_010_642);
  or2  I021_256(w_021_256, w_001_002, w_015_432);
  not1 I021_257(w_021_257, w_020_539);
  nand2 I021_259(w_021_259, w_012_250, w_005_047);
  nand2 I021_261(w_021_261, w_017_291, w_010_338);
  nand2 I021_262(w_021_262, w_006_091, w_018_035);
  or2  I021_263(w_021_263, w_020_028, w_020_562);
  not1 I021_264(w_021_264, w_017_653);
  or2  I021_265(w_021_265, w_006_242, w_003_074);
  or2  I021_266(w_021_266, w_006_210, w_019_013);
  not1 I021_267(w_021_267, w_010_245);
  not1 I021_270(w_021_270, w_008_522);
  or2  I021_271(w_021_271, w_020_396, w_009_084);
  or2  I021_272(w_021_272, w_014_211, w_015_372);
  or2  I021_273(w_021_273, w_020_288, w_006_228);
  not1 I021_274(w_021_274, w_014_025);
  and2 I021_275(w_020_622, w_009_154, w_020_617);
  nand2 I022_000(w_022_000, w_001_029, w_017_333);
  not1 I022_001(w_022_001, w_008_149);
  nand2 I022_003(w_022_003, w_003_015, w_005_025);
  not1 I022_005(w_022_005, w_015_501);
  not1 I022_006(w_022_006, w_007_102);
  nand2 I022_009(w_022_009, w_000_477, w_006_169);
  or2  I022_010(w_022_010, w_009_162, w_000_741);
  or2  I022_011(w_022_011, w_002_599, w_017_364);
  or2  I022_012(w_022_012, w_008_417, w_015_054);
  nand2 I022_013(w_022_013, w_016_004, w_020_031);
  not1 I022_017(w_022_017, w_005_125);
  or2  I022_020(w_022_020, w_013_175, w_014_044);
  not1 I022_021(w_022_021, w_007_178);
  and2 I022_023(w_022_023, w_017_130, w_003_021);
  or2  I022_024(w_022_024, w_003_075, w_002_046);
  and2 I022_026(w_022_026, w_020_271, w_010_587);
  nand2 I022_029(w_022_029, w_004_088, w_013_507);
  not1 I022_030(w_022_030, w_015_408);
  nand2 I022_031(w_022_031, w_018_041, w_010_660);
  or2  I022_032(w_022_032, w_008_179, w_021_210);
  nand2 I022_033(w_022_033, w_019_015, w_021_037);
  nand2 I022_034(w_022_034, w_021_220, w_018_043);
  not1 I022_035(w_022_035, w_018_008);
  not1 I022_036(w_022_036, w_000_448);
  or2  I022_037(w_022_037, w_019_008, w_006_244);
  or2  I022_038(w_022_038, w_001_000, w_009_469);
  nand2 I022_039(w_022_039, w_018_018, w_000_151);
  and2 I022_041(w_022_041, w_005_054, w_008_027);
  nand2 I022_042(w_022_042, w_004_387, w_011_063);
  nand2 I022_043(w_022_043, w_001_034, w_009_377);
  not1 I022_044(w_022_044, w_011_634);
  and2 I022_045(w_022_045, w_018_034, w_011_172);
  not1 I022_048(w_022_048, w_002_428);
  nand2 I022_050(w_022_050, w_006_150, w_008_428);
  or2  I022_051(w_022_051, w_012_081, w_002_706);
  nand2 I022_052(w_022_052, w_020_562, w_009_031);
  nand2 I022_053(w_022_053, w_020_091, w_007_397);
  nand2 I022_054(w_022_054, w_019_007, w_012_271);
  or2  I022_055(w_022_055, w_012_252, w_011_281);
  nand2 I022_056(w_022_056, w_017_657, w_006_241);
  or2  I022_058(w_022_058, w_021_022, w_012_092);
  not1 I022_059(w_022_059, w_021_025);
  nand2 I022_061(w_022_061, w_010_450, w_005_111);
  and2 I022_062(w_022_062, w_016_005, w_007_181);
  or2  I022_064(w_022_064, w_013_297, w_004_424);
  or2  I022_065(w_022_065, w_016_004, w_008_274);
  nand2 I022_066(w_022_066, w_015_180, w_017_462);
  not1 I022_068(w_022_068, w_004_286);
  and2 I022_071(w_022_071, w_021_150, w_000_688);
  or2  I022_074(w_022_074, w_007_294, w_000_620);
  and2 I022_076(w_022_076, w_011_193, w_007_131);
  and2 I022_077(w_022_077, w_015_029, w_020_267);
  or2  I022_079(w_022_079, w_001_016, w_015_073);
  and2 I022_080(w_022_080, w_005_144, w_020_461);
  not1 I022_081(w_022_081, w_020_084);
  and2 I022_082(w_022_082, w_000_743, w_010_355);
  nand2 I022_083(w_022_083, w_017_487, w_016_001);
  not1 I022_084(w_022_084, w_012_116);
  and2 I022_086(w_022_086, w_016_001, w_014_258);
  nand2 I022_087(w_022_087, w_017_240, w_015_134);
  nand2 I022_088(w_022_088, w_011_387, w_005_212);
  or2  I022_089(w_022_089, w_016_007, w_002_473);
  not1 I022_090(w_022_090, w_018_007);
  or2  I022_093(w_022_093, w_006_139, w_019_019);
  and2 I022_094(w_022_094, w_010_377, w_019_010);
  nand2 I022_097(w_022_097, w_007_103, w_015_139);
  nand2 I022_098(w_022_098, w_009_318, w_013_573);
  not1 I022_100(w_022_100, w_001_030);
  not1 I022_102(w_022_102, w_015_084);
  not1 I022_103(w_022_103, w_017_151);
  or2  I022_104(w_022_104, w_014_214, w_000_565);
  nand2 I022_111(w_022_111, w_000_288, w_002_709);
  or2  I022_112(w_022_112, w_013_066, w_008_018);
  nand2 I022_114(w_022_114, w_000_427, w_013_322);
  nand2 I022_115(w_022_115, w_013_118, w_018_015);
  or2  I022_117(w_022_117, w_004_273, w_011_554);
  and2 I022_118(w_022_118, w_009_183, w_000_591);
  and2 I022_119(w_022_119, w_005_061, w_021_174);
  nand2 I022_120(w_022_120, w_002_148, w_018_006);
  and2 I022_123(w_022_123, w_012_225, w_015_222);
  nand2 I022_124(w_022_124, w_005_009, w_005_315);
  and2 I022_125(w_022_125, w_003_000, w_012_054);
  or2  I022_126(w_022_126, w_011_130, w_013_413);
  or2  I022_128(w_022_128, w_019_005, w_019_007);
  and2 I022_129(w_022_129, w_020_158, w_014_284);
  and2 I022_130(w_022_130, w_007_176, w_000_418);
  not1 I022_131(w_022_131, w_014_042);
  nand2 I022_132(w_022_132, w_004_082, w_015_015);
  and2 I022_134(w_022_134, w_006_033, w_019_020);
  and2 I022_135(w_022_135, w_015_671, w_001_016);
  or2  I022_136(w_022_136, w_013_426, w_017_597);
  nand2 I022_137(w_022_137, w_017_215, w_001_029);
  nand2 I022_138(w_022_138, w_009_342, w_014_009);
  nand2 I022_140(w_022_140, w_003_026, w_017_089);
  and2 I022_141(w_022_141, w_015_396, w_013_158);
  nand2 I022_142(w_022_142, w_012_003, w_000_023);
  and2 I022_144(w_022_144, w_020_136, w_021_263);
  nand2 I022_145(w_022_145, w_013_121, w_015_210);
  not1 I022_148(w_022_148, w_005_092);
  or2  I022_149(w_022_149, w_005_305, w_013_036);
  not1 I022_150(w_022_150, w_007_059);
  not1 I022_151(w_022_151, w_003_023);
  or2  I022_152(w_022_152, w_008_210, w_005_170);
  nand2 I022_153(w_022_153, w_007_078, w_009_603);
  or2  I022_154(w_022_154, w_005_231, w_020_571);
  and2 I022_155(w_022_155, w_018_033, w_021_059);
  not1 I022_158(w_022_158, w_011_108);
  and2 I022_160(w_022_160, w_003_080, w_015_370);
  and2 I022_161(w_022_161, w_011_494, w_000_437);
  not1 I022_163(w_022_163, w_012_022);
  and2 I022_164(w_022_164, w_004_116, w_013_339);
  not1 I022_165(w_022_165, w_002_087);
  or2  I022_167(w_022_167, w_016_000, w_010_773);
  and2 I022_168(w_022_168, w_019_019, w_002_116);
  or2  I022_170(w_022_170, w_018_024, w_015_396);
  nand2 I022_172(w_022_172, w_002_120, w_010_453);
  and2 I022_173(w_022_173, w_005_056, w_014_162);
  or2  I022_174(w_022_174, w_019_012, w_006_033);
  not1 I022_175(w_022_175, w_011_057);
  and2 I022_177(w_022_177, w_020_446, w_001_015);
  and2 I022_181(w_022_181, w_005_097, w_007_212);
  or2  I022_183(w_022_183, w_007_330, w_020_131);
  or2  I022_185(w_022_185, w_015_641, w_012_086);
  nand2 I022_186(w_022_186, w_020_513, w_010_779);
  and2 I022_187(w_022_187, w_002_292, w_011_637);
  not1 I022_188(w_022_188, w_002_211);
  or2  I022_193(w_022_193, w_020_622, w_001_001);
  not1 I022_194(w_022_194, w_016_003);
  and2 I022_195(w_022_195, w_016_004, w_021_082);
  not1 I022_196(w_022_196, w_021_018);
  and2 I022_198(w_022_198, w_008_298, w_008_033);
  not1 I022_199(w_022_199, w_015_374);
  not1 I022_200(w_022_200, w_020_123);
  nand2 I022_201(w_022_201, w_002_034, w_014_178);
  and2 I022_202(w_022_202, w_006_236, w_018_033);
  and2 I022_204(w_022_204, w_005_159, w_018_014);
  nand2 I022_205(w_022_205, w_004_402, w_000_644);
  or2  I022_206(w_022_206, w_013_570, w_007_225);
  or2  I022_207(w_022_207, w_020_107, w_001_026);
  or2  I022_210(w_022_210, w_004_425, w_018_001);
  or2  I022_211(w_022_211, w_009_071, w_014_165);
  not1 I022_213(w_022_213, w_010_009);
  not1 I022_214(w_022_214, w_009_109);
  and2 I022_219(w_022_219, w_021_100, w_011_269);
  or2  I022_220(w_022_220, w_019_007, w_017_620);
  not1 I022_221(w_022_221, w_015_232);
  and2 I022_226(w_022_226, w_012_306, w_003_031);
  nand2 I022_227(w_022_227, w_000_744, w_007_353);
  not1 I022_229(w_022_229, w_021_055);
  or2  I022_231(w_022_231, w_007_098, w_005_135);
  not1 I022_232(w_022_232, w_001_021);
  nand2 I022_234(w_022_234, w_014_194, w_009_500);
  or2  I022_235(w_022_235, w_001_000, w_005_087);
  nand2 I022_236(w_022_236, w_005_302, w_010_094);
  not1 I022_237(w_022_237, w_021_210);
  and2 I022_238(w_022_238, w_004_169, w_011_035);
  and2 I022_239(w_022_239, w_009_047, w_011_128);
  nand2 I022_240(w_022_240, w_000_599, w_015_230);
  or2  I022_241(w_022_241, w_002_018, w_019_011);
  and2 I022_243(w_022_243, w_009_359, w_010_724);
  nand2 I022_245(w_022_245, w_020_000, w_014_176);
  or2  I022_247(w_022_247, w_017_475, w_021_140);
  not1 I022_248(w_022_248, w_006_215);
  or2  I022_249(w_022_249, w_003_030, w_017_028);
  or2  I022_251(w_022_251, w_021_168, w_002_253);
  nand2 I022_252(w_022_252, w_016_006, w_007_211);
  or2  I022_253(w_022_253, w_019_007, w_010_408);
  and2 I022_255(w_022_255, w_010_653, w_011_169);
  or2  I022_256(w_022_256, w_019_019, w_000_745);
  not1 I022_258(w_022_258, w_007_407);
  and2 I022_259(w_022_259, w_012_170, w_016_001);
  or2  I022_261(w_022_261, w_021_041, w_011_441);
  and2 I022_262(w_022_262, w_000_163, w_020_192);
  nand2 I022_263(w_022_263, w_018_004, w_001_031);
  nand2 I022_264(w_022_264, w_021_168, w_005_108);
  or2  I022_265(w_022_265, w_010_130, w_003_071);
  and2 I022_266(w_022_266, w_004_174, w_017_329);
  nand2 I022_267(w_022_267, w_015_222, w_014_247);
  and2 I022_268(w_022_268, w_006_135, w_009_100);
  nand2 I022_269(w_022_269, w_006_013, w_020_427);
  nand2 I022_270(w_022_270, w_003_039, w_019_017);
  and2 I022_271(w_022_271, w_016_003, w_021_042);
  or2  I022_272(w_022_272, w_021_050, w_021_161);
  nand2 I022_276(w_022_276, w_007_175, w_017_295);
  and2 I022_277(w_022_277, w_002_025, w_017_611);
  not1 I022_279(w_022_279, w_001_024);
  not1 I022_280(w_022_280, w_019_010);
  not1 I022_281(w_022_281, w_013_160);
  or2  I022_282(w_022_282, w_014_220, w_015_029);
  nand2 I022_283(w_022_283, w_001_004, w_011_560);
  nand2 I022_287(w_022_287, w_005_310, w_008_524);
  nand2 I022_288(w_022_288, w_019_012, w_010_245);
  or2  I022_290(w_022_290, w_002_423, w_002_711);
  nand2 I022_291(w_022_291, w_016_003, w_011_180);
  nand2 I022_293(w_022_293, w_019_017, w_006_234);
  nand2 I022_294(w_022_294, w_012_316, w_011_198);
  and2 I022_295(w_022_295, w_009_435, w_002_574);
  or2  I022_296(w_022_296, w_002_401, w_006_000);
  or2  I022_297(w_022_297, w_009_417, w_006_150);
  or2  I022_298(w_022_298, w_018_043, w_002_518);
  or2  I022_300(w_022_300, w_003_011, w_009_504);
  and2 I022_303(w_022_303, w_000_632, w_020_071);
  nand2 I022_304(w_022_304, w_015_647, w_003_019);
  or2  I022_305(w_022_305, w_009_543, w_017_111);
  nand2 I022_307(w_022_307, w_003_064, w_020_525);
  and2 I022_309(w_022_309, w_012_090, w_016_002);
  nand2 I022_310(w_022_310, w_016_000, w_016_005);
  or2  I022_311(w_022_311, w_004_446, w_006_057);
  and2 I022_313(w_022_313, w_020_506, w_001_021);
  and2 I022_315(w_022_315, w_000_747, w_018_006);
  nand2 I022_316(w_022_316, w_011_440, w_000_265);
  and2 I022_319(w_022_319, w_018_004, w_017_146);
  not1 I022_320(w_022_320, w_016_006);
  and2 I022_321(w_022_321, w_014_058, w_005_025);
  not1 I022_322(w_022_322, w_005_011);
  not1 I022_323(w_022_323, w_016_000);
  and2 I022_328(w_022_328, w_010_685, w_000_748);
  nand2 I022_330(w_022_330, w_010_342, w_001_027);
  not1 I022_331(w_022_331, w_009_167);
  not1 I022_332(w_022_332, w_014_102);
  nand2 I022_333(w_022_333, w_003_062, w_000_548);
  not1 I022_334(w_022_334, w_009_390);
  and2 I022_336(w_022_336, w_011_383, w_005_233);
  or2  I022_337(w_022_337, w_006_201, w_011_291);
  or2  I022_341(w_022_341, w_001_034, w_004_370);
  or2  I022_342(w_022_342, w_018_029, w_011_124);
  and2 I022_343(w_022_343, w_016_000, w_011_329);
  nand2 I022_344(w_022_344, w_000_172, w_008_745);
  nand2 I022_345(w_022_345, w_017_651, w_003_050);
  and2 I022_347(w_022_347, w_007_328, w_007_441);
  not1 I022_348(w_022_348, w_010_005);
  nand2 I022_349(w_022_349, w_021_203, w_021_144);
  nand2 I022_351(w_022_351, w_006_227, w_006_245);
  not1 I022_352(w_022_352, w_007_236);
  or2  I022_353(w_022_353, w_000_573, w_009_109);
  nand2 I022_355(w_022_355, w_014_269, w_016_006);
  nand2 I022_356(w_022_356, w_015_008, w_009_389);
  nand2 I022_357(w_022_357, w_009_041, w_018_001);
  and2 I022_360(w_022_360, w_010_250, w_021_017);
  nand2 I022_361(w_022_361, w_002_072, w_014_289);
  not1 I022_362(w_022_362, w_006_194);
  nand2 I022_364(w_022_364, w_020_043, w_010_097);
  not1 I022_365(w_022_365, w_002_099);
  nand2 I022_366(w_022_366, w_018_039, w_009_537);
  nand2 I022_367(w_022_367, w_018_014, w_013_034);
  not1 I022_368(w_022_368, w_015_043);
  and2 I022_369(w_022_369, w_002_047, w_013_452);
  nand2 I022_370(w_022_370, w_017_043, w_010_736);
  nand2 I022_373(w_022_373, w_012_316, w_016_001);
  nand2 I022_376(w_022_376, w_015_566, w_006_212);
  not1 I022_378(w_022_378, w_015_506);
  and2 I022_380(w_022_380, w_018_022, w_019_013);
  not1 I022_381(w_022_381, w_002_563);
  or2  I022_382(w_022_382, w_001_020, w_009_124);
  and2 I022_383(w_022_383, w_004_144, w_021_131);
  and2 I022_384(w_022_384, w_001_004, w_015_386);
  nand2 I022_385(w_022_385, w_009_092, w_009_607);
  or2  I022_386(w_022_386, w_015_448, w_019_017);
  nand2 I022_388(w_022_388, w_002_470, w_011_306);
  or2  I022_389(w_022_389, w_017_670, w_013_210);
  or2  I022_390(w_022_390, w_011_198, w_013_214);
  not1 I022_392(w_022_392, w_003_079);
  not1 I022_393(w_022_393, w_000_619);
  not1 I022_395(w_022_395, w_003_052);
  and2 I022_397(w_022_397, w_012_018, w_019_010);
  and2 I022_399(w_022_399, w_000_396, w_019_008);
  not1 I022_401(w_022_401, w_009_231);
  not1 I022_404(w_022_404, w_004_265);
  nand2 I022_407(w_022_407, w_002_319, w_014_031);
  nand2 I022_408(w_022_408, w_012_168, w_002_183);
  nand2 I023_000(w_023_000, w_021_032, w_010_347);
  nand2 I023_002(w_023_002, w_002_401, w_006_081);
  and2 I023_003(w_023_003, w_003_060, w_016_000);
  and2 I023_005(w_023_005, w_010_099, w_012_239);
  or2  I023_006(w_023_006, w_010_259, w_008_486);
  not1 I023_007(w_023_007, w_002_306);
  or2  I023_008(w_023_008, w_021_010, w_007_038);
  or2  I023_009(w_023_009, w_007_119, w_017_483);
  or2  I023_011(w_023_011, w_009_462, w_012_058);
  or2  I023_012(w_023_012, w_001_014, w_022_328);
  not1 I023_013(w_023_013, w_001_036);
  nand2 I023_015(w_023_015, w_004_002, w_017_141);
  and2 I023_016(w_023_016, w_005_305, w_013_159);
  and2 I023_017(w_023_017, w_012_350, w_013_194);
  and2 I023_018(w_023_018, w_002_155, w_017_422);
  not1 I023_019(w_023_019, w_010_713);
  or2  I023_020(w_023_020, w_006_183, w_010_471);
  and2 I023_021(w_023_021, w_007_111, w_002_570);
  not1 I023_023(w_023_023, w_019_003);
  not1 I023_024(w_023_024, w_000_548);
  not1 I023_025(w_023_025, w_008_621);
  and2 I023_026(w_023_026, w_017_496, w_001_025);
  not1 I023_027(w_023_027, w_016_001);
  nand2 I023_028(w_023_028, w_015_633, w_015_023);
  or2  I023_029(w_023_029, w_022_037, w_013_565);
  or2  I023_031(w_023_031, w_019_015, w_000_610);
  not1 I023_032(w_023_032, w_008_432);
  nand2 I023_033(w_023_033, w_003_055, w_002_303);
  not1 I023_034(w_023_034, w_012_179);
  not1 I023_035(w_023_035, w_021_090);
  and2 I023_037(w_023_037, w_020_281, w_015_114);
  and2 I023_038(w_023_038, w_019_003, w_004_190);
  or2  I023_039(w_023_039, w_022_094, w_015_561);
  or2  I023_040(w_023_040, w_012_241, w_007_198);
  nand2 I023_041(w_023_041, w_013_411, w_007_154);
  and2 I023_042(w_023_042, w_009_090, w_016_006);
  not1 I023_043(w_023_043, w_005_098);
  nand2 I023_044(w_023_044, w_014_267, w_005_144);
  and2 I023_045(w_023_045, w_009_085, w_016_008);
  not1 I023_046(w_023_046, w_002_435);
  nand2 I023_047(w_023_047, w_008_228, w_006_172);
  and2 I023_048(w_023_048, w_014_287, w_001_035);
  and2 I023_049(w_023_049, w_005_140, w_017_055);
  or2  I023_051(w_023_051, w_007_140, w_013_001);
  not1 I023_052(w_023_052, w_000_501);
  nand2 I023_053(w_023_053, w_019_000, w_004_086);
  not1 I023_054(w_023_054, w_012_024);
  not1 I023_055(w_023_055, w_007_162);
  not1 I023_056(w_023_056, w_001_035);
  not1 I023_058(w_023_058, w_018_011);
  or2  I023_059(w_023_059, w_011_428, w_021_144);
  not1 I023_060(w_023_060, w_012_206);
  or2  I023_062(w_023_062, w_017_297, w_000_406);
  not1 I023_063(w_023_063, w_004_020);
  not1 I023_064(w_023_064, w_005_023);
  and2 I023_065(w_023_065, w_020_003, w_002_308);
  not1 I023_066(w_023_066, w_018_025);
  and2 I023_067(w_023_067, w_012_080, w_000_330);
  not1 I023_068(w_023_068, w_007_293);
  nand2 I023_069(w_023_069, w_017_419, w_001_016);
  not1 I023_070(w_023_070, w_012_347);
  and2 I023_071(w_023_071, w_001_033, w_019_020);
  and2 I023_073(w_023_073, w_014_043, w_001_036);
  nand2 I023_074(w_023_074, w_013_106, w_002_070);
  and2 I023_075(w_023_075, w_004_397, w_003_009);
  and2 I023_076(w_023_076, w_021_165, w_003_023);
  and2 I023_077(w_023_077, w_014_252, w_017_589);
  nand2 I023_078(w_023_078, w_018_022, w_000_238);
  nand2 I023_079(w_023_079, w_012_029, w_014_225);
  not1 I023_080(w_023_080, w_010_261);
  and2 I023_081(w_023_081, w_007_331, w_021_009);
  and2 I023_082(w_023_082, w_001_004, w_000_641);
  or2  I023_083(w_023_083, w_003_035, w_020_149);
  or2  I023_084(w_023_084, w_009_554, w_018_010);
  and2 I023_086(w_023_086, w_011_059, w_006_075);
  and2 I023_087(w_023_087, w_000_053, w_007_094);
  and2 I023_088(w_023_088, w_009_507, w_008_015);
  and2 I023_090(w_023_090, w_012_345, w_013_118);
  and2 I023_091(w_023_091, w_015_067, w_010_581);
  not1 I023_092(w_023_092, w_005_233);
  or2  I023_093(w_023_093, w_011_014, w_005_168);
  not1 I023_095(w_023_095, w_001_006);
  not1 I023_096(w_023_096, w_014_016);
  not1 I023_098(w_023_098, w_013_022);
  not1 I023_099(w_023_099, w_010_539);
  and2 I023_100(w_023_100, w_003_082, w_002_261);
  not1 I023_101(w_023_101, w_019_000);
  not1 I023_102(w_023_102, w_007_218);
  or2  I023_103(w_023_103, w_017_035, w_015_624);
  or2  I023_104(w_023_104, w_006_006, w_000_710);
  nand2 I023_105(w_023_105, w_018_020, w_009_022);
  or2  I023_106(w_023_106, w_008_747, w_010_014);
  nand2 I023_107(w_023_107, w_007_032, w_006_084);
  and2 I023_108(w_023_108, w_019_015, w_007_149);
  nand2 I023_109(w_023_109, w_001_026, w_007_340);
  not1 I023_110(w_023_110, w_009_478);
  and2 I023_111(w_023_111, w_009_388, w_013_032);
  and2 I023_112(w_023_112, w_000_684, w_004_197);
  nand2 I023_113(w_023_113, w_008_192, w_020_569);
  not1 I023_114(w_023_114, w_020_205);
  nand2 I023_115(w_023_115, w_016_004, w_009_046);
  nand2 I023_116(w_023_116, w_004_072, w_022_320);
  nand2 I023_117(w_023_117, w_002_408, w_021_125);
  or2  I023_120(w_023_120, w_020_425, w_012_094);
  nand2 I023_121(w_023_121, w_014_196, w_019_009);
  or2  I023_122(w_023_122, w_006_210, w_006_047);
  or2  I023_123(w_023_123, w_014_125, w_018_003);
  not1 I023_124(w_023_124, w_014_081);
  not1 I023_125(w_023_125, w_020_095);
  or2  I023_128(w_023_128, w_019_020, w_006_147);
  nand2 I023_129(w_023_129, w_011_551, w_010_009);
  not1 I023_130(w_023_130, w_003_023);
  or2  I023_131(w_023_131, w_012_312, w_017_306);
  nand2 I023_132(w_023_132, w_019_014, w_002_243);
  and2 I023_134(w_023_134, w_016_002, w_006_030);
  nand2 I023_135(w_023_135, w_012_178, w_020_072);
  and2 I023_136(w_023_136, w_001_027, w_018_003);
  and2 I023_137(w_023_137, w_011_368, w_022_265);
  not1 I023_138(w_023_138, w_005_113);
  not1 I023_139(w_023_139, w_008_708);
  or2  I023_141(w_023_141, w_013_095, w_001_011);
  and2 I023_142(w_023_142, w_008_318, w_001_019);
  and2 I023_143(w_023_143, w_019_007, w_017_121);
  or2  I023_144(w_023_144, w_022_336, w_003_054);
  not1 I023_145(w_023_145, w_002_620);
  or2  I023_146(w_023_146, w_015_158, w_021_067);
  or2  I023_147(w_023_147, w_010_272, w_011_572);
  nand2 I023_148(w_023_148, w_012_232, w_000_485);
  not1 I023_149(w_023_149, w_018_034);
  not1 I023_150(w_023_150, w_014_071);
  and2 I023_151(w_023_151, w_012_298, w_007_013);
  nand2 I023_152(w_023_152, w_011_033, w_010_240);
  nand2 I023_153(w_023_153, w_019_000, w_007_143);
  and2 I023_154(w_023_154, w_017_097, w_016_000);
  nand2 I023_155(w_023_155, w_022_183, w_010_691);
  nand2 I023_156(w_023_156, w_005_183, w_016_003);
  and2 I023_157(w_023_157, w_019_009, w_000_568);
  and2 I023_158(w_023_158, w_008_541, w_003_013);
  or2  I023_159(w_023_159, w_018_039, w_021_039);
  nand2 I023_160(w_023_160, w_003_034, w_018_030);
  not1 I023_161(w_023_161, w_011_589);
  nand2 I023_162(w_023_162, w_022_032, w_001_006);
  not1 I023_164(w_023_164, w_001_020);
  not1 I023_165(w_023_165, w_003_024);
  and2 I023_166(w_023_166, w_015_613, w_014_049);
  and2 I023_169(w_023_169, w_012_119, w_022_003);
  or2  I023_170(w_023_170, w_017_006, w_015_236);
  and2 I023_171(w_023_171, w_010_327, w_008_729);
  not1 I023_172(w_023_172, w_011_003);
  nand2 I023_173(w_023_173, w_002_247, w_014_288);
  and2 I023_175(w_023_175, w_013_269, w_006_121);
  nand2 I023_176(w_023_176, w_005_273, w_011_317);
  not1 I023_178(w_023_178, w_007_432);
  or2  I023_179(w_023_179, w_021_041, w_018_025);
  nand2 I023_181(w_023_181, w_005_077, w_002_249);
  not1 I023_183(w_023_183, w_009_123);
  not1 I023_184(w_023_184, w_000_004);
  or2  I023_186(w_023_186, w_002_066, w_017_315);
  nand2 I023_188(w_023_188, w_004_401, w_000_308);
  nand2 I023_189(w_023_189, w_014_081, w_012_227);
  not1 I023_191(w_023_191, w_000_739);
  or2  I023_192(w_023_192, w_005_293, w_003_083);
  nand2 I023_193(w_023_193, w_020_109, w_000_630);
  nand2 I023_194(w_023_194, w_002_690, w_013_432);
  nand2 I023_195(w_023_195, w_007_258, w_021_061);
  nand2 I023_196(w_023_196, w_011_639, w_018_008);
  nand2 I023_197(w_023_197, w_019_000, w_017_428);
  and2 I023_198(w_023_198, w_001_012, w_014_116);
  or2  I023_199(w_023_199, w_004_190, w_019_001);
  and2 I023_200(w_023_200, w_014_084, w_018_034);
  not1 I023_201(w_023_201, w_012_209);
  not1 I023_202(w_023_202, w_011_622);
  or2  I023_203(w_023_203, w_016_004, w_004_163);
  or2  I023_205(w_023_205, w_018_015, w_012_331);
  not1 I023_206(w_023_206, w_016_002);
  and2 I023_207(w_023_207, w_015_445, w_000_588);
  and2 I023_208(w_023_208, w_021_231, w_008_050);
  or2  I023_210(w_023_210, w_005_261, w_011_136);
  and2 I023_212(w_023_212, w_001_025, w_021_110);
  not1 I023_213(w_023_213, w_014_285);
  nand2 I023_214(w_023_214, w_006_030, w_019_018);
  nand2 I023_215(w_023_215, w_017_165, w_021_149);
  not1 I023_216(w_023_216, w_005_054);
  or2  I023_217(w_023_217, w_005_163, w_009_259);
  and2 I024_000(w_024_000, w_018_025, w_008_118);
  nand2 I024_003(w_024_003, w_017_037, w_005_254);
  not1 I024_004(w_024_004, w_002_337);
  or2  I024_005(w_024_005, w_008_418, w_019_009);
  not1 I024_007(w_024_007, w_017_657);
  not1 I024_008(w_024_008, w_023_175);
  nand2 I024_009(w_024_009, w_015_111, w_002_070);
  not1 I024_010(w_024_010, w_020_148);
  nand2 I024_013(w_024_013, w_023_056, w_010_185);
  not1 I024_015(w_024_015, w_017_408);
  or2  I024_016(w_024_016, w_000_397, w_023_092);
  and2 I024_017(w_024_017, w_011_011, w_023_090);
  and2 I024_018(w_024_018, w_014_101, w_020_335);
  or2  I024_020(w_024_020, w_008_360, w_007_314);
  and2 I024_022(w_024_022, w_020_501, w_006_247);
  not1 I024_024(w_024_024, w_009_373);
  or2  I024_025(w_024_025, w_011_174, w_003_066);
  not1 I024_026(w_024_026, w_003_056);
  and2 I024_027(w_024_027, w_009_621, w_004_227);
  and2 I024_028(w_024_028, w_006_010, w_009_320);
  or2  I024_029(w_024_029, w_022_393, w_017_315);
  nand2 I024_030(w_024_030, w_005_127, w_004_311);
  nand2 I024_032(w_024_032, w_013_539, w_005_224);
  not1 I024_034(w_024_034, w_006_234);
  and2 I024_035(w_024_035, w_007_131, w_001_009);
  not1 I024_036(w_024_036, w_010_264);
  nand2 I024_039(w_024_039, w_000_254, w_008_587);
  and2 I024_040(w_024_040, w_016_006, w_013_561);
  or2  I024_041(w_024_041, w_011_203, w_015_104);
  nand2 I024_042(w_024_042, w_022_307, w_008_404);
  not1 I024_044(w_024_044, w_009_144);
  and2 I024_045(w_024_045, w_008_339, w_016_001);
  nand2 I024_048(w_024_048, w_018_007, w_007_094);
  nand2 I024_049(w_024_049, w_015_301, w_002_676);
  and2 I024_051(w_024_051, w_010_311, w_002_013);
  or2  I024_054(w_024_054, w_003_005, w_009_109);
  or2  I024_055(w_024_055, w_008_555, w_001_010);
  or2  I024_056(w_024_056, w_019_002, w_023_041);
  not1 I024_057(w_024_057, w_007_017);
  not1 I024_059(w_024_059, w_010_177);
  nand2 I024_060(w_024_060, w_012_336, w_021_115);
  not1 I024_061(w_024_061, w_000_210);
  nand2 I024_062(w_024_062, w_014_215, w_015_161);
  or2  I024_064(w_024_064, w_013_123, w_001_036);
  and2 I024_065(w_024_065, w_010_249, w_021_080);
  and2 I024_068(w_024_068, w_020_314, w_016_000);
  not1 I024_070(w_024_070, w_000_749);
  or2  I024_071(w_024_071, w_001_014, w_001_024);
  and2 I024_073(w_024_073, w_005_212, w_000_577);
  and2 I024_077(w_024_077, w_015_123, w_011_392);
  not1 I024_079(w_024_079, w_017_107);
  and2 I024_081(w_024_081, w_018_024, w_000_179);
  not1 I024_082(w_024_082, w_020_020);
  or2  I024_083(w_024_083, w_023_059, w_014_273);
  and2 I024_086(w_024_086, w_005_158, w_013_318);
  or2  I024_088(w_024_088, w_000_613, w_011_532);
  or2  I024_089(w_024_089, w_016_001, w_020_591);
  or2  I024_090(w_024_090, w_000_588, w_010_478);
  and2 I024_092(w_024_092, w_018_034, w_004_050);
  or2  I024_093(w_024_093, w_009_078, w_008_737);
  and2 I024_095(w_024_095, w_004_278, w_017_053);
  and2 I024_096(w_024_096, w_014_196, w_021_211);
  and2 I024_097(w_024_097, w_023_164, w_011_114);
  and2 I024_098(w_024_098, w_003_035, w_021_060);
  nand2 I024_099(w_024_099, w_015_376, w_022_237);
  nand2 I024_101(w_024_101, w_004_095, w_012_088);
  and2 I024_102(w_024_102, w_020_604, w_008_137);
  not1 I024_103(w_024_103, w_000_264);
  not1 I024_105(w_024_105, w_006_148);
  not1 I024_107(w_024_107, w_018_036);
  nand2 I024_108(w_024_108, w_002_588, w_006_247);
  and2 I024_109(w_024_109, w_005_230, w_006_041);
  or2  I024_110(w_024_110, w_010_289, w_018_008);
  not1 I024_115(w_024_115, w_011_166);
  nand2 I024_116(w_024_116, w_008_268, w_017_321);
  or2  I024_117(w_024_117, w_020_610, w_008_592);
  and2 I024_118(w_024_118, w_002_699, w_017_410);
  or2  I024_119(w_024_119, w_004_256, w_002_629);
  not1 I024_120(w_024_120, w_011_121);
  and2 I024_121(w_024_121, w_014_099, w_013_171);
  or2  I024_122(w_024_122, w_001_004, w_008_409);
  or2  I024_123(w_024_123, w_018_011, w_011_142);
  not1 I024_125(w_024_125, w_010_487);
  nand2 I024_126(w_024_126, w_015_005, w_001_029);
  nand2 I024_127(w_024_127, w_012_050, w_011_130);
  and2 I024_128(w_024_128, w_001_005, w_017_242);
  nand2 I024_129(w_024_129, w_002_651, w_004_036);
  not1 I024_130(w_024_130, w_007_178);
  or2  I024_133(w_024_133, w_015_357, w_011_072);
  nand2 I024_137(w_024_137, w_016_000, w_002_402);
  or2  I024_139(w_024_139, w_018_014, w_022_055);
  or2  I024_141(w_024_141, w_022_219, w_018_037);
  not1 I024_142(w_024_142, w_012_051);
  or2  I024_143(w_024_143, w_008_348, w_012_129);
  or2  I024_144(w_024_144, w_006_082, w_018_000);
  and2 I024_145(w_024_145, w_005_248, w_017_543);
  or2  I024_146(w_024_146, w_008_561, w_014_272);
  nand2 I024_151(w_024_151, w_000_143, w_012_189);
  nand2 I024_155(w_024_155, w_023_092, w_007_368);
  and2 I024_157(w_024_157, w_012_021, w_015_440);
  not1 I024_164(w_024_164, w_007_128);
  nand2 I024_166(w_024_166, w_009_512, w_022_310);
  nand2 I024_171(w_024_171, w_000_434, w_014_281);
  not1 I024_172(w_024_172, w_012_058);
  and2 I024_173(w_024_173, w_022_213, w_001_028);
  not1 I024_175(w_024_175, w_002_205);
  nand2 I024_176(w_024_176, w_017_447, w_007_306);
  not1 I024_178(w_024_178, w_007_190);
  and2 I024_180(w_024_180, w_003_017, w_018_013);
  and2 I024_181(w_024_181, w_004_179, w_001_001);
  nand2 I024_182(w_024_182, w_004_104, w_018_005);
  or2  I024_183(w_024_183, w_002_664, w_005_140);
  not1 I024_184(w_024_184, w_004_215);
  not1 I024_186(w_024_186, w_002_711);
  nand2 I024_187(w_024_187, w_005_184, w_001_011);
  and2 I024_188(w_024_188, w_021_236, w_021_122);
  not1 I024_189(w_024_189, w_017_211);
  and2 I024_190(w_024_190, w_023_024, w_018_017);
  not1 I024_191(w_024_191, w_021_179);
  not1 I024_192(w_024_192, w_005_048);
  not1 I024_193(w_024_193, w_019_011);
  not1 I024_194(w_024_194, w_017_125);
  not1 I024_195(w_024_195, w_016_004);
  not1 I024_197(w_024_197, w_006_029);
  not1 I024_200(w_024_200, w_005_054);
  or2  I024_202(w_024_202, w_009_247, w_010_059);
  and2 I024_205(w_024_205, w_011_211, w_022_295);
  nand2 I024_206(w_024_206, w_014_258, w_017_171);
  nand2 I024_207(w_024_207, w_017_438, w_009_328);
  nand2 I024_208(w_024_208, w_007_145, w_002_465);
  and2 I024_209(w_024_209, w_002_374, w_017_075);
  not1 I024_210(w_024_210, w_004_020);
  not1 I024_211(w_024_211, w_002_182);
  not1 I024_212(w_024_212, w_014_151);
  and2 I024_213(w_024_213, w_005_006, w_010_528);
  or2  I024_214(w_024_214, w_014_085, w_022_020);
  and2 I024_215(w_024_215, w_006_245, w_023_155);
  not1 I024_216(w_024_216, w_017_347);
  and2 I024_218(w_024_218, w_001_018, w_003_063);
  not1 I024_219(w_024_219, w_017_240);
  or2  I024_221(w_024_221, w_006_161, w_019_009);
  and2 I024_222(w_024_222, w_015_142, w_006_060);
  or2  I024_223(w_024_223, w_006_190, w_014_120);
  and2 I024_224(w_024_224, w_021_110, w_019_001);
  not1 I024_225(w_024_225, w_021_131);
  nand2 I024_227(w_024_227, w_017_009, w_020_039);
  nand2 I024_229(w_024_229, w_017_564, w_016_000);
  or2  I024_230(w_024_230, w_007_287, w_017_356);
  nand2 I024_231(w_024_231, w_013_123, w_013_034);
  or2  I024_243(w_024_243, w_013_122, w_008_735);
  nand2 I024_244(w_024_244, w_011_095, w_011_064);
  not1 I024_247(w_024_247, w_018_003);
  and2 I024_253(w_024_253, w_002_034, w_003_015);
  and2 I024_254(w_024_254, w_014_104, w_008_595);
  and2 I024_257(w_024_257, w_007_026, w_010_288);
  or2  I024_258(w_024_258, w_023_148, w_010_518);
  or2  I024_260(w_024_260, w_023_143, w_010_567);
  not1 I024_262(w_024_262, w_013_195);
  or2  I024_263(w_024_263, w_017_443, w_003_040);
  not1 I024_265(w_024_265, w_012_011);
  not1 I024_268(w_024_268, w_005_087);
  nand2 I024_272(w_024_272, w_022_255, w_019_004);
  nand2 I024_273(w_024_273, w_022_304, w_009_122);
  and2 I024_275(w_024_275, w_012_038, w_006_145);
  not1 I024_276(w_024_276, w_007_219);
  or2  I024_277(w_024_277, w_011_338, w_021_044);
  and2 I024_280(w_024_280, w_002_622, w_022_102);
  or2  I024_283(w_024_283, w_002_553, w_008_399);
  not1 I024_284(w_024_284, w_019_002);
  or2  I024_286(w_024_286, w_011_057, w_014_022);
  not1 I024_292(w_024_292, w_001_029);
  not1 I024_295(w_024_295, w_015_016);
  or2  I024_299(w_024_299, w_008_623, w_011_504);
  nand2 I024_300(w_024_300, w_016_000, w_012_099);
  or2  I024_301(w_024_301, w_006_146, w_005_087);
  or2  I024_305(w_024_305, w_020_080, w_007_428);
  not1 I024_307(w_024_307, w_003_063);
  or2  I024_311(w_024_311, w_022_320, w_006_181);
  not1 I024_312(w_024_312, w_013_414);
  not1 I024_313(w_024_313, w_007_098);
  or2  I024_316(w_024_316, w_002_170, w_019_016);
  or2  I024_317(w_024_317, w_008_096, w_020_076);
  or2  I024_319(w_024_319, w_005_202, w_011_108);
  not1 I024_324(w_024_324, w_014_202);
  not1 I024_326(w_024_326, w_021_217);
  nand2 I024_327(w_024_327, w_008_541, w_008_647);
  and2 I024_329(w_024_329, w_014_284, w_006_208);
  nand2 I024_339(w_024_339, w_004_059, w_019_011);
  nand2 I024_342(w_024_342, w_015_665, w_005_210);
  or2  I024_346(w_024_346, w_006_108, w_007_218);
  or2  I024_347(w_024_347, w_014_226, w_000_478);
  and2 I024_354(w_024_354, w_020_123, w_012_171);
  and2 I024_355(w_024_355, w_023_018, w_005_248);
  nand2 I024_358(w_024_358, w_002_082, w_005_192);
  nand2 I024_359(w_024_359, w_012_340, w_021_010);
  and2 I024_361(w_024_361, w_004_101, w_009_049);
  not1 I024_365(w_024_365, w_005_303);
  nand2 I024_367(w_024_367, w_023_044, w_008_715);
  or2  I024_369(w_024_369, w_022_144, w_005_207);
  or2  I024_371(w_024_371, w_016_005, w_023_012);
  not1 I024_372(w_024_372, w_010_217);
  and2 I024_373(w_024_373, w_002_141, w_019_019);
  not1 I024_377(w_024_377, w_013_116);
  and2 I024_378(w_024_378, w_021_181, w_012_088);
  nand2 I024_386(w_024_386, w_021_127, w_007_064);
  or2  I024_387(w_024_387, w_002_041, w_013_256);
  not1 I024_388(w_024_388, w_022_344);
  and2 I024_389(w_024_389, w_022_214, w_012_126);
  not1 I024_391(w_024_391, w_022_081);
  not1 I024_392(w_024_392, w_003_067);
  not1 I024_395(w_024_395, w_008_169);
  and2 I024_399(w_024_399, w_017_189, w_001_034);
  and2 I024_401(w_024_401, w_010_763, w_007_050);
  and2 I024_404(w_024_404, w_007_454, w_002_158);
  or2  I024_411(w_024_411, w_004_394, w_007_042);
  not1 I024_413(w_024_413, w_012_000);
  and2 I024_418(w_024_418, w_002_561, w_011_372);
  nand2 I024_419(w_024_419, w_004_247, w_014_215);
  not1 I024_421(w_024_421, w_005_014);
  or2  I024_422(w_024_422, w_013_158, w_018_021);
  and2 I024_424(w_024_424, w_014_081, w_018_012);
  not1 I024_426(w_024_426, w_015_023);
  or2  I024_430(w_024_430, w_010_149, w_013_016);
  or2  I024_433(w_024_433, w_000_426, w_012_127);
  not1 I024_434(w_024_434, w_007_043);
  and2 I024_435(w_024_435, w_015_259, w_004_157);
  not1 I024_436(w_024_436, w_018_005);
  nand2 I024_439(w_024_439, w_000_208, w_019_008);
  nand2 I024_441(w_024_441, w_004_286, w_012_203);
  not1 I024_444(w_024_444, w_017_257);
  or2  I024_445(w_024_445, w_014_205, w_020_134);
  or2  I024_447(w_024_447, w_011_036, w_001_027);
  and2 I024_452(w_024_452, w_001_023, w_013_392);
  or2  I024_456(w_024_456, w_003_059, w_008_030);
  or2  I024_457(w_024_457, w_023_020, w_000_703);
  and2 I024_461(w_024_461, w_008_699, w_010_672);
  nand2 I024_464(w_024_464, w_014_104, w_013_422);
  not1 I024_473(w_024_473, w_002_059);
  not1 I024_477(w_024_477, w_018_020);
  not1 I024_478(w_024_478, w_014_102);
  not1 I024_481(w_024_481, w_022_323);
  not1 I024_482(w_024_482, w_006_001);
  or2  I024_483(w_024_483, w_007_261, w_018_006);
  or2  I024_489(w_024_489, w_016_003, w_002_504);
  nand2 I024_491(w_024_491, w_003_050, w_019_005);
  nand2 I024_492(w_024_492, w_009_251, w_014_126);
  or2  I024_493(w_024_493, w_002_257, w_001_013);
  nand2 I024_496(w_024_496, w_006_243, w_013_542);
  and2 I024_499(w_024_499, w_017_402, w_021_259);
  and2 I024_503(w_024_503, w_017_051, w_023_207);
  nand2 I024_506(w_024_506, w_010_196, w_011_360);
  not1 I024_507(w_024_507, w_007_045);
  not1 I024_509(w_024_509, w_015_058);
  not1 I024_510(w_024_510, w_008_461);
  or2  I024_513(w_024_513, w_008_221, w_011_041);
  and2 I024_516(w_024_516, w_008_199, w_002_504);
  and2 I024_517(w_024_517, w_020_067, w_022_298);
  not1 I024_518(w_024_518, w_013_309);
  or2  I024_521(w_024_521, w_009_362, w_010_716);
  nand2 I024_523(w_024_523, w_001_036, w_010_201);
  nand2 I024_524(w_024_524, w_022_084, w_018_022);
  not1 I024_525(w_024_525, w_007_423);
  and2 I024_528(w_024_528, w_022_033, w_014_250);
  or2  I024_530(w_024_530, w_021_174, w_003_010);
  nand2 I024_534(w_024_534, w_020_065, w_011_339);
  and2 I024_535(w_024_535, w_017_086, w_016_004);
  nand2 I024_537(w_024_537, w_005_056, w_001_011);
  nand2 I024_541(w_024_541, w_013_004, w_005_134);
  or2  I024_542(w_024_542, w_021_183, w_013_158);
  and2 I024_545(w_024_545, w_015_523, w_000_207);
  or2  I024_549(w_024_549, w_011_118, w_019_015);
  nand2 I024_551(w_024_551, w_009_463, w_003_070);
  nand2 I024_557(w_024_557, w_012_227, w_020_465);
  not1 I024_558(w_024_558, w_005_161);
  not1 I024_559(w_024_559, w_013_219);
  nand2 I024_563(w_024_563, w_016_006, w_015_072);
  not1 I024_565(w_024_565, w_009_162);
  nand2 I024_566(w_024_566, w_017_144, w_017_085);
  nand2 I024_569(w_024_569, w_010_525, w_023_020);
  nand2 I024_571(w_024_571, w_004_487, w_019_000);
  nand2 I024_574(w_024_574, w_001_004, w_013_169);
  or2  I024_577(w_024_577, w_006_020, w_013_401);
  and2 I024_579(w_024_579, w_016_008, w_022_357);
  not1 I024_580(w_024_582, w_024_581);
  or2  I024_581(w_024_583, w_006_258, w_024_582);
  or2  I024_582(w_024_584, w_024_599, w_024_583);
  not1 I024_583(w_024_585, w_024_584);
  nand2 I024_584(w_024_586, w_024_585, w_021_195);
  and2 I024_585(w_024_587, w_021_146, w_024_586);
  not1 I024_586(w_024_581, w_024_587);
  nand2 I024_587(w_024_592, w_024_591, w_010_635);
  not1 I024_588(w_024_593, w_024_592);
  not1 I024_589(w_024_594, w_024_593);
  nand2 I024_590(w_024_595, w_021_115, w_024_594);
  nand2 I024_591(w_024_596, w_024_595, w_013_188);
  and2 I024_592(w_024_597, w_024_596, w_023_027);
  not1 I024_593(w_024_591, w_024_584);
  and2 I024_594(w_024_599, w_013_199, w_024_597);
  not1 I025_000(w_025_000, w_018_012);
  nand2 I025_001(w_025_001, w_021_246, w_008_036);
  not1 I025_002(w_025_002, w_016_005);
  and2 I025_003(w_025_003, w_014_225, w_010_049);
  and2 I025_004(w_025_004, w_009_126, w_012_332);
  or2  I025_005(w_025_005, w_010_166, w_014_025);
  not1 I025_006(w_025_006, w_016_002);
  not1 I025_007(w_025_007, w_000_448);
  not1 I025_008(w_025_008, w_022_249);
  and2 I025_009(w_025_009, w_020_320, w_006_239);
  and2 I025_010(w_025_010, w_014_183, w_000_638);
  nand2 I025_011(w_025_011, w_002_174, w_024_128);
  nand2 I025_012(w_025_012, w_006_055, w_022_024);
  not1 I025_013(w_025_013, w_018_023);
  nand2 I025_015(w_025_015, w_016_006, w_000_513);
  and2 I025_016(w_025_016, w_007_459, w_007_396);
  and2 I025_018(w_025_018, w_002_367, w_021_235);
  or2  I025_019(w_025_019, w_020_260, w_007_289);
  not1 I025_021(w_025_021, w_009_058);
  not1 I025_023(w_025_023, w_019_013);
  not1 I025_024(w_025_024, w_015_401);
  nand2 I025_025(w_025_025, w_001_004, w_023_073);
  not1 I025_026(w_025_026, w_018_040);
  or2  I025_027(w_025_027, w_024_051, w_006_152);
  and2 I025_028(w_025_028, w_001_009, w_020_016);
  nand2 I025_029(w_025_029, w_015_644, w_019_009);
  or2  I025_032(w_025_032, w_018_012, w_013_327);
  not1 I025_034(w_025_034, w_006_067);
  not1 I025_035(w_025_035, w_010_428);
  and2 I025_036(w_025_036, w_017_059, w_019_015);
  not1 I025_037(w_025_037, w_006_066);
  not1 I025_038(w_025_038, w_009_169);
  nand2 I025_039(w_025_039, w_014_092, w_000_452);
  and2 I025_040(w_025_040, w_020_592, w_008_696);
  nand2 I025_042(w_025_042, w_007_248, w_003_084);
  not1 I025_043(w_025_043, w_006_168);
  not1 I025_044(w_025_044, w_017_087);
  not1 I025_048(w_025_048, w_017_119);
  nand2 I025_049(w_025_049, w_019_007, w_008_428);
  nand2 I025_050(w_025_050, w_015_606, w_011_057);
  and2 I025_051(w_025_051, w_006_191, w_006_070);
  and2 I025_053(w_025_053, w_002_475, w_023_062);
  or2  I025_054(w_025_054, w_024_107, w_007_236);
  or2  I025_055(w_025_055, w_019_000, w_017_352);
  and2 I025_056(w_025_056, w_012_217, w_002_025);
  or2  I025_057(w_025_057, w_016_006, w_021_150);
  or2  I025_059(w_025_059, w_004_281, w_021_256);
  not1 I025_060(w_025_060, w_020_011);
  and2 I025_061(w_025_061, w_021_250, w_021_114);
  and2 I025_062(w_025_062, w_015_254, w_022_009);
  nand2 I025_063(w_025_063, w_011_539, w_002_338);
  or2  I025_064(w_025_064, w_018_029, w_013_170);
  nand2 I025_066(w_025_066, w_015_568, w_017_660);
  and2 I025_067(w_025_067, w_006_056, w_007_220);
  and2 I025_069(w_025_069, w_002_574, w_003_059);
  not1 I025_072(w_025_072, w_002_503);
  not1 I025_073(w_025_073, w_017_272);
  and2 I025_074(w_025_074, w_005_085, w_024_133);
  not1 I025_075(w_025_075, w_001_029);
  or2  I025_076(w_025_076, w_022_356, w_016_002);
  not1 I025_077(w_025_077, w_018_015);
  or2  I025_078(w_025_078, w_005_095, w_004_016);
  not1 I025_079(w_025_079, w_001_025);
  and2 I025_080(w_025_080, w_004_066, w_024_280);
  and2 I025_081(w_025_081, w_021_098, w_000_052);
  not1 I025_082(w_025_082, w_014_093);
  not1 I025_083(w_025_083, w_002_695);
  nand2 I025_084(w_025_084, w_018_012, w_009_616);
  not1 I025_086(w_025_086, w_003_045);
  nand2 I025_088(w_025_088, w_011_024, w_013_175);
  or2  I025_089(w_025_089, w_015_333, w_015_057);
  not1 I025_092(w_025_092, w_011_641);
  and2 I025_093(w_025_093, w_017_312, w_020_094);
  nand2 I025_094(w_025_094, w_001_010, w_018_015);
  not1 I025_095(w_025_095, w_008_424);
  nand2 I025_096(w_025_096, w_023_092, w_018_027);
  or2  I025_097(w_025_097, w_011_162, w_005_111);
  or2  I025_098(w_025_098, w_024_099, w_003_044);
  or2  I025_099(w_025_099, w_017_565, w_000_209);
  or2  I025_100(w_025_100, w_022_245, w_007_225);
  or2  I025_101(w_025_101, w_000_690, w_010_383);
  nand2 I025_102(w_025_102, w_013_183, w_002_583);
  or2  I025_103(w_025_103, w_022_361, w_005_283);
  and2 I025_104(w_025_104, w_012_253, w_003_070);
  or2  I025_105(w_025_105, w_007_382, w_020_091);
  nand2 I025_106(w_025_106, w_024_579, w_024_457);
  nand2 I025_108(w_025_108, w_014_110, w_003_036);
  or2  I025_110(w_025_110, w_004_020, w_010_668);
  or2  I025_111(w_025_111, w_014_108, w_005_279);
  nand2 I025_112(w_025_112, w_000_505, w_013_574);
  and2 I025_113(w_025_113, w_012_231, w_017_546);
  nand2 I025_114(w_025_114, w_014_093, w_013_105);
  or2  I025_115(w_025_115, w_018_036, w_016_006);
  not1 I025_116(w_025_116, w_004_123);
  not1 I025_117(w_025_117, w_014_197);
  nand2 I025_118(w_025_118, w_005_132, w_014_131);
  not1 I025_119(w_025_119, w_016_008);
  or2  I025_120(w_025_120, w_016_007, w_024_574);
  not1 I025_121(w_025_121, w_020_169);
  or2  I025_122(w_025_122, w_012_056, w_013_127);
  and2 I025_123(w_025_123, w_011_002, w_020_109);
  not1 I025_124(w_025_124, w_018_021);
  and2 I025_125(w_025_125, w_011_571, w_005_099);
  or2  I025_126(w_025_126, w_009_154, w_004_244);
  or2  I025_127(w_025_127, w_022_118, w_020_023);
  and2 I025_130(w_025_130, w_023_031, w_003_066);
  or2  I025_131(w_025_131, w_001_033, w_009_481);
  nand2 I025_132(w_025_132, w_021_042, w_003_017);
  or2  I025_133(w_025_133, w_024_424, w_009_271);
  and2 I025_134(w_025_134, w_022_239, w_016_004);
  not1 I025_135(w_025_135, w_018_010);
  not1 I025_137(w_025_137, w_013_514);
  nand2 I025_138(w_025_138, w_016_007, w_000_500);
  not1 I025_139(w_025_139, w_024_292);
  or2  I025_140(w_025_140, w_001_015, w_018_021);
  and2 I025_141(w_025_141, w_015_201, w_014_059);
  not1 I025_142(w_025_142, w_009_126);
  nand2 I025_143(w_025_143, w_014_193, w_011_018);
  and2 I025_145(w_025_145, w_006_034, w_017_581);
  nand2 I025_147(w_025_147, w_019_009, w_001_007);
  nand2 I025_148(w_025_148, w_016_003, w_020_075);
  nand2 I025_149(w_025_149, w_009_064, w_011_146);
  not1 I025_151(w_025_151, w_004_270);
  not1 I025_152(w_025_152, w_012_325);
  not1 I025_154(w_025_154, w_020_311);
  nand2 I025_155(w_025_155, w_004_382, w_007_381);
  not1 I025_157(w_025_157, w_005_280);
  or2  I025_158(w_025_158, w_015_215, w_020_036);
  not1 I025_160(w_025_160, w_008_654);
  nand2 I025_161(w_025_161, w_002_599, w_011_123);
  not1 I025_162(w_025_162, w_024_326);
  nand2 I025_163(w_025_163, w_006_182, w_011_024);
  and2 I025_164(w_025_164, w_010_434, w_001_000);
  and2 I025_165(w_025_165, w_018_011, w_013_379);
  nand2 I025_166(w_025_166, w_022_349, w_011_465);
  nand2 I025_167(w_025_167, w_019_004, w_002_173);
  nand2 I025_168(w_025_168, w_015_491, w_016_003);
  or2  I025_169(w_025_169, w_021_147, w_005_095);
  not1 I025_170(w_025_170, w_003_013);
  and2 I025_171(w_025_171, w_006_005, w_002_050);
  nand2 I025_172(w_025_172, w_015_429, w_011_047);
  nand2 I025_173(w_025_173, w_022_355, w_005_105);
  not1 I025_174(w_025_174, w_009_468);
  or2  I025_176(w_025_176, w_010_139, w_011_168);
  or2  I025_177(w_025_177, w_014_061, w_022_235);
  not1 I025_178(w_025_178, w_024_115);
  not1 I025_179(w_025_179, w_017_006);
  or2  I025_180(w_025_180, w_007_208, w_012_088);
  not1 I025_181(w_025_181, w_007_183);
  and2 I025_182(w_025_182, w_000_211, w_001_024);
  and2 I025_184(w_025_184, w_004_086, w_015_318);
  and2 I025_186(w_025_186, w_008_590, w_013_037);
  nand2 I025_187(w_025_187, w_022_187, w_019_015);
  and2 I025_188(w_025_188, w_001_020, w_015_478);
  not1 I025_189(w_025_189, w_018_015);
  nand2 I025_191(w_025_191, w_009_089, w_024_354);
  or2  I025_192(w_025_192, w_012_292, w_010_248);
  nand2 I025_194(w_025_194, w_012_212, w_023_080);
  not1 I025_199(w_025_199, w_018_011);
  not1 I025_201(w_025_201, w_006_025);
  or2  I025_202(w_025_202, w_022_175, w_023_065);
  not1 I025_204(w_025_204, w_012_027);
  not1 I025_205(w_025_205, w_001_027);
  not1 I025_207(w_025_207, w_019_001);
  or2  I025_209(w_025_209, w_001_007, w_007_003);
  or2  I025_210(w_025_210, w_001_000, w_019_016);
  nand2 I025_211(w_025_211, w_003_056, w_007_258);
  or2  I025_216(w_025_216, w_024_369, w_016_003);
  and2 I025_217(w_025_217, w_012_072, w_009_244);
  or2  I025_218(w_025_218, w_013_555, w_011_465);
  nand2 I025_219(w_025_219, w_023_122, w_000_159);
  and2 I025_221(w_025_221, w_012_060, w_018_033);
  nand2 I025_222(w_025_222, w_001_028, w_000_492);
  nand2 I025_223(w_025_223, w_005_156, w_022_131);
  or2  I025_227(w_025_227, w_009_232, w_013_404);
  nand2 I025_228(w_025_228, w_019_012, w_014_201);
  or2  I025_229(w_025_229, w_012_076, w_008_561);
  nand2 I025_231(w_025_231, w_023_141, w_003_036);
  and2 I025_233(w_025_233, w_012_209, w_009_601);
  or2  I025_234(w_025_234, w_020_495, w_021_061);
  not1 I025_235(w_025_235, w_023_189);
  not1 I025_236(w_025_236, w_006_134);
  not1 I025_239(w_025_239, w_002_007);
  nand2 I025_240(w_025_240, w_002_096, w_020_045);
  or2  I025_241(w_025_241, w_023_161, w_002_569);
  or2  I025_242(w_025_242, w_013_163, w_000_413);
  or2  I025_243(w_025_243, w_006_099, w_024_171);
  or2  I025_247(w_025_247, w_019_010, w_020_221);
  nand2 I025_249(w_025_249, w_021_056, w_006_146);
  nand2 I025_251(w_025_251, w_001_000, w_016_007);
  and2 I025_253(w_025_253, w_012_215, w_013_126);
  nand2 I025_257(w_025_257, w_003_031, w_012_044);
  not1 I025_258(w_025_258, w_005_081);
  nand2 I025_261(w_025_261, w_017_019, w_021_249);
  and2 I025_263(w_025_263, w_011_310, w_018_034);
  and2 I025_264(w_025_264, w_007_163, w_014_212);
  and2 I025_265(w_025_265, w_023_104, w_001_010);
  not1 I025_269(w_025_269, w_018_038);
  and2 I025_271(w_025_271, w_015_632, w_008_439);
  and2 I025_272(w_025_272, w_009_408, w_009_284);
  and2 I025_277(w_025_277, w_001_008, w_021_194);
  or2  I025_279(w_025_279, w_015_004, w_001_004);
  not1 I025_280(w_025_280, w_002_414);
  or2  I025_281(w_025_281, w_009_059, w_003_082);
  nand2 I025_282(w_025_282, w_020_063, w_014_062);
  not1 I025_283(w_025_283, w_015_103);
  or2  I025_287(w_025_287, w_006_219, w_014_193);
  or2  I025_288(w_025_288, w_005_181, w_008_519);
  not1 I025_290(w_025_290, w_009_233);
  nand2 I025_291(w_025_291, w_015_363, w_020_393);
  and2 I025_294(w_025_294, w_015_369, w_005_277);
  and2 I025_296(w_025_296, w_005_316, w_020_453);
  or2  I025_297(w_025_297, w_008_015, w_020_341);
  or2  I025_303(w_025_303, w_010_263, w_004_083);
  not1 I025_304(w_025_304, w_002_135);
  and2 I025_305(w_025_305, w_017_392, w_011_525);
  nand2 I025_306(w_025_306, w_009_235, w_019_007);
  nand2 I025_307(w_025_307, w_004_259, w_022_319);
  nand2 I025_308(w_025_308, w_015_658, w_007_395);
  and2 I025_309(w_024_589, w_017_093, w_024_581);
  and2 I026_000(w_026_000, w_009_210, w_024_372);
  not1 I026_002(w_026_002, w_008_434);
  nand2 I026_004(w_026_004, w_010_597, w_021_009);
  not1 I026_005(w_026_005, w_016_002);
  and2 I026_006(w_026_006, w_013_138, w_010_407);
  or2  I026_007(w_026_007, w_017_131, w_016_006);
  or2  I026_008(w_026_008, w_018_030, w_003_030);
  not1 I026_009(w_026_009, w_005_088);
  not1 I026_010(w_026_010, w_014_191);
  nand2 I026_012(w_026_012, w_021_177, w_002_406);
  nand2 I026_013(w_026_013, w_015_328, w_007_010);
  nand2 I026_015(w_026_015, w_015_258, w_002_013);
  not1 I026_018(w_026_018, w_025_036);
  and2 I026_023(w_026_023, w_025_188, w_019_014);
  and2 I026_025(w_026_025, w_008_277, w_017_613);
  and2 I026_026(w_026_026, w_007_071, w_025_179);
  and2 I026_027(w_026_027, w_005_270, w_005_098);
  nand2 I026_028(w_026_028, w_000_378, w_016_002);
  not1 I026_033(w_026_033, w_013_536);
  or2  I026_038(w_026_038, w_012_253, w_024_181);
  and2 I026_039(w_026_039, w_000_154, w_008_587);
  not1 I026_042(w_026_042, w_006_218);
  and2 I026_044(w_026_044, w_014_122, w_002_050);
  nand2 I026_045(w_026_045, w_016_008, w_005_027);
  not1 I026_048(w_026_048, w_007_067);
  and2 I026_049(w_026_049, w_020_447, w_000_343);
  or2  I026_050(w_026_050, w_014_198, w_015_013);
  not1 I026_051(w_026_051, w_003_062);
  or2  I026_055(w_026_055, w_024_065, w_022_311);
  not1 I026_056(w_026_056, w_006_232);
  nand2 I026_058(w_026_058, w_006_163, w_004_348);
  not1 I026_059(w_026_059, w_005_103);
  or2  I026_060(w_026_060, w_013_528, w_010_452);
  or2  I026_061(w_026_061, w_024_122, w_023_193);
  or2  I026_064(w_026_064, w_002_646, w_018_039);
  and2 I026_067(w_026_067, w_006_023, w_014_121);
  not1 I026_068(w_026_068, w_002_311);
  not1 I026_070(w_026_070, w_013_053);
  nand2 I026_071(w_026_071, w_017_484, w_015_020);
  and2 I026_072(w_026_072, w_013_332, w_010_442);
  not1 I026_074(w_026_074, w_008_581);
  not1 I026_076(w_026_076, w_004_163);
  and2 I026_077(w_026_077, w_016_005, w_021_207);
  or2  I026_082(w_026_082, w_012_257, w_006_002);
  and2 I026_088(w_026_088, w_000_541, w_023_188);
  or2  I026_090(w_026_090, w_016_007, w_010_211);
  and2 I026_092(w_026_092, w_021_192, w_013_016);
  or2  I026_093(w_026_093, w_016_001, w_015_043);
  nand2 I026_098(w_026_098, w_006_065, w_005_051);
  nand2 I026_105(w_026_105, w_015_467, w_002_688);
  or2  I026_107(w_026_107, w_019_010, w_019_019);
  nand2 I026_109(w_026_109, w_009_009, w_011_120);
  or2  I026_110(w_026_110, w_010_118, w_025_027);
  not1 I026_112(w_026_112, w_020_062);
  or2  I026_113(w_026_113, w_001_004, w_010_216);
  or2  I026_114(w_026_114, w_005_236, w_008_351);
  not1 I026_115(w_026_115, w_021_204);
  or2  I026_117(w_026_117, w_021_248, w_002_536);
  and2 I026_118(w_026_118, w_004_479, w_012_153);
  or2  I026_121(w_026_121, w_008_728, w_008_271);
  nand2 I026_122(w_026_122, w_003_047, w_015_394);
  or2  I026_123(w_026_123, w_016_005, w_019_019);
  or2  I026_125(w_026_125, w_000_594, w_001_003);
  or2  I026_126(w_026_126, w_013_077, w_010_326);
  not1 I026_127(w_026_127, w_014_203);
  nand2 I026_128(w_026_128, w_024_200, w_007_145);
  or2  I026_130(w_026_130, w_007_268, w_003_020);
  not1 I026_132(w_026_132, w_011_551);
  and2 I026_136(w_026_136, w_019_017, w_019_014);
  and2 I026_139(w_026_139, w_005_266, w_025_122);
  not1 I026_140(w_026_140, w_006_103);
  nand2 I026_144(w_026_144, w_025_062, w_001_034);
  nand2 I026_145(w_026_145, w_022_066, w_001_027);
  not1 I026_146(w_026_146, w_000_708);
  and2 I026_149(w_026_149, w_019_013, w_016_002);
  or2  I026_152(w_026_152, w_017_499, w_025_077);
  not1 I026_154(w_026_154, w_023_082);
  or2  I026_160(w_026_160, w_000_194, w_009_379);
  and2 I026_161(w_026_161, w_002_013, w_003_081);
  and2 I026_163(w_026_163, w_019_018, w_009_141);
  and2 I026_169(w_026_169, w_000_177, w_011_144);
  nand2 I026_172(w_026_172, w_009_183, w_020_177);
  and2 I026_173(w_026_173, w_016_006, w_002_013);
  or2  I026_174(w_026_174, w_002_316, w_016_008);
  and2 I026_178(w_026_178, w_008_745, w_012_181);
  and2 I026_179(w_026_179, w_006_205, w_023_017);
  nand2 I026_181(w_026_181, w_005_259, w_017_248);
  and2 I026_182(w_026_182, w_003_067, w_012_135);
  not1 I026_184(w_026_184, w_012_069);
  and2 I026_187(w_026_187, w_004_184, w_019_019);
  nand2 I026_188(w_026_188, w_024_218, w_019_012);
  not1 I026_189(w_026_189, w_022_251);
  nand2 I026_191(w_026_191, w_022_076, w_010_343);
  nand2 I026_192(w_026_192, w_005_150, w_012_125);
  or2  I026_193(w_026_193, w_006_102, w_020_180);
  and2 I026_196(w_026_196, w_003_011, w_002_069);
  nand2 I026_198(w_026_198, w_003_067, w_003_024);
  or2  I026_201(w_026_201, w_013_159, w_023_161);
  and2 I026_211(w_026_211, w_019_016, w_017_338);
  or2  I026_216(w_026_216, w_014_249, w_001_018);
  or2  I026_217(w_026_217, w_005_247, w_012_340);
  or2  I026_223(w_026_223, w_013_562, w_005_072);
  and2 I026_224(w_026_224, w_024_589, w_020_411);
  or2  I026_225(w_026_225, w_006_106, w_011_136);
  or2  I026_226(w_026_226, w_012_043, w_000_754);
  and2 I026_227(w_026_227, w_025_207, w_008_749);
  nand2 I026_229(w_026_229, w_005_160, w_015_144);
  not1 I026_231(w_026_231, w_015_263);
  nand2 I026_234(w_026_234, w_009_055, w_009_120);
  and2 I026_237(w_026_237, w_003_025, w_001_009);
  nand2 I026_238(w_026_238, w_008_130, w_015_458);
  or2  I026_239(w_026_239, w_011_492, w_001_009);
  nand2 I026_250(w_026_250, w_013_518, w_005_153);
  and2 I026_257(w_026_257, w_017_012, w_023_121);
  nand2 I026_261(w_026_261, w_020_290, w_020_356);
  not1 I026_267(w_026_267, w_024_077);
  not1 I026_268(w_026_268, w_019_016);
  and2 I026_273(w_026_273, w_025_162, w_009_164);
  not1 I026_274(w_026_274, w_004_295);
  nand2 I026_275(w_026_275, w_016_004, w_012_350);
  nand2 I026_283(w_026_283, w_021_126, w_004_025);
  not1 I026_286(w_026_286, w_003_081);
  not1 I026_287(w_026_287, w_002_128);
  and2 I026_288(w_026_288, w_009_136, w_013_028);
  and2 I026_289(w_026_289, w_005_215, w_002_076);
  or2  I026_290(w_026_290, w_025_168, w_017_636);
  not1 I026_291(w_026_291, w_005_289);
  not1 I026_294(w_026_294, w_008_118);
  not1 I026_295(w_026_295, w_017_607);
  nand2 I026_296(w_026_296, w_021_192, w_012_204);
  nand2 I026_297(w_026_297, w_024_577, w_008_425);
  nand2 I026_298(w_026_298, w_019_018, w_008_574);
  or2  I026_299(w_026_299, w_019_005, w_012_054);
  or2  I026_304(w_026_304, w_010_489, w_014_182);
  and2 I026_305(w_026_305, w_009_603, w_006_161);
  or2  I026_310(w_026_310, w_008_310, w_012_271);
  not1 I026_311(w_026_311, w_008_209);
  or2  I026_315(w_026_315, w_004_030, w_020_529);
  and2 I026_317(w_026_317, w_002_654, w_014_209);
  and2 I026_321(w_026_321, w_008_683, w_001_012);
  or2  I026_322(w_026_322, w_021_040, w_005_089);
  or2  I026_326(w_026_326, w_012_091, w_002_496);
  or2  I026_328(w_026_328, w_019_008, w_000_703);
  or2  I026_331(w_026_331, w_021_152, w_003_077);
  and2 I026_332(w_026_332, w_012_311, w_015_652);
  not1 I026_333(w_026_333, w_019_008);
  not1 I026_343(w_026_343, w_000_041);
  nand2 I026_344(w_026_344, w_010_083, w_011_061);
  not1 I026_346(w_026_346, w_005_296);
  and2 I026_348(w_026_348, w_012_213, w_017_131);
  or2  I026_351(w_026_351, w_007_179, w_000_389);
  and2 I026_354(w_026_354, w_017_640, w_012_067);
  nand2 I026_357(w_026_357, w_024_173, w_005_124);
  nand2 I026_358(w_026_358, w_012_141, w_019_016);
  and2 I026_361(w_026_361, w_000_381, w_019_003);
  not1 I026_364(w_026_364, w_009_539);
  nand2 I026_366(w_026_366, w_002_178, w_018_014);
  or2  I026_371(w_026_371, w_007_295, w_002_056);
  nand2 I026_380(w_026_380, w_012_304, w_017_022);
  or2  I026_381(w_026_381, w_023_202, w_022_291);
  and2 I026_382(w_026_382, w_011_087, w_023_065);
  and2 I026_383(w_026_383, w_010_419, w_014_182);
  not1 I026_393(w_026_393, w_000_355);
  not1 I026_394(w_026_394, w_004_400);
  not1 I026_395(w_026_395, w_007_188);
  nand2 I026_396(w_026_396, w_019_020, w_012_019);
  not1 I026_400(w_026_400, w_014_059);
  or2  I026_404(w_026_404, w_018_002, w_001_021);
  and2 I026_410(w_026_410, w_010_583, w_003_013);
  or2  I026_411(w_026_411, w_004_223, w_022_193);
  and2 I026_413(w_026_413, w_018_034, w_022_277);
  and2 I026_415(w_026_415, w_023_141, w_002_302);
  or2  I026_420(w_026_420, w_021_118, w_019_014);
  nand2 I026_424(w_026_424, w_017_598, w_006_216);
  not1 I026_427(w_026_427, w_024_061);
  or2  I026_430(w_026_430, w_020_022, w_024_525);
  and2 I026_431(w_026_431, w_004_289, w_013_077);
  and2 I026_433(w_026_433, w_011_579, w_016_006);
  nand2 I026_439(w_026_439, w_005_090, w_021_189);
  and2 I026_441(w_026_441, w_003_010, w_020_430);
  nand2 I026_442(w_026_442, w_013_461, w_019_007);
  or2  I026_447(w_026_447, w_011_060, w_000_327);
  nand2 I026_448(w_026_448, w_020_447, w_004_007);
  or2  I026_449(w_026_449, w_015_082, w_024_042);
  not1 I026_451(w_026_451, w_018_003);
  or2  I026_453(w_026_453, w_019_002, w_018_039);
  nand2 I026_455(w_026_455, w_021_238, w_000_372);
  nand2 I026_457(w_026_457, w_000_756, w_015_033);
  and2 I026_459(w_026_459, w_019_011, w_024_137);
  not1 I026_466(w_026_466, w_007_115);
  or2  I026_471(w_026_471, w_024_422, w_004_215);
  nand2 I026_477(w_026_477, w_015_590, w_022_269);
  and2 I026_480(w_026_480, w_022_331, w_001_002);
  not1 I026_483(w_026_483, w_011_124);
  and2 I026_488(w_026_488, w_015_194, w_014_059);
  not1 I026_489(w_026_489, w_000_191);
  and2 I026_490(w_026_490, w_007_307, w_017_559);
  not1 I026_491(w_026_491, w_006_216);
  and2 I026_493(w_026_493, w_017_590, w_009_082);
  nand2 I026_494(w_026_494, w_012_214, w_019_019);
  not1 I026_499(w_026_499, w_001_034);
  and2 I026_500(w_026_500, w_013_102, w_024_439);
  and2 I026_502(w_026_502, w_019_013, w_007_049);
  nand2 I026_506(w_026_506, w_016_003, w_024_125);
  nand2 I026_507(w_026_507, w_013_363, w_015_308);
  nand2 I026_508(w_026_508, w_010_571, w_018_026);
  nand2 I026_513(w_026_513, w_015_134, w_003_016);
  or2  I026_514(w_026_514, w_017_271, w_004_125);
  not1 I026_515(w_026_515, w_017_248);
  nand2 I026_517(w_026_517, w_002_494, w_025_308);
  and2 I026_519(w_026_519, w_016_000, w_017_518);
  not1 I026_520(w_026_520, w_006_147);
  and2 I026_523(w_026_523, w_025_303, w_018_009);
  not1 I026_527(w_026_527, w_004_128);
  or2  I026_530(w_026_530, w_010_570, w_019_016);
  nand2 I026_531(w_026_531, w_016_003, w_007_090);
  nand2 I026_532(w_026_532, w_008_669, w_010_456);
  or2  I026_534(w_026_534, w_017_045, w_025_095);
  not1 I026_535(w_026_535, w_002_504);
  and2 I026_536(w_026_536, w_019_006, w_005_065);
  nand2 I026_538(w_026_538, w_012_101, w_008_580);
  not1 I026_539(w_026_539, w_020_588);
  nand2 I026_541(w_026_541, w_003_043, w_014_072);
  or2  I026_544(w_026_544, w_004_284, w_018_007);
  nand2 I026_548(w_026_548, w_016_008, w_023_087);
  or2  I026_549(w_026_549, w_015_651, w_001_025);
  or2  I026_550(w_026_550, w_008_484, w_005_168);
  and2 I026_551(w_026_551, w_023_053, w_001_012);
  and2 I026_555(w_026_555, w_001_007, w_013_468);
  and2 I026_561(w_026_561, w_024_059, w_012_145);
  nand2 I026_564(w_026_564, w_000_379, w_015_110);
  and2 I026_566(w_026_566, w_023_162, w_024_313);
  and2 I026_570(w_026_570, w_007_021, w_025_062);
  not1 I026_572(w_026_572, w_001_026);
  and2 I026_579(w_026_579, w_022_086, w_025_034);
  not1 I026_580(w_026_580, w_005_046);
  or2  I026_585(w_026_585, w_000_189, w_022_050);
  and2 I026_591(w_026_591, w_023_069, w_023_015);
  not1 I026_593(w_026_593, w_000_571);
  nand2 I026_595(w_026_595, w_016_001, w_003_043);
  and2 I026_597(w_026_597, w_002_669, w_004_413);
  and2 I026_598(w_026_598, w_001_006, w_016_006);
  and2 I026_600(w_026_600, w_018_030, w_019_005);
  nand2 I026_604(w_026_604, w_001_033, w_023_136);
  nand2 I026_605(w_026_605, w_015_107, w_020_305);
  nand2 I026_606(w_026_606, w_010_095, w_011_089);
  nand2 I026_608(w_026_608, w_006_085, w_016_005);
  or2  I026_613(w_026_613, w_024_110, w_024_215);
  and2 I026_614(w_026_614, w_005_302, w_004_181);
  and2 I026_617(w_026_617, w_024_200, w_025_151);
  or2  I026_620(w_026_620, w_008_640, w_004_235);
  and2 I026_621(w_026_621, w_009_056, w_020_036);
  not1 I026_630(w_026_630, w_016_006);
  and2 I026_632(w_026_632, w_014_029, w_002_478);
  nand2 I026_635(w_026_635, w_021_073, w_009_250);
  and2 I026_642(w_026_642, w_011_298, w_011_284);
  and2 I026_643(w_026_643, w_015_042, w_006_137);
  and2 I026_645(w_026_645, w_014_289, w_021_016);
  or2  I026_648(w_026_648, w_013_109, w_022_074);
  or2  I026_649(w_026_649, w_008_011, w_020_022);
  not1 I026_655(w_026_655, w_010_432);
  not1 I026_657(w_026_657, w_005_002);
  or2  I026_660(w_026_660, w_015_210, w_001_015);
  nand2 I026_661(w_026_661, w_016_005, w_022_300);
  or2  I026_662(w_026_662, w_008_284, w_009_391);
  not1 I026_663(w_026_663, w_001_013);
  nand2 I026_665(w_026_665, w_003_019, w_022_283);
  nand2 I026_668(w_026_668, w_002_337, w_007_171);
  or2  I026_669(w_026_669, w_016_006, w_001_002);
  not1 I026_670(w_026_670, w_002_234);
  and2 I026_675(w_026_675, w_016_008, w_007_087);
  not1 I026_681(w_026_681, w_024_430);
  nand2 I026_683(w_026_683, w_018_003, w_010_520);
  or2  I026_684(w_026_684, w_005_124, w_012_052);
  nand2 I026_687(w_026_687, w_002_019, w_003_024);
  and2 I026_692(w_026_692, w_019_019, w_012_264);
  or2  I026_693(w_026_693, w_017_506, w_009_525);
  or2  I026_694(w_026_694, w_012_008, w_002_285);
  not1 I026_695(w_026_695, w_005_195);
  or2  I026_698(w_026_698, w_024_491, w_025_049);
  and2 I026_699(w_026_699, w_013_313, w_000_738);
  and2 I026_701(w_026_701, w_016_007, w_000_197);
  and2 I026_702(w_026_702, w_024_034, w_018_040);
  or2  I026_703(w_026_703, w_024_022, w_004_083);
  not1 I026_705(w_026_705, w_017_024);
  and2 I026_706(w_026_706, w_019_003, w_004_418);
  nand2 I026_708(w_026_708, w_015_137, w_009_253);
  nand2 I026_709(w_026_709, w_003_010, w_016_005);
  not1 I026_711(w_026_711, w_017_613);
  and2 I026_712(w_026_712, w_014_172, w_011_329);
  not1 I026_718(w_026_718, w_001_010);
  not1 I026_720(w_026_720, w_019_005);
  nand2 I027_000(w_027_000, w_024_223, w_015_325);
  or2  I027_001(w_027_001, w_014_059, w_004_209);
  nand2 I027_002(w_027_002, w_016_001, w_023_203);
  and2 I027_004(w_027_004, w_024_062, w_022_390);
  not1 I027_006(w_027_006, w_005_010);
  or2  I027_007(w_027_007, w_009_024, w_017_337);
  nand2 I027_008(w_027_008, w_021_098, w_014_103);
  nand2 I027_009(w_027_009, w_010_670, w_021_102);
  nand2 I027_011(w_027_011, w_004_259, w_007_209);
  not1 I027_012(w_027_012, w_024_178);
  or2  I027_014(w_027_014, w_013_112, w_021_181);
  nand2 I027_015(w_027_015, w_005_313, w_014_043);
  nand2 I027_016(w_027_016, w_013_265, w_021_139);
  not1 I027_018(w_027_018, w_024_521);
  and2 I027_019(w_027_019, w_021_149, w_004_130);
  nand2 I027_020(w_027_020, w_008_097, w_025_086);
  and2 I027_023(w_027_023, w_016_002, w_004_406);
  nand2 I027_024(w_027_024, w_005_236, w_024_516);
  or2  I027_026(w_027_026, w_012_269, w_020_124);
  or2  I027_027(w_027_027, w_018_024, w_002_647);
  nand2 I027_028(w_027_028, w_024_411, w_015_099);
  and2 I027_030(w_027_030, w_001_010, w_009_074);
  nand2 I027_031(w_027_031, w_006_168, w_022_407);
  or2  I027_032(w_027_032, w_021_154, w_014_027);
  or2  I027_033(w_027_033, w_026_161, w_020_161);
  or2  I027_034(w_027_034, w_013_061, w_018_009);
  or2  I027_035(w_027_035, w_011_251, w_006_226);
  and2 I027_036(w_027_036, w_012_074, w_006_101);
  or2  I027_037(w_027_037, w_003_029, w_009_302);
  nand2 I027_039(w_027_039, w_001_033, w_019_006);
  not1 I027_040(w_027_040, w_012_305);
  nand2 I027_041(w_027_041, w_025_053, w_008_383);
  not1 I027_042(w_027_042, w_019_018);
  nand2 I027_043(w_027_043, w_017_038, w_017_121);
  or2  I027_044(w_027_044, w_016_000, w_004_115);
  nand2 I027_045(w_027_045, w_019_007, w_024_566);
  and2 I027_046(w_027_046, w_014_113, w_004_242);
  and2 I027_047(w_027_047, w_016_007, w_026_332);
  not1 I027_048(w_027_048, w_023_049);
  and2 I027_049(w_027_049, w_016_003, w_013_578);
  and2 I027_050(w_027_050, w_003_060, w_016_007);
  nand2 I027_051(w_027_051, w_020_348, w_023_156);
  or2  I027_053(w_027_053, w_023_147, w_024_359);
  nand2 I027_054(w_027_054, w_013_243, w_025_137);
  not1 I027_055(w_027_055, w_023_070);
  nand2 I027_056(w_027_056, w_009_019, w_022_305);
  nand2 I027_057(w_027_057, w_000_537, w_025_035);
  or2  I027_058(w_027_058, w_021_136, w_009_418);
  nand2 I027_059(w_027_059, w_017_260, w_007_287);
  nand2 I027_060(w_027_060, w_004_136, w_016_007);
  or2  I027_061(w_027_061, w_014_045, w_008_434);
  and2 I027_062(w_027_062, w_016_004, w_018_007);
  or2  I027_063(w_027_063, w_003_055, w_021_104);
  nand2 I027_064(w_027_064, w_024_401, w_011_267);
  nand2 I027_065(w_027_065, w_019_020, w_016_008);
  nand2 I027_066(w_027_066, w_016_003, w_024_182);
  not1 I027_067(w_027_067, w_012_207);
  and2 I027_068(w_027_068, w_021_091, w_002_018);
  nand2 I027_070(w_027_070, w_023_141, w_016_004);
  or2  I027_071(w_027_071, w_001_003, w_002_616);
  and2 I027_072(w_027_072, w_018_005, w_024_068);
  nand2 I027_073(w_027_073, w_021_162, w_011_189);
  or2  I027_074(w_027_074, w_021_073, w_020_055);
  not1 I027_075(w_027_075, w_010_609);
  not1 I027_076(w_027_076, w_012_149);
  not1 I027_077(w_027_077, w_024_496);
  and2 I027_078(w_027_078, w_006_192, w_000_305);
  not1 I027_079(w_027_079, w_026_113);
  not1 I027_080(w_027_080, w_013_536);
  not1 I027_081(w_027_081, w_009_270);
  or2  I027_082(w_027_082, w_009_011, w_022_404);
  nand2 I027_083(w_027_083, w_015_459, w_013_086);
  or2  I027_084(w_027_084, w_006_215, w_006_021);
  and2 I027_086(w_027_086, w_018_017, w_004_472);
  not1 I027_088(w_027_088, w_009_345);
  or2  I027_089(w_027_089, w_004_301, w_000_540);
  or2  I027_090(w_027_090, w_002_178, w_005_102);
  nand2 I027_091(w_027_091, w_000_442, w_005_122);
  and2 I027_092(w_027_092, w_008_138, w_025_093);
  and2 I027_093(w_027_093, w_002_565, w_020_514);
  or2  I027_094(w_027_094, w_007_120, w_022_010);
  or2  I027_095(w_027_095, w_014_090, w_002_350);
  not1 I027_096(w_027_096, w_024_491);
  and2 I027_097(w_027_097, w_018_022, w_018_025);
  nand2 I027_098(w_027_098, w_023_192, w_016_003);
  nand2 I027_099(w_027_099, w_014_222, w_019_009);
  nand2 I027_101(w_027_101, w_001_001, w_018_035);
  nand2 I027_102(w_027_102, w_020_520, w_009_516);
  and2 I027_103(w_027_103, w_009_130, w_013_361);
  and2 I027_104(w_027_104, w_010_757, w_020_131);
  not1 I027_105(w_027_105, w_025_074);
  nand2 I027_107(w_027_107, w_016_003, w_009_190);
  or2  I027_109(w_027_109, w_020_180, w_012_111);
  not1 I027_110(w_027_110, w_015_024);
  not1 I027_111(w_027_111, w_025_163);
  not1 I027_112(w_027_112, w_014_123);
  not1 I027_113(w_027_113, w_023_063);
  or2  I027_114(w_027_114, w_021_110, w_012_000);
  nand2 I027_115(w_027_115, w_002_479, w_014_037);
  nand2 I027_116(w_027_116, w_014_215, w_025_092);
  or2  I027_117(w_027_117, w_002_289, w_016_003);
  nand2 I027_118(w_027_118, w_013_027, w_000_294);
  or2  I027_119(w_027_119, w_003_034, w_013_053);
  nand2 I027_120(w_027_120, w_006_157, w_005_095);
  not1 I027_121(w_027_121, w_013_197);
  or2  I027_122(w_027_122, w_016_001, w_001_022);
  nand2 I027_123(w_027_123, w_015_010, w_020_158);
  or2  I027_124(w_027_124, w_010_707, w_015_374);
  not1 I027_125(w_027_125, w_015_668);
  nand2 I027_126(w_027_126, w_018_000, w_020_417);
  not1 I027_127(w_027_127, w_026_027);
  not1 I027_129(w_027_129, w_011_097);
  not1 I027_130(w_027_130, w_004_081);
  or2  I027_131(w_027_131, w_020_100, w_009_054);
  or2  I027_132(w_027_132, w_018_012, w_017_616);
  not1 I027_134(w_027_134, w_024_493);
  not1 I027_135(w_027_135, w_014_060);
  not1 I027_136(w_027_136, w_016_008);
  not1 I027_138(w_027_138, w_002_067);
  nand2 I027_139(w_027_139, w_008_258, w_018_011);
  and2 I027_140(w_027_140, w_002_536, w_017_142);
  and2 I027_141(w_027_141, w_009_487, w_009_032);
  or2  I027_142(w_027_142, w_000_152, w_011_576);
  not1 I027_143(w_027_143, w_000_244);
  nand2 I027_145(w_027_145, w_000_005, w_003_063);
  nand2 I027_146(w_027_146, w_021_239, w_015_384);
  not1 I027_148(w_027_148, w_025_249);
  and2 I027_149(w_027_149, w_015_401, w_006_175);
  nand2 I027_150(w_027_150, w_007_477, w_012_073);
  not1 I027_151(w_027_151, w_010_714);
  nand2 I027_153(w_027_153, w_000_726, w_012_259);
  and2 I027_155(w_027_155, w_018_033, w_023_143);
  nand2 I027_156(w_027_156, w_003_024, w_013_030);
  or2  I027_157(w_027_157, w_026_005, w_009_439);
  nand2 I027_158(w_027_158, w_012_067, w_026_239);
  not1 I027_159(w_027_159, w_023_113);
  or2  I027_160(w_027_160, w_008_724, w_010_242);
  not1 I027_161(w_027_161, w_003_006);
  nand2 I027_162(w_027_162, w_010_421, w_011_020);
  and2 I027_163(w_027_163, w_014_099, w_016_004);
  or2  I027_164(w_027_164, w_004_068, w_026_591);
  or2  I027_165(w_027_165, w_000_210, w_007_351);
  and2 I027_166(w_027_166, w_003_016, w_015_319);
  or2  I027_167(w_027_167, w_026_561, w_026_531);
  or2  I027_168(w_027_168, w_014_166, w_019_006);
  and2 I027_169(w_027_169, w_011_616, w_010_486);
  or2  I027_170(w_027_170, w_016_007, w_006_213);
  or2  I027_171(w_027_171, w_025_059, w_007_231);
  not1 I027_173(w_027_173, w_011_177);
  and2 I027_175(w_027_175, w_007_071, w_017_218);
  not1 I027_176(w_027_176, w_000_704);
  nand2 I027_177(w_027_177, w_016_002, w_000_270);
  and2 I027_178(w_027_178, w_014_147, w_003_074);
  nand2 I027_179(w_027_179, w_019_016, w_023_215);
  or2  I027_180(w_027_180, w_007_128, w_000_714);
  nand2 I027_181(w_027_181, w_015_042, w_022_198);
  nand2 I027_182(w_027_182, w_013_184, w_002_076);
  or2  I027_183(w_027_183, w_012_134, w_022_058);
  and2 I027_184(w_027_184, w_018_035, w_015_407);
  and2 I027_185(w_027_185, w_012_203, w_021_011);
  nand2 I027_187(w_027_187, w_001_000, w_012_169);
  nand2 I027_188(w_027_188, w_010_468, w_005_158);
  or2  I027_189(w_027_189, w_016_001, w_020_448);
  not1 I027_191(w_027_191, w_007_131);
  or2  I027_192(w_027_192, w_001_013, w_012_179);
  nand2 I027_194(w_027_194, w_000_757, w_012_346);
  and2 I027_195(w_027_195, w_017_408, w_004_200);
  or2  I027_197(w_027_197, w_006_018, w_025_038);
  not1 I027_198(w_027_198, w_021_182);
  or2  I027_199(w_027_199, w_022_054, w_017_017);
  and2 I027_202(w_027_202, w_000_461, w_008_278);
  not1 I027_204(w_027_204, w_012_142);
  not1 I028_000(w_028_000, w_000_291);
  not1 I028_001(w_028_001, w_013_236);
  and2 I028_003(w_028_003, w_001_036, w_021_121);
  and2 I028_005(w_028_005, w_009_105, w_020_339);
  and2 I028_006(w_028_006, w_017_561, w_018_020);
  not1 I028_008(w_028_008, w_019_000);
  nand2 I028_011(w_028_011, w_023_037, w_011_632);
  or2  I028_012(w_028_012, w_004_119, w_014_203);
  nand2 I028_013(w_028_013, w_003_084, w_013_025);
  not1 I028_014(w_028_014, w_001_007);
  and2 I028_018(w_028_018, w_010_505, w_025_120);
  and2 I028_021(w_028_021, w_005_228, w_007_085);
  and2 I028_022(w_028_022, w_018_014, w_024_054);
  nand2 I028_025(w_028_025, w_018_019, w_012_210);
  not1 I028_026(w_028_026, w_021_067);
  nand2 I028_027(w_028_027, w_027_180, w_003_070);
  or2  I028_028(w_028_028, w_020_034, w_012_143);
  not1 I028_029(w_028_029, w_002_285);
  not1 I028_030(w_028_030, w_008_419);
  and2 I028_033(w_028_033, w_006_102, w_020_183);
  not1 I028_034(w_028_034, w_018_020);
  nand2 I028_035(w_028_035, w_014_075, w_004_059);
  or2  I028_036(w_028_036, w_021_255, w_016_008);
  and2 I028_037(w_028_037, w_010_644, w_017_197);
  or2  I028_038(w_028_038, w_020_395, w_006_092);
  or2  I028_039(w_028_039, w_025_176, w_025_103);
  not1 I028_040(w_028_040, w_002_286);
  and2 I028_041(w_028_041, w_004_398, w_019_005);
  or2  I028_042(w_028_042, w_007_148, w_023_149);
  not1 I028_044(w_028_044, w_005_137);
  nand2 I028_045(w_028_045, w_002_088, w_019_004);
  and2 I028_050(w_028_050, w_018_004, w_027_084);
  or2  I028_052(w_028_052, w_003_025, w_020_521);
  nand2 I028_053(w_028_053, w_025_229, w_011_544);
  or2  I028_056(w_028_056, w_010_129, w_018_003);
  or2  I028_057(w_028_057, w_020_152, w_001_030);
  not1 I028_058(w_028_058, w_018_009);
  not1 I028_060(w_028_060, w_005_077);
  and2 I028_064(w_028_064, w_017_575, w_013_010);
  or2  I028_065(w_028_065, w_015_559, w_001_012);
  not1 I028_068(w_028_068, w_020_609);
  or2  I028_069(w_028_069, w_010_031, w_012_105);
  not1 I028_070(w_028_070, w_010_551);
  or2  I028_072(w_028_072, w_018_035, w_013_266);
  nand2 I028_074(w_028_074, w_002_028, w_025_114);
  or2  I028_076(w_028_076, w_015_033, w_013_464);
  and2 I028_077(w_028_077, w_008_567, w_007_071);
  nand2 I028_078(w_028_078, w_024_389, w_021_130);
  not1 I028_079(w_028_079, w_018_028);
  or2  I028_080(w_028_080, w_008_014, w_012_174);
  not1 I028_084(w_028_084, w_002_053);
  or2  I028_085(w_028_085, w_003_072, w_005_081);
  not1 I028_086(w_028_086, w_004_207);
  and2 I028_087(w_028_087, w_024_524, w_024_373);
  and2 I028_088(w_028_088, w_018_013, w_014_045);
  nand2 I028_089(w_028_089, w_001_029, w_001_033);
  nand2 I028_090(w_028_090, w_027_053, w_017_345);
  or2  I028_091(w_028_091, w_020_135, w_003_047);
  not1 I028_094(w_028_094, w_015_090);
  and2 I028_096(w_028_096, w_020_012, w_023_123);
  and2 I028_097(w_028_097, w_012_021, w_021_208);
  and2 I028_098(w_028_098, w_008_608, w_000_341);
  and2 I028_099(w_028_099, w_006_037, w_015_340);
  and2 I028_101(w_028_101, w_009_478, w_020_067);
  and2 I028_102(w_028_102, w_010_550, w_000_170);
  nand2 I028_104(w_028_104, w_008_188, w_003_055);
  and2 I028_105(w_028_105, w_003_033, w_004_117);
  nand2 I028_106(w_028_106, w_003_009, w_022_315);
  nand2 I028_107(w_028_107, w_026_090, w_001_002);
  and2 I028_109(w_028_109, w_013_191, w_019_003);
  or2  I028_110(w_028_110, w_018_042, w_012_093);
  nand2 I028_111(w_028_111, w_015_112, w_015_202);
  or2  I028_113(w_028_113, w_006_075, w_003_002);
  and2 I028_115(w_028_115, w_005_067, w_008_730);
  not1 I028_117(w_028_117, w_019_010);
  or2  I028_118(w_028_118, w_006_183, w_017_018);
  nand2 I028_119(w_028_119, w_020_208, w_005_196);
  or2  I028_120(w_028_120, w_020_142, w_000_126);
  and2 I028_121(w_028_121, w_005_260, w_024_010);
  and2 I028_122(w_028_122, w_005_293, w_021_257);
  nand2 I028_123(w_028_123, w_000_039, w_021_221);
  not1 I028_125(w_028_125, w_010_168);
  nand2 I028_126(w_028_126, w_027_068, w_012_072);
  not1 I028_127(w_028_127, w_024_102);
  not1 I028_128(w_028_128, w_001_011);
  nand2 I028_129(w_028_129, w_024_137, w_016_007);
  nand2 I028_130(w_028_130, w_005_293, w_003_018);
  not1 I028_131(w_028_131, w_006_191);
  or2  I028_132(w_028_132, w_027_103, w_005_071);
  not1 I028_133(w_028_133, w_017_497);
  or2  I028_134(w_028_134, w_013_013, w_020_595);
  or2  I028_135(w_028_135, w_014_289, w_011_043);
  and2 I028_136(w_028_136, w_019_019, w_020_144);
  and2 I028_137(w_028_137, w_009_124, w_003_075);
  nand2 I028_139(w_028_139, w_020_087, w_020_158);
  or2  I028_140(w_028_140, w_010_471, w_026_223);
  and2 I028_141(w_028_141, w_003_030, w_022_011);
  nand2 I028_142(w_028_142, w_005_017, w_012_090);
  not1 I028_143(w_028_143, w_004_304);
  not1 I028_144(w_028_144, w_014_131);
  or2  I028_145(w_028_145, w_016_003, w_006_118);
  nand2 I028_147(w_028_147, w_005_061, w_009_516);
  nand2 I028_149(w_028_149, w_007_077, w_008_636);
  or2  I028_150(w_028_150, w_016_005, w_010_000);
  and2 I028_151(w_028_151, w_008_428, w_009_150);
  nand2 I028_152(w_028_152, w_015_351, w_018_008);
  nand2 I028_154(w_028_154, w_026_211, w_022_098);
  or2  I028_156(w_028_156, w_019_007, w_027_139);
  nand2 I028_160(w_028_160, w_026_517, w_010_724);
  not1 I028_162(w_028_162, w_020_015);
  and2 I028_163(w_028_163, w_012_111, w_023_007);
  or2  I028_165(w_028_165, w_017_267, w_021_110);
  not1 I028_170(w_028_170, w_003_037);
  not1 I028_171(w_028_171, w_026_595);
  or2  I028_173(w_028_173, w_009_584, w_020_083);
  and2 I028_175(w_028_175, w_014_027, w_014_072);
  or2  I028_177(w_028_177, w_003_033, w_025_042);
  nand2 I028_178(w_028_178, w_009_564, w_002_580);
  or2  I028_181(w_028_181, w_026_351, w_010_120);
  nand2 I028_182(w_028_182, w_024_489, w_004_187);
  or2  I028_183(w_028_183, w_017_522, w_023_047);
  nand2 I028_184(w_028_184, w_004_307, w_002_318);
  nand2 I028_185(w_028_185, w_004_450, w_014_210);
  not1 I028_186(w_028_186, w_009_407);
  or2  I028_187(w_028_187, w_025_124, w_003_051);
  or2  I028_190(w_028_190, w_021_191, w_024_430);
  not1 I028_191(w_028_191, w_010_300);
  or2  I028_196(w_028_196, w_011_262, w_014_069);
  and2 I028_197(w_028_197, w_005_084, w_014_054);
  not1 I028_198(w_028_198, w_024_119);
  or2  I028_200(w_028_200, w_006_028, w_006_079);
  or2  I028_201(w_028_201, w_021_119, w_002_466);
  not1 I028_202(w_028_202, w_020_527);
  and2 I028_203(w_028_203, w_003_001, w_002_256);
  not1 I028_204(w_028_204, w_019_011);
  and2 I028_205(w_028_205, w_004_305, w_008_467);
  not1 I028_206(w_028_206, w_012_041);
  and2 I028_208(w_028_208, w_025_110, w_003_051);
  and2 I028_209(w_028_209, w_005_228, w_019_010);
  and2 I028_215(w_028_215, w_022_270, w_010_361);
  or2  I028_216(w_028_216, w_000_450, w_003_018);
  nand2 I028_222(w_028_222, w_016_001, w_013_527);
  or2  I028_224(w_028_224, w_002_413, w_011_039);
  not1 I028_226(w_028_226, w_024_151);
  and2 I028_228(w_028_228, w_027_157, w_023_173);
  and2 I028_231(w_028_231, w_027_012, w_006_091);
  not1 I028_232(w_028_232, w_001_022);
  and2 I028_234(w_028_234, w_007_018, w_019_005);
  nand2 I028_240(w_028_240, w_004_474, w_019_016);
  nand2 I028_244(w_028_244, w_000_758, w_003_071);
  or2  I028_245(w_028_245, w_021_249, w_008_721);
  or2  I028_248(w_028_248, w_021_123, w_006_224);
  or2  I028_251(w_028_251, w_022_268, w_001_031);
  nand2 I028_252(w_028_252, w_012_215, w_015_131);
  nand2 I028_254(w_028_254, w_019_019, w_018_030);
  not1 I028_255(w_028_255, w_001_011);
  nand2 I028_256(w_028_256, w_019_006, w_014_216);
  and2 I028_258(w_028_258, w_023_009, w_023_175);
  not1 I028_260(w_028_260, w_001_010);
  and2 I028_262(w_028_262, w_002_435, w_025_264);
  not1 I028_263(w_028_263, w_017_430);
  and2 I028_264(w_028_264, w_022_011, w_020_536);
  not1 I028_267(w_028_267, w_012_007);
  and2 I028_268(w_028_268, w_014_095, w_002_396);
  not1 I028_270(w_028_270, w_011_616);
  nand2 I028_274(w_028_274, w_010_625, w_023_194);
  and2 I028_275(w_028_275, w_009_361, w_000_080);
  not1 I028_277(w_028_277, w_006_095);
  or2  I028_279(w_028_279, w_002_073, w_018_004);
  or2  I028_283(w_028_283, w_025_127, w_025_271);
  nand2 I028_284(w_028_284, w_015_620, w_014_219);
  nand2 I028_287(w_028_287, w_014_125, w_020_129);
  not1 I028_296(w_028_296, w_019_013);
  nand2 I028_299(w_028_299, w_000_522, w_004_402);
  nand2 I028_300(w_028_300, w_011_611, w_016_006);
  not1 I028_301(w_028_301, w_020_399);
  or2  I028_302(w_028_302, w_001_033, w_025_182);
  not1 I028_304(w_028_304, w_011_090);
  not1 I028_310(w_028_310, w_023_070);
  or2  I028_313(w_028_313, w_020_280, w_014_279);
  not1 I028_317(w_028_317, w_020_116);
  and2 I028_321(w_028_321, w_015_023, w_016_007);
  not1 I028_324(w_028_324, w_003_017);
  not1 I028_325(w_028_325, w_015_006);
  nand2 I028_326(w_028_326, w_003_027, w_006_073);
  not1 I028_335(w_028_335, w_002_030);
  nand2 I028_336(w_028_336, w_023_101, w_003_006);
  or2  I028_340(w_028_340, w_023_081, w_006_096);
  or2  I028_345(w_028_345, w_007_310, w_024_254);
  not1 I028_350(w_028_350, w_027_086);
  and2 I028_354(w_028_354, w_018_017, w_004_350);
  not1 I028_361(w_028_361, w_000_523);
  not1 I028_362(w_028_362, w_019_010);
  and2 I028_366(w_028_366, w_027_121, w_021_247);
  nand2 I028_368(w_028_368, w_016_007, w_025_043);
  nand2 I028_374(w_028_374, w_012_068, w_016_003);
  not1 I028_376(w_028_376, w_008_573);
  not1 I028_380(w_028_380, w_002_604);
  not1 I028_390(w_028_390, w_005_178);
  or2  I028_392(w_028_392, w_003_016, w_001_008);
  and2 I028_393(w_028_393, w_009_591, w_008_200);
  or2  I028_397(w_028_397, w_004_045, w_019_011);
  and2 I028_400(w_028_400, w_022_059, w_004_349);
  or2  I028_402(w_028_402, w_009_403, w_014_124);
  and2 I028_405(w_028_405, w_013_042, w_009_113);
  or2  I028_408(w_028_408, w_004_428, w_006_108);
  nand2 I028_409(w_028_409, w_021_084, w_010_158);
  or2  I028_411(w_028_411, w_004_221, w_001_001);
  or2  I028_413(w_028_413, w_002_162, w_027_012);
  and2 I028_415(w_028_415, w_011_163, w_012_158);
  not1 I028_416(w_028_416, w_024_189);
  not1 I028_425(w_028_425, w_020_162);
  or2  I028_427(w_028_427, w_014_209, w_016_001);
  or2  I028_433(w_028_433, w_024_117, w_005_236);
  nand2 I028_436(w_028_436, w_010_061, w_026_701);
  nand2 I028_437(w_028_437, w_023_165, w_002_204);
  and2 I028_438(w_028_438, w_004_225, w_016_004);
  not1 I028_440(w_028_440, w_015_652);
  and2 I028_441(w_028_441, w_014_081, w_015_124);
  nand2 I028_446(w_028_446, w_020_248, w_018_039);
  not1 I028_449(w_028_449, w_010_675);
  and2 I028_456(w_028_456, w_015_007, w_016_008);
  and2 I028_458(w_028_458, w_013_466, w_011_050);
  not1 I028_462(w_028_462, w_006_222);
  not1 I028_463(w_028_463, w_005_287);
  not1 I028_464(w_028_464, w_018_039);
  and2 I028_465(w_028_465, w_009_422, w_000_759);
  or2  I028_470(w_028_470, w_020_277, w_023_179);
  and2 I028_473(w_028_473, w_026_074, w_005_128);
  nand2 I028_474(w_028_474, w_026_274, w_016_001);
  nand2 I028_475(w_028_475, w_013_468, w_022_226);
  or2  I028_479(w_028_479, w_003_078, w_009_481);
  or2  I028_483(w_028_483, w_008_661, w_021_127);
  or2  I028_488(w_028_488, w_012_080, w_000_437);
  and2 I028_489(w_028_489, w_025_184, w_013_125);
  not1 I028_490(w_028_490, w_018_029);
  nand2 I028_491(w_028_491, w_012_155, w_027_167);
  or2  I028_497(w_028_497, w_004_346, w_000_192);
  or2  I028_499(w_028_499, w_026_163, w_022_045);
  nand2 I028_503(w_028_503, w_014_080, w_016_001);
  and2 I028_505(w_028_505, w_023_217, w_022_088);
  and2 I028_512(w_028_512, w_017_218, w_012_066);
  and2 I028_517(w_028_517, w_008_239, w_011_592);
  nand2 I028_521(w_028_521, w_000_297, w_019_013);
  nand2 I028_522(w_028_522, w_022_042, w_000_337);
  and2 I028_523(w_028_523, w_017_549, w_008_117);
  and2 I028_526(w_028_526, w_015_057, w_018_021);
  nand2 I028_527(w_028_527, w_010_209, w_008_729);
  or2  I028_528(w_028_528, w_023_076, w_009_121);
  or2  I028_536(w_028_536, w_017_235, w_003_009);
  nand2 I028_541(w_028_541, w_011_158, w_018_019);
  not1 I028_542(w_028_542, w_020_603);
  or2  I028_543(w_028_543, w_007_193, w_004_015);
  and2 I028_547(w_028_547, w_000_679, w_007_135);
  and2 I028_550(w_028_550, w_006_128, w_027_110);
  or2  I028_551(w_028_551, w_000_024, w_013_437);
  nand2 I028_554(w_028_554, w_020_125, w_020_074);
  or2  I028_559(w_028_559, w_007_017, w_022_071);
  and2 I028_560(w_028_560, w_008_287, w_007_052);
  nand2 I028_564(w_028_564, w_010_039, w_023_216);
  and2 I028_565(w_028_565, w_015_093, w_015_065);
  not1 I028_567(w_028_567, w_010_386);
  not1 I028_569(w_028_569, w_009_081);
  and2 I028_574(w_028_574, w_027_150, w_008_402);
  or2  I028_575(w_028_575, w_018_024, w_016_002);
  nand2 I028_578(w_028_578, w_017_108, w_023_139);
  or2  I028_586(w_028_586, w_008_097, w_022_059);
  and2 I028_587(w_028_589, w_001_029, w_028_588);
  or2  I028_588(w_028_590, w_028_589, w_019_012);
  or2  I028_589(w_028_591, w_001_005, w_028_590);
  not1 I028_590(w_028_592, w_028_591);
  nand2 I028_591(w_028_593, w_001_012, w_028_592);
  nand2 I028_592(w_028_594, w_028_593, w_013_311);
  or2  I028_593(w_028_595, w_020_576, w_028_594);
  not1 I028_594(w_028_596, w_028_595);
  and2 I028_595(w_028_597, w_028_596, w_028_607);
  nand2 I028_596(w_028_588, w_018_015, w_028_597);
  not1 I028_597(w_028_602, w_028_601);
  nand2 I028_598(w_028_603, w_013_256, w_028_602);
  nand2 I028_599(w_028_604, w_028_603, w_015_116);
  and2 I028_600(w_028_605, w_027_136, w_028_604);
  not1 I028_601(w_028_601, w_028_597);
  and2 I028_602(w_028_607, w_019_003, w_028_605);
  or2  I029_000(w_029_000, w_022_313, w_024_342);
  not1 I029_001(w_029_001, w_002_587);
  or2  I029_002(w_029_002, w_002_620, w_027_171);
  not1 I029_003(w_029_003, w_005_190);
  nand2 I029_004(w_029_004, w_023_054, w_027_070);
  and2 I029_005(w_029_005, w_025_305, w_005_079);
  or2  I029_006(w_029_006, w_027_188, w_024_478);
  or2  I029_007(w_029_007, w_017_343, w_028_483);
  or2  I029_008(w_029_008, w_022_270, w_023_214);
  nand2 I029_009(w_029_009, w_014_189, w_001_022);
  or2  I029_010(w_029_010, w_026_420, w_017_609);
  or2  I029_011(w_029_011, w_023_110, w_006_097);
  and2 I029_012(w_029_012, w_012_278, w_014_218);
  and2 I029_013(w_029_013, w_018_000, w_009_075);
  nand2 I029_014(w_029_014, w_011_085, w_016_006);
  not1 I029_015(w_029_015, w_000_459);
  or2  I029_016(w_029_016, w_022_293, w_004_443);
  nand2 I029_017(w_029_017, w_021_054, w_000_403);
  not1 I029_018(w_029_018, w_027_001);
  nand2 I029_019(w_029_019, w_011_036, w_018_007);
  or2  I029_020(w_029_020, w_007_332, w_001_002);
  and2 I029_021(w_029_021, w_012_260, w_014_150);
  not1 I029_022(w_029_022, w_006_103);
  and2 I029_023(w_029_023, w_028_065, w_008_737);
  and2 I029_024(w_029_024, w_000_541, w_018_025);
  and2 I029_025(w_029_025, w_008_681, w_016_008);
  not1 I029_026(w_029_026, w_005_031);
  nand2 I029_027(w_029_027, w_004_172, w_021_106);
  not1 I029_028(w_029_028, w_025_023);
  and2 I029_029(w_029_029, w_028_231, w_001_034);
  and2 I029_031(w_029_031, w_011_031, w_021_179);
  nand2 I029_032(w_029_032, w_000_163, w_012_314);
  or2  I029_033(w_029_033, w_009_216, w_019_018);
  or2  I029_035(w_029_035, w_028_317, w_015_047);
  and2 I029_036(w_029_036, w_017_003, w_021_022);
  or2  I029_037(w_029_037, w_003_057, w_000_377);
  nand2 I029_038(w_029_038, w_021_108, w_011_607);
  or2  I029_039(w_029_039, w_023_037, w_008_135);
  not1 I029_041(w_029_041, w_007_257);
  nand2 I029_042(w_029_042, w_023_086, w_004_295);
  not1 I029_043(w_029_043, w_017_669);
  and2 I029_044(w_029_044, w_021_181, w_006_161);
  and2 I029_045(w_029_045, w_020_525, w_023_095);
  nand2 I029_046(w_029_046, w_018_024, w_013_576);
  or2  I029_047(w_029_047, w_004_006, w_017_138);
  and2 I029_048(w_029_048, w_025_086, w_025_006);
  and2 I029_049(w_029_049, w_021_060, w_011_082);
  nand2 I029_050(w_029_050, w_017_372, w_012_333);
  nand2 I029_051(w_029_051, w_003_075, w_001_007);
  nand2 I029_052(w_029_052, w_027_076, w_019_001);
  or2  I029_053(w_029_053, w_012_082, w_014_035);
  nand2 I029_054(w_029_054, w_015_373, w_017_366);
  and2 I029_055(w_029_055, w_012_281, w_013_049);
  not1 I029_056(w_029_056, w_019_008);
  not1 I029_057(w_029_057, w_023_116);
  or2  I029_058(w_029_058, w_019_003, w_004_072);
  nand2 I029_059(w_029_059, w_023_197, w_026_530);
  and2 I029_060(w_029_060, w_009_163, w_000_142);
  nand2 I029_061(w_029_061, w_015_068, w_026_684);
  and2 I029_062(w_029_062, w_009_516, w_008_474);
  nand2 I029_063(w_029_063, w_019_013, w_025_233);
  not1 I029_064(w_029_064, w_007_132);
  not1 I029_065(w_029_065, w_003_034);
  or2  I029_066(w_029_066, w_018_014, w_010_289);
  or2  I029_067(w_029_067, w_011_004, w_000_392);
  nand2 I029_068(w_029_068, w_007_460, w_026_098);
  and2 I029_069(w_029_069, w_027_166, w_018_037);
  or2  I029_070(w_029_070, w_009_303, w_003_075);
  not1 I029_071(w_029_071, w_002_002);
  and2 I029_072(w_029_072, w_026_268, w_001_026);
  or2  I029_073(w_029_073, w_011_079, w_009_531);
  nand2 I029_074(w_029_074, w_001_012, w_008_612);
  nand2 I029_075(w_029_075, w_006_204, w_009_438);
  and2 I029_076(w_029_076, w_020_035, w_014_015);
  nand2 I029_077(w_029_077, w_009_237, w_012_131);
  nand2 I029_078(w_029_078, w_020_006, w_013_043);
  nand2 I029_079(w_029_079, w_022_267, w_003_019);
  and2 I029_080(w_029_080, w_011_564, w_023_109);
  and2 I029_081(w_029_081, w_022_031, w_004_163);
  not1 I029_082(w_029_082, w_019_007);
  or2  I029_083(w_029_083, w_025_170, w_019_002);
  not1 I029_085(w_029_085, w_023_108);
  not1 I029_086(w_029_086, w_008_639);
  and2 I029_087(w_029_087, w_002_599, w_027_051);
  not1 I029_088(w_029_088, w_009_184);
  and2 I029_089(w_029_089, w_019_017, w_017_014);
  or2  I029_090(w_029_090, w_010_423, w_017_470);
  and2 I029_091(w_029_091, w_015_060, w_019_018);
  not1 I029_092(w_029_092, w_005_270);
  and2 I029_093(w_029_093, w_013_256, w_007_418);
  and2 I029_094(w_029_094, w_001_015, w_019_019);
  and2 I029_095(w_029_095, w_020_576, w_022_201);
  nand2 I029_096(w_029_096, w_002_567, w_006_014);
  nand2 I029_097(w_029_097, w_015_443, w_013_484);
  not1 I029_098(w_029_098, w_003_057);
  and2 I029_099(w_029_099, w_001_023, w_025_142);
  not1 I029_100(w_029_100, w_024_378);
  not1 I029_101(w_029_101, w_026_500);
  nand2 I029_102(w_029_102, w_009_505, w_005_091);
  not1 I029_103(w_029_103, w_008_594);
  or2  I029_104(w_029_104, w_006_042, w_004_172);
  and2 I029_105(w_029_105, w_026_191, w_010_496);
  and2 I029_106(w_029_106, w_003_076, w_004_466);
  and2 I029_107(w_029_107, w_010_408, w_023_095);
  not1 I029_108(w_029_108, w_020_232);
  or2  I029_109(w_029_109, w_021_187, w_014_040);
  nand2 I029_110(w_029_110, w_022_074, w_004_357);
  not1 I029_111(w_029_111, w_008_530);
  not1 I029_112(w_029_112, w_026_273);
  nand2 I029_113(w_029_113, w_009_103, w_001_008);
  not1 I029_114(w_029_114, w_003_033);
  nand2 I029_115(w_029_115, w_023_067, w_027_088);
  and2 I029_116(w_029_116, w_028_111, w_008_180);
  and2 I029_117(w_029_117, w_018_001, w_017_068);
  and2 I029_118(w_028_599, w_023_096, w_028_588);
  nand2 I030_004(w_030_004, w_009_604, w_000_577);
  not1 I030_006(w_030_006, w_000_688);
  not1 I030_007(w_030_007, w_029_020);
  and2 I030_008(w_030_008, w_002_022, w_004_046);
  nand2 I030_009(w_030_009, w_004_203, w_010_315);
  not1 I030_011(w_030_011, w_023_181);
  nand2 I030_012(w_030_012, w_007_180, w_010_484);
  nand2 I030_013(w_030_013, w_003_008, w_016_004);
  nand2 I030_015(w_030_015, w_016_005, w_012_302);
  not1 I030_016(w_030_016, w_008_408);
  and2 I030_017(w_030_017, w_028_599, w_010_067);
  or2  I030_020(w_030_020, w_012_321, w_018_038);
  not1 I030_021(w_030_021, w_006_129);
  and2 I030_022(w_030_022, w_013_158, w_007_461);
  not1 I030_024(w_030_024, w_020_064);
  not1 I030_031(w_030_031, w_026_593);
  and2 I030_033(w_030_033, w_011_152, w_006_024);
  not1 I030_035(w_030_035, w_001_028);
  and2 I030_036(w_030_036, w_001_028, w_020_296);
  nand2 I030_037(w_030_037, w_006_142, w_025_098);
  nand2 I030_040(w_030_040, w_008_434, w_010_413);
  and2 I030_041(w_030_041, w_021_137, w_025_219);
  not1 I030_044(w_030_044, w_027_055);
  nand2 I030_047(w_030_047, w_006_051, w_013_166);
  or2  I030_048(w_030_048, w_009_521, w_012_013);
  and2 I030_049(w_030_049, w_025_145, w_005_091);
  and2 I030_050(w_030_050, w_015_045, w_028_522);
  nand2 I030_051(w_030_051, w_009_136, w_006_072);
  and2 I030_052(w_030_052, w_029_080, w_029_018);
  and2 I030_053(w_030_053, w_002_694, w_011_468);
  and2 I030_055(w_030_055, w_010_655, w_002_167);
  not1 I030_056(w_030_056, w_026_364);
  nand2 I030_057(w_030_057, w_016_005, w_028_175);
  nand2 I030_061(w_030_061, w_019_016, w_011_641);
  nand2 I030_064(w_030_064, w_005_017, w_002_591);
  or2  I030_067(w_030_067, w_017_032, w_010_308);
  or2  I030_069(w_030_069, w_004_134, w_021_103);
  and2 I030_070(w_030_070, w_014_236, w_026_411);
  or2  I030_071(w_030_071, w_028_202, w_003_020);
  or2  I030_073(w_030_073, w_001_008, w_010_623);
  or2  I030_074(w_030_074, w_029_031, w_025_247);
  and2 I030_076(w_030_076, w_015_582, w_009_241);
  or2  I030_077(w_030_077, w_010_421, w_007_123);
  not1 I030_078(w_030_078, w_009_026);
  or2  I030_080(w_030_080, w_017_092, w_012_216);
  nand2 I030_083(w_030_083, w_003_016, w_024_386);
  or2  I030_086(w_030_086, w_019_017, w_010_468);
  and2 I030_088(w_030_088, w_011_148, w_018_036);
  and2 I030_089(w_030_089, w_011_056, w_018_026);
  not1 I030_090(w_030_090, w_009_133);
  or2  I030_091(w_030_091, w_029_013, w_026_657);
  not1 I030_097(w_030_097, w_002_042);
  not1 I030_099(w_030_099, w_011_269);
  nand2 I030_100(w_030_100, w_015_309, w_029_079);
  not1 I030_101(w_030_101, w_017_404);
  and2 I030_102(w_030_102, w_012_281, w_018_021);
  and2 I030_104(w_030_104, w_028_030, w_008_602);
  or2  I030_105(w_030_105, w_006_140, w_010_061);
  or2  I030_106(w_030_106, w_013_330, w_000_371);
  nand2 I030_107(w_030_107, w_022_238, w_022_269);
  not1 I030_108(w_030_108, w_020_067);
  and2 I030_112(w_030_112, w_006_058, w_008_257);
  or2  I030_113(w_030_113, w_013_139, w_028_147);
  not1 I030_117(w_030_117, w_028_122);
  nand2 I030_119(w_030_119, w_010_703, w_009_444);
  or2  I030_121(w_030_121, w_019_019, w_012_040);
  not1 I030_123(w_030_123, w_009_226);
  or2  I030_125(w_030_125, w_021_243, w_023_121);
  and2 I030_132(w_030_132, w_010_726, w_026_224);
  and2 I030_134(w_030_134, w_020_359, w_018_026);
  nand2 I030_136(w_030_136, w_008_616, w_005_095);
  and2 I030_137(w_030_137, w_008_255, w_006_153);
  not1 I030_138(w_030_138, w_023_139);
  nand2 I030_143(w_030_143, w_023_125, w_004_067);
  nand2 I030_144(w_030_144, w_013_091, w_029_081);
  or2  I030_145(w_030_145, w_022_155, w_012_074);
  not1 I030_146(w_030_146, w_015_516);
  not1 I030_148(w_030_148, w_005_112);
  not1 I030_149(w_030_149, w_013_136);
  or2  I030_151(w_030_151, w_021_116, w_018_013);
  nand2 I030_152(w_030_152, w_012_181, w_010_591);
  and2 I030_155(w_030_155, w_028_076, w_016_008);
  nand2 I030_157(w_030_157, w_005_078, w_026_198);
  or2  I030_159(w_030_159, w_002_150, w_022_353);
  nand2 I030_161(w_030_161, w_026_527, w_013_246);
  not1 I030_162(w_030_162, w_000_660);
  and2 I030_163(w_030_163, w_010_633, w_024_327);
  not1 I030_167(w_030_167, w_009_089);
  or2  I030_168(w_030_168, w_027_001, w_017_314);
  not1 I030_171(w_030_171, w_027_008);
  not1 I030_172(w_030_172, w_024_434);
  nand2 I030_174(w_030_174, w_021_153, w_028_258);
  and2 I030_177(w_030_177, w_013_081, w_014_062);
  and2 I030_178(w_030_178, w_012_070, w_019_002);
  and2 I030_179(w_030_179, w_022_321, w_003_073);
  nand2 I030_180(w_030_180, w_001_033, w_024_082);
  nand2 I030_183(w_030_183, w_011_094, w_007_025);
  nand2 I030_184(w_030_184, w_025_079, w_023_042);
  and2 I030_185(w_030_185, w_023_021, w_028_458);
  or2  I030_188(w_030_188, w_000_311, w_023_017);
  nand2 I030_191(w_030_191, w_007_271, w_018_037);
  nand2 I030_192(w_030_192, w_007_049, w_013_274);
  nand2 I030_194(w_030_194, w_007_386, w_022_130);
  and2 I030_196(w_030_196, w_003_062, w_018_019);
  not1 I030_198(w_030_198, w_019_001);
  or2  I030_199(w_030_199, w_027_027, w_022_351);
  and2 I030_200(w_030_200, w_001_024, w_024_207);
  not1 I030_201(w_030_201, w_023_071);
  and2 I030_202(w_030_202, w_023_015, w_002_261);
  and2 I030_203(w_030_203, w_005_037, w_004_097);
  and2 I030_204(w_030_204, w_017_015, w_009_009);
  and2 I030_205(w_030_205, w_029_027, w_011_508);
  and2 I030_207(w_030_207, w_008_686, w_004_091);
  nand2 I030_208(w_030_208, w_018_006, w_025_025);
  or2  I030_210(w_030_210, w_007_367, w_015_116);
  or2  I030_212(w_030_212, w_021_103, w_013_489);
  nand2 I030_213(w_030_213, w_028_036, w_023_130);
  not1 I030_214(w_030_214, w_027_177);
  or2  I030_215(w_030_215, w_008_628, w_022_253);
  and2 I030_219(w_030_219, w_000_611, w_001_016);
  and2 I030_220(w_030_220, w_010_190, w_024_056);
  nand2 I030_222(w_030_222, w_013_115, w_002_666);
  not1 I030_223(w_030_223, w_027_184);
  not1 I030_224(w_030_224, w_022_052);
  nand2 I030_225(w_030_225, w_002_711, w_002_518);
  nand2 I030_226(w_030_226, w_024_101, w_002_045);
  not1 I030_227(w_030_227, w_012_235);
  and2 I030_228(w_030_228, w_020_288, w_009_452);
  nand2 I030_229(w_030_229, w_016_006, w_005_173);
  and2 I030_231(w_030_231, w_019_011, w_011_511);
  not1 I030_235(w_030_235, w_014_143);
  and2 I030_236(w_030_236, w_011_133, w_018_008);
  or2  I030_239(w_030_239, w_018_026, w_022_024);
  not1 I030_240(w_030_240, w_002_646);
  nand2 I030_241(w_030_241, w_010_569, w_025_125);
  nand2 I030_242(w_030_242, w_001_001, w_007_121);
  and2 I030_243(w_030_243, w_017_613, w_019_005);
  or2  I030_244(w_030_244, w_006_175, w_022_145);
  or2  I030_247(w_030_247, w_026_439, w_019_002);
  not1 I030_248(w_030_248, w_000_495);
  or2  I030_249(w_030_249, w_000_650, w_013_237);
  and2 I030_250(w_030_250, w_002_383, w_027_158);
  and2 I030_251(w_030_251, w_011_033, w_010_106);
  nand2 I030_252(w_030_252, w_023_091, w_012_338);
  nand2 I030_257(w_030_257, w_012_274, w_019_010);
  and2 I030_258(w_030_258, w_026_305, w_003_015);
  nand2 I030_259(w_030_259, w_028_427, w_002_319);
  and2 I030_261(w_030_261, w_009_551, w_008_023);
  nand2 I030_262(w_030_262, w_020_475, w_014_052);
  not1 I030_263(w_030_263, w_027_051);
  and2 I030_264(w_030_264, w_008_103, w_004_064);
  or2  I030_265(w_030_265, w_029_106, w_006_058);
  nand2 I030_267(w_030_267, w_020_037, w_006_191);
  and2 I030_268(w_030_268, w_014_180, w_002_486);
  nand2 I030_269(w_030_269, w_008_333, w_025_149);
  and2 I030_270(w_030_270, w_027_040, w_009_553);
  and2 I030_273(w_030_273, w_005_058, w_013_067);
  or2  I030_274(w_030_274, w_014_176, w_012_298);
  not1 I030_275(w_030_275, w_029_116);
  nand2 I030_276(w_030_276, w_025_083, w_023_090);
  nand2 I030_278(w_030_278, w_005_223, w_008_136);
  not1 I030_279(w_030_279, w_008_258);
  not1 I030_280(w_030_280, w_008_142);
  not1 I030_284(w_030_284, w_023_034);
  or2  I030_287(w_030_287, w_005_184, w_010_539);
  and2 I030_288(w_030_288, w_014_252, w_012_243);
  nand2 I030_290(w_030_290, w_013_176, w_004_226);
  and2 I030_291(w_030_291, w_027_011, w_015_092);
  nand2 I030_292(w_030_292, w_010_553, w_011_116);
  not1 I030_293(w_030_293, w_019_017);
  nand2 I030_295(w_030_295, w_000_397, w_004_365);
  nand2 I030_296(w_030_296, w_026_093, w_020_131);
  not1 I030_298(w_030_298, w_014_126);
  not1 I030_300(w_030_300, w_001_028);
  nand2 I030_301(w_030_301, w_022_148, w_023_120);
  and2 I030_302(w_030_302, w_000_270, w_002_444);
  or2  I030_305(w_030_305, w_019_009, w_027_070);
  and2 I030_307(w_030_307, w_014_155, w_005_116);
  and2 I030_308(w_030_308, w_020_442, w_017_433);
  and2 I030_309(w_030_309, w_011_077, w_005_311);
  not1 I030_311(w_030_311, w_028_226);
  or2  I030_312(w_030_312, w_018_009, w_026_018);
  nand2 I030_313(w_030_313, w_017_016, w_019_010);
  not1 I030_315(w_030_315, w_021_180);
  nand2 I030_316(w_030_316, w_003_014, w_014_126);
  and2 I030_317(w_030_317, w_028_497, w_015_548);
  nand2 I030_318(w_030_318, w_005_136, w_014_153);
  and2 I030_319(w_030_319, w_010_097, w_006_040);
  or2  I030_320(w_030_320, w_017_283, w_017_294);
  nand2 I030_324(w_030_324, w_023_052, w_029_039);
  and2 I030_325(w_030_325, w_020_300, w_003_018);
  nand2 I030_326(w_030_326, w_018_020, w_026_287);
  nand2 I030_327(w_030_327, w_001_028, w_012_103);
  and2 I030_328(w_030_328, w_027_143, w_018_011);
  and2 I030_330(w_030_330, w_006_042, w_005_175);
  not1 I030_331(w_030_331, w_021_167);
  not1 I030_332(w_030_332, w_024_155);
  and2 I030_337(w_030_337, w_005_271, w_009_172);
  or2  I030_338(w_030_338, w_000_090, w_003_004);
  or2  I030_339(w_030_339, w_027_169, w_012_089);
  and2 I030_340(w_030_340, w_017_034, w_023_098);
  nand2 I030_341(w_030_341, w_017_162, w_007_060);
  nand2 I030_345(w_030_345, w_019_005, w_007_021);
  or2  I030_346(w_030_346, w_001_013, w_010_756);
  and2 I030_348(w_030_348, w_017_093, w_014_167);
  nand2 I030_349(w_030_349, w_005_140, w_008_417);
  not1 I030_350(w_030_350, w_027_086);
  or2  I030_352(w_030_352, w_018_034, w_015_071);
  and2 I030_353(w_030_353, w_017_257, w_014_245);
  or2  I030_354(w_030_354, w_023_062, w_009_073);
  or2  I030_355(w_030_355, w_015_070, w_004_170);
  and2 I030_358(w_030_358, w_017_176, w_023_073);
  and2 I030_359(w_030_359, w_008_676, w_016_002);
  or2  I030_360(w_030_360, w_000_257, w_028_376);
  or2  I030_364(w_030_364, w_014_258, w_003_021);
  nand2 I030_365(w_030_365, w_018_028, w_025_147);
  nand2 I030_367(w_030_367, w_003_047, w_010_119);
  and2 I030_369(w_030_369, w_016_001, w_023_145);
  and2 I030_370(w_030_370, w_001_022, w_009_435);
  and2 I030_372(w_030_372, w_005_000, w_026_346);
  not1 I030_374(w_030_374, w_010_113);
  and2 I030_375(w_030_375, w_011_064, w_024_247);
  not1 I030_377(w_030_377, w_013_520);
  and2 I030_378(w_030_378, w_020_034, w_012_049);
  not1 I030_379(w_030_379, w_005_249);
  not1 I030_382(w_030_382, w_026_400);
  not1 I030_385(w_030_385, w_003_037);
  not1 I030_391(w_030_391, w_018_027);
  and2 I030_392(w_030_392, w_013_002, w_003_072);
  and2 I030_393(w_030_393, w_009_045, w_021_027);
  or2  I030_396(w_030_396, w_018_027, w_009_464);
  and2 I030_399(w_030_399, w_029_012, w_012_070);
  nand2 I030_408(w_030_408, w_013_076, w_004_355);
  and2 I030_409(w_030_409, w_025_249, w_017_464);
  or2  I030_410(w_030_410, w_005_048, w_024_172);
  not1 I030_411(w_030_411, w_018_018);
  nand2 I030_413(w_030_413, w_026_074, w_013_515);
  not1 I030_414(w_030_414, w_011_130);
  or2  I030_417(w_030_417, w_017_095, w_018_022);
  nand2 I030_419(w_030_419, w_027_159, w_018_003);
  not1 I031_001(w_031_001, w_020_012);
  nand2 I031_002(w_031_002, w_027_092, w_018_006);
  or2  I031_008(w_031_008, w_029_113, w_001_024);
  not1 I031_009(w_031_009, w_019_018);
  nand2 I031_011(w_031_011, w_002_648, w_013_171);
  or2  I031_012(w_031_012, w_006_108, w_000_207);
  nand2 I031_014(w_031_014, w_015_092, w_005_052);
  not1 I031_015(w_031_015, w_006_008);
  and2 I031_016(w_031_016, w_026_130, w_029_095);
  nand2 I031_017(w_031_017, w_016_005, w_019_001);
  or2  I031_020(w_031_020, w_014_129, w_009_335);
  not1 I031_021(w_031_021, w_015_258);
  not1 I031_026(w_031_026, w_010_540);
  not1 I031_027(w_031_027, w_001_005);
  and2 I031_030(w_031_030, w_004_295, w_000_331);
  and2 I031_032(w_031_032, w_027_092, w_008_724);
  or2  I031_033(w_031_033, w_030_123, w_009_109);
  and2 I031_034(w_031_034, w_008_115, w_023_201);
  nand2 I031_040(w_031_040, w_024_260, w_003_062);
  nand2 I031_043(w_031_043, w_026_288, w_008_460);
  or2  I031_049(w_031_049, w_000_213, w_002_582);
  and2 I031_050(w_031_050, w_014_217, w_011_248);
  not1 I031_054(w_031_054, w_005_260);
  nand2 I031_055(w_031_055, w_003_079, w_026_163);
  nand2 I031_058(w_031_058, w_015_023, w_022_029);
  not1 I031_059(w_031_059, w_019_018);
  nand2 I031_065(w_031_065, w_009_527, w_013_296);
  not1 I031_066(w_031_066, w_017_390);
  or2  I031_068(w_031_068, w_028_119, w_015_393);
  not1 I031_069(w_031_069, w_026_291);
  nand2 I031_070(w_031_070, w_013_178, w_028_156);
  and2 I031_072(w_031_072, w_024_265, w_017_279);
  nand2 I031_074(w_031_074, w_029_009, w_011_027);
  nand2 I031_076(w_031_076, w_024_139, w_003_065);
  or2  I031_081(w_031_081, w_007_214, w_012_203);
  and2 I031_082(w_031_082, w_030_024, w_014_074);
  nand2 I031_083(w_031_083, w_016_003, w_018_009);
  or2  I031_086(w_031_086, w_004_283, w_016_006);
  or2  I031_088(w_031_088, w_006_005, w_029_008);
  or2  I031_090(w_031_090, w_015_249, w_010_457);
  and2 I031_092(w_031_092, w_018_037, w_019_004);
  and2 I031_093(w_031_093, w_004_224, w_004_397);
  not1 I031_095(w_031_095, w_001_013);
  and2 I031_097(w_031_097, w_011_021, w_025_223);
  nand2 I031_100(w_031_100, w_007_112, w_017_010);
  or2  I031_101(w_031_101, w_018_040, w_030_191);
  or2  I031_102(w_031_102, w_017_025, w_020_571);
  nand2 I031_103(w_031_103, w_009_398, w_030_226);
  and2 I031_105(w_031_105, w_009_422, w_023_059);
  or2  I031_107(w_031_107, w_004_067, w_010_074);
  and2 I031_111(w_031_111, w_001_022, w_030_369);
  and2 I031_112(w_031_112, w_028_400, w_002_023);
  nand2 I031_116(w_031_116, w_011_102, w_005_108);
  nand2 I031_118(w_031_118, w_002_489, w_021_230);
  and2 I031_119(w_031_119, w_003_028, w_030_249);
  or2  I031_120(w_031_120, w_019_020, w_009_308);
  or2  I031_121(w_031_121, w_004_462, w_013_243);
  not1 I031_122(w_031_122, w_027_072);
  and2 I031_124(w_031_124, w_025_306, w_011_290);
  and2 I031_125(w_031_125, w_001_018, w_029_027);
  or2  I031_126(w_031_126, w_026_491, w_020_015);
  not1 I031_127(w_031_127, w_029_019);
  nand2 I031_128(w_031_128, w_000_153, w_027_112);
  nand2 I031_129(w_031_129, w_021_007, w_000_180);
  not1 I031_130(w_031_130, w_016_006);
  nand2 I031_131(w_031_131, w_008_523, w_003_073);
  and2 I031_133(w_031_133, w_026_125, w_019_001);
  nand2 I031_134(w_031_134, w_016_000, w_005_141);
  or2  I031_136(w_031_136, w_019_004, w_019_013);
  and2 I031_138(w_031_138, w_025_191, w_015_155);
  nand2 I031_143(w_031_143, w_010_530, w_004_392);
  or2  I031_144(w_031_144, w_014_163, w_028_198);
  and2 I031_145(w_031_145, w_022_251, w_014_268);
  nand2 I031_147(w_031_147, w_025_059, w_016_006);
  nand2 I031_148(w_031_148, w_021_230, w_013_372);
  or2  I031_150(w_031_150, w_007_328, w_024_065);
  not1 I031_151(w_031_151, w_025_166);
  or2  I031_153(w_031_153, w_007_038, w_003_015);
  not1 I031_154(w_031_154, w_020_272);
  or2  I031_155(w_031_155, w_010_777, w_023_092);
  not1 I031_156(w_031_156, w_021_083);
  or2  I031_160(w_031_160, w_013_210, w_002_418);
  not1 I031_161(w_031_161, w_002_368);
  nand2 I031_162(w_031_162, w_009_378, w_002_374);
  or2  I031_163(w_031_163, w_025_201, w_002_080);
  and2 I031_165(w_031_165, w_028_171, w_008_157);
  not1 I031_168(w_031_168, w_004_454);
  and2 I031_171(w_031_171, w_025_080, w_000_212);
  nand2 I031_174(w_031_174, w_001_006, w_009_032);
  nand2 I031_175(w_031_175, w_016_008, w_021_060);
  or2  I031_176(w_031_176, w_005_094, w_004_164);
  nand2 I031_177(w_031_177, w_002_184, w_022_140);
  or2  I031_178(w_031_178, w_015_095, w_017_512);
  or2  I031_179(w_031_179, w_029_091, w_020_543);
  nand2 I031_182(w_031_182, w_014_290, w_026_404);
  nand2 I031_186(w_031_186, w_027_063, w_026_632);
  or2  I031_188(w_031_188, w_026_548, w_030_259);
  not1 I031_193(w_031_193, w_021_072);
  not1 I031_195(w_031_195, w_008_449);
  or2  I031_202(w_031_202, w_014_004, w_016_004);
  nand2 I031_204(w_031_204, w_013_092, w_006_025);
  not1 I031_205(w_031_205, w_001_003);
  not1 I031_206(w_031_206, w_029_062);
  and2 I031_213(w_031_213, w_012_191, w_027_187);
  not1 I031_214(w_031_214, w_015_080);
  not1 I031_218(w_031_218, w_002_214);
  nand2 I031_223(w_031_223, w_009_074, w_001_026);
  not1 I031_231(w_031_231, w_002_033);
  nand2 I031_234(w_031_234, w_021_184, w_021_137);
  or2  I031_235(w_031_235, w_005_087, w_007_118);
  or2  I031_236(w_031_236, w_012_121, w_028_181);
  and2 I031_239(w_031_239, w_027_033, w_018_026);
  not1 I031_251(w_031_251, w_001_018);
  not1 I031_253(w_031_253, w_007_213);
  not1 I031_256(w_031_256, w_028_084);
  nand2 I031_259(w_031_259, w_009_611, w_001_021);
  or2  I031_260(w_031_260, w_006_247, w_025_126);
  not1 I031_265(w_031_265, w_002_195);
  and2 I031_268(w_031_268, w_005_136, w_023_079);
  and2 I031_271(w_031_271, w_002_696, w_006_168);
  and2 I031_272(w_031_272, w_004_081, w_001_014);
  not1 I031_273(w_031_273, w_027_122);
  not1 I031_276(w_031_276, w_012_034);
  nand2 I031_277(w_031_277, w_029_066, w_014_215);
  and2 I031_281(w_031_281, w_021_017, w_027_198);
  and2 I031_287(w_031_287, w_002_591, w_025_303);
  or2  I031_290(w_031_290, w_013_260, w_002_625);
  or2  I031_295(w_031_295, w_007_129, w_020_334);
  and2 I031_297(w_031_297, w_026_140, w_011_477);
  nand2 I031_302(w_031_302, w_001_015, w_001_006);
  or2  I031_308(w_031_308, w_021_180, w_010_612);
  and2 I031_309(w_031_309, w_018_001, w_001_014);
  nand2 I031_315(w_031_315, w_015_288, w_023_008);
  or2  I031_319(w_031_319, w_014_241, w_012_217);
  or2  I031_330(w_031_330, w_005_096, w_021_192);
  and2 I031_336(w_031_336, w_017_072, w_020_031);
  not1 I031_340(w_031_340, w_025_143);
  and2 I031_343(w_031_343, w_014_192, w_004_470);
  and2 I031_346(w_031_346, w_000_739, w_005_085);
  nand2 I031_356(w_031_356, w_001_010, w_019_007);
  nand2 I031_362(w_031_362, w_022_188, w_030_163);
  or2  I031_366(w_031_366, w_005_141, w_012_053);
  or2  I031_367(w_031_367, w_004_449, w_018_029);
  and2 I031_370(w_031_370, w_017_379, w_015_283);
  or2  I031_375(w_031_375, w_015_408, w_015_117);
  not1 I031_377(w_031_377, w_019_004);
  not1 I031_380(w_031_380, w_011_439);
  and2 I031_382(w_031_382, w_015_556, w_012_090);
  not1 I031_386(w_031_386, w_030_007);
  nand2 I031_387(w_031_387, w_001_015, w_017_376);
  and2 I031_389(w_031_389, w_024_107, w_021_265);
  nand2 I031_390(w_031_390, w_009_396, w_003_004);
  and2 I031_392(w_031_392, w_017_154, w_001_021);
  not1 I031_410(w_031_410, w_011_333);
  not1 I031_413(w_031_413, w_023_083);
  or2  I031_415(w_031_415, w_029_112, w_030_179);
  and2 I031_417(w_031_417, w_022_352, w_011_312);
  or2  I031_419(w_031_419, w_009_253, w_017_349);
  nand2 I031_420(w_031_420, w_009_068, w_001_015);
  and2 I031_422(w_031_422, w_030_227, w_024_222);
  nand2 I031_423(w_031_423, w_024_200, w_025_073);
  nand2 I031_425(w_031_425, w_001_021, w_002_072);
  and2 I031_434(w_031_434, w_004_088, w_011_135);
  nand2 I031_437(w_031_437, w_006_168, w_026_229);
  nand2 I031_439(w_031_439, w_014_009, w_013_296);
  and2 I031_440(w_031_440, w_028_397, w_020_033);
  nand2 I031_442(w_031_442, w_006_179, w_021_043);
  nand2 I031_444(w_031_444, w_016_004, w_017_047);
  nand2 I031_445(w_031_445, w_009_330, w_020_000);
  not1 I031_446(w_031_446, w_007_312);
  not1 I031_453(w_031_453, w_022_061);
  nand2 I031_456(w_031_456, w_009_093, w_026_172);
  not1 I031_457(w_031_457, w_021_237);
  and2 I031_460(w_031_460, w_017_178, w_006_117);
  nand2 I031_462(w_031_462, w_020_008, w_012_006);
  nand2 I031_463(w_031_463, w_019_003, w_003_036);
  and2 I031_465(w_031_465, w_020_005, w_027_089);
  or2  I031_466(w_031_466, w_011_098, w_013_121);
  not1 I031_467(w_031_467, w_002_221);
  or2  I031_469(w_031_469, w_006_113, w_023_150);
  and2 I031_470(w_031_470, w_011_201, w_006_226);
  and2 I031_471(w_031_471, w_029_000, w_022_144);
  not1 I031_472(w_031_472, w_011_111);
  nand2 I031_476(w_031_476, w_016_006, w_021_209);
  not1 I031_482(w_031_482, w_016_004);
  and2 I031_483(w_031_483, w_016_003, w_008_471);
  nand2 I031_487(w_031_487, w_011_295, w_028_187);
  or2  I031_488(w_031_488, w_018_012, w_020_122);
  nand2 I031_489(w_031_489, w_012_083, w_003_002);
  not1 I031_490(w_031_490, w_009_024);
  nand2 I031_494(w_031_494, w_024_181, w_030_037);
  nand2 I031_495(w_031_495, w_017_159, w_013_385);
  or2  I031_497(w_031_497, w_026_643, w_010_743);
  not1 I031_498(w_031_498, w_022_043);
  nand2 I031_499(w_031_499, w_030_358, w_015_445);
  and2 I031_501(w_031_501, w_012_059, w_010_408);
  or2  I031_508(w_031_508, w_030_337, w_007_285);
  or2  I031_509(w_031_509, w_012_095, w_015_443);
  nand2 I031_511(w_031_511, w_029_102, w_024_036);
  not1 I031_514(w_031_514, w_008_262);
  or2  I031_518(w_031_518, w_001_013, w_030_410);
  and2 I031_520(w_031_520, w_021_092, w_030_250);
  or2  I031_528(w_031_528, w_019_012, w_009_350);
  not1 I031_531(w_031_531, w_020_511);
  not1 I031_539(w_031_539, w_006_058);
  and2 I031_540(w_031_540, w_013_575, w_021_045);
  or2  I031_541(w_031_541, w_004_149, w_027_077);
  not1 I031_543(w_031_543, w_000_649);
  nand2 I031_546(w_031_546, w_004_508, w_006_153);
  not1 I031_548(w_031_548, w_001_011);
  and2 I031_553(w_031_553, w_024_441, w_029_008);
  or2  I031_555(w_031_555, w_020_198, w_003_019);
  and2 I031_556(w_031_556, w_019_005, w_007_234);
  or2  I031_557(w_031_557, w_001_022, w_014_067);
  and2 I031_558(w_031_558, w_003_076, w_016_006);
  or2  I031_561(w_031_561, w_023_150, w_006_122);
  nand2 I031_566(w_031_566, w_021_128, w_000_046);
  not1 I031_570(w_031_570, w_002_496);
  or2  I031_571(w_031_571, w_017_412, w_019_011);
  nand2 I031_574(w_031_574, w_017_157, w_023_083);
  and2 I031_581(w_031_581, w_013_061, w_030_061);
  nand2 I031_582(w_031_582, w_007_284, w_025_161);
  or2  I031_588(w_031_588, w_023_024, w_024_477);
  or2  I031_590(w_031_590, w_015_366, w_007_190);
  nand2 I031_593(w_031_593, w_017_118, w_009_255);
  nand2 I031_595(w_031_595, w_024_230, w_001_023);
  or2  I031_596(w_031_596, w_018_011, w_023_183);
  nand2 I031_599(w_031_599, w_023_052, w_028_183);
  not1 I031_601(w_031_601, w_015_484);
  and2 I031_602(w_031_602, w_015_577, w_013_097);
  or2  I031_604(w_031_604, w_012_254, w_020_043);
  not1 I031_605(w_031_605, w_003_059);
  and2 I031_609(w_031_611, w_031_610, w_029_048);
  or2  I031_610(w_031_612, w_031_611, w_002_537);
  not1 I031_611(w_031_613, w_031_612);
  nand2 I031_612(w_031_614, w_031_613, w_020_425);
  not1 I031_613(w_031_615, w_031_614);
  and2 I031_614(w_031_616, w_031_615, w_031_631);
  not1 I031_615(w_031_610, w_031_616);
  and2 I031_616(w_031_621, w_013_431, w_031_620);
  or2  I031_617(w_031_622, w_025_072, w_031_621);
  or2  I031_618(w_031_623, w_024_513, w_031_622);
  and2 I031_619(w_031_624, w_005_031, w_031_623);
  nand2 I031_620(w_031_625, w_031_624, w_026_703);
  not1 I031_621(w_031_626, w_031_625);
  nand2 I031_622(w_031_627, w_031_626, w_018_038);
  or2  I031_623(w_031_628, w_031_627, w_007_408);
  and2 I031_624(w_031_629, w_031_628, w_016_007);
  not1 I031_625(w_031_620, w_031_616);
  and2 I031_626(w_031_631, w_012_320, w_031_629);
  or2  I032_000(w_032_000, w_012_335, w_012_068);
  and2 I032_011(w_032_011, w_007_438, w_025_009);
  or2  I032_013(w_032_013, w_001_031, w_020_340);
  not1 I032_019(w_032_019, w_009_149);
  nand2 I032_021(w_032_021, w_004_388, w_019_003);
  and2 I032_022(w_032_022, w_010_633, w_002_083);
  or2  I032_025(w_032_025, w_000_275, w_027_138);
  and2 I032_028(w_032_028, w_027_197, w_028_101);
  and2 I032_030(w_032_030, w_007_295, w_006_167);
  not1 I032_031(w_032_031, w_031_143);
  and2 I032_033(w_032_033, w_001_007, w_016_004);
  and2 I032_037(w_032_037, w_018_002, w_014_106);
  and2 I032_039(w_032_039, w_015_059, w_024_081);
  not1 I032_041(w_032_041, w_029_037);
  not1 I032_042(w_032_042, w_015_087);
  not1 I032_043(w_032_043, w_020_515);
  and2 I032_044(w_032_044, w_005_135, w_026_039);
  or2  I032_045(w_032_045, w_013_509, w_013_190);
  or2  I032_046(w_032_046, w_007_223, w_013_000);
  and2 I032_049(w_032_049, w_029_085, w_027_120);
  or2  I032_051(w_032_051, w_029_060, w_010_459);
  or2  I032_052(w_032_052, w_024_433, w_015_511);
  and2 I032_053(w_032_053, w_028_296, w_008_026);
  and2 I032_057(w_032_057, w_007_345, w_025_164);
  or2  I032_060(w_032_060, w_010_579, w_025_016);
  nand2 I032_064(w_032_064, w_022_100, w_009_058);
  and2 I032_065(w_032_065, w_009_629, w_021_023);
  and2 I032_066(w_032_066, w_006_168, w_019_001);
  nand2 I032_067(w_032_067, w_010_603, w_022_332);
  and2 I032_068(w_032_068, w_002_597, w_023_105);
  and2 I032_072(w_032_072, w_005_165, w_030_280);
  and2 I032_073(w_032_073, w_005_069, w_000_092);
  or2  I032_074(w_032_074, w_020_030, w_031_235);
  not1 I032_076(w_032_076, w_011_555);
  nand2 I032_077(w_032_077, w_029_002, w_012_281);
  nand2 I032_078(w_032_078, w_021_267, w_003_062);
  nand2 I032_083(w_032_083, w_013_041, w_019_010);
  not1 I032_084(w_032_084, w_002_526);
  or2  I032_085(w_032_085, w_005_035, w_028_302);
  and2 I032_086(w_032_086, w_021_041, w_020_084);
  or2  I032_088(w_032_088, w_013_148, w_024_525);
  and2 I032_089(w_032_089, w_014_167, w_023_071);
  not1 I032_090(w_032_090, w_010_468);
  and2 I032_091(w_032_091, w_012_194, w_005_147);
  nand2 I032_092(w_032_092, w_001_010, w_028_140);
  and2 I032_095(w_032_095, w_015_253, w_028_060);
  nand2 I032_097(w_032_097, w_018_006, w_028_350);
  or2  I032_098(w_032_098, w_001_003, w_001_029);
  nand2 I032_099(w_032_099, w_029_002, w_030_194);
  or2  I032_102(w_032_102, w_031_076, w_002_231);
  not1 I032_103(w_032_103, w_026_442);
  and2 I032_105(w_032_105, w_012_346, w_024_133);
  and2 I032_106(w_032_106, w_022_086, w_026_693);
  nand2 I032_108(w_032_108, w_002_608, w_020_545);
  and2 I032_109(w_032_109, w_023_123, w_030_273);
  nand2 I032_110(w_032_110, w_012_167, w_027_023);
  nand2 I032_114(w_032_114, w_002_638, w_028_001);
  not1 I032_115(w_032_115, w_031_161);
  not1 I032_116(w_032_116, w_000_397);
  nand2 I032_118(w_032_118, w_009_050, w_014_022);
  not1 I032_120(w_032_120, w_026_010);
  not1 I032_121(w_032_121, w_001_024);
  and2 I032_122(w_032_122, w_000_548, w_025_113);
  nand2 I032_123(w_032_123, w_026_192, w_003_031);
  not1 I032_124(w_032_124, w_013_114);
  nand2 I032_129(w_032_129, w_028_087, w_022_214);
  or2  I032_132(w_032_132, w_018_000, w_015_604);
  or2  I032_133(w_032_133, w_004_036, w_030_009);
  nand2 I032_134(w_032_134, w_010_165, w_026_055);
  or2  I032_136(w_032_136, w_003_000, w_004_221);
  not1 I032_137(w_032_137, w_014_195);
  not1 I032_138(w_032_138, w_012_035);
  and2 I032_143(w_032_143, w_018_031, w_025_165);
  or2  I032_144(w_032_144, w_007_178, w_031_178);
  not1 I032_148(w_032_148, w_005_037);
  nand2 I032_149(w_032_149, w_014_013, w_010_577);
  or2  I032_150(w_032_150, w_028_340, w_026_555);
  not1 I032_151(w_032_151, w_001_026);
  or2  I032_152(w_032_152, w_020_403, w_013_367);
  not1 I032_153(w_032_153, w_015_468);
  or2  I032_154(w_032_154, w_008_556, w_005_221);
  nand2 I032_158(w_032_158, w_003_068, w_009_288);
  nand2 I032_160(w_032_160, w_013_386, w_006_100);
  not1 I032_163(w_032_163, w_008_648);
  not1 I032_165(w_032_165, w_016_004);
  nand2 I032_167(w_032_167, w_030_171, w_016_000);
  and2 I032_168(w_032_168, w_017_065, w_010_351);
  or2  I032_169(w_032_169, w_020_155, w_003_020);
  and2 I032_172(w_032_172, w_029_100, w_013_025);
  or2  I032_173(w_032_173, w_002_063, w_015_513);
  not1 I032_174(w_032_174, w_013_311);
  not1 I032_175(w_032_175, w_014_211);
  or2  I032_177(w_032_177, w_006_090, w_005_298);
  nand2 I032_178(w_032_178, w_012_052, w_031_514);
  nand2 I032_180(w_032_180, w_031_437, w_019_016);
  nand2 I032_183(w_032_183, w_015_497, w_024_182);
  and2 I032_184(w_032_184, w_029_115, w_000_202);
  not1 I032_185(w_032_185, w_031_268);
  not1 I032_186(w_032_186, w_028_554);
  nand2 I032_187(w_032_187, w_018_044, w_030_391);
  nand2 I032_189(w_032_189, w_015_607, w_019_013);
  not1 I032_191(w_032_191, w_025_038);
  and2 I032_192(w_032_192, w_024_130, w_006_112);
  or2  I032_193(w_032_193, w_018_017, w_001_034);
  and2 I032_194(w_032_194, w_019_017, w_011_474);
  not1 I032_195(w_032_195, w_009_472);
  nand2 I032_197(w_032_197, w_007_453, w_022_266);
  not1 I032_204(w_032_204, w_006_219);
  and2 I032_207(w_032_207, w_000_245, w_023_029);
  not1 I032_208(w_032_208, w_013_049);
  or2  I032_209(w_032_209, w_013_239, w_011_523);
  and2 I032_210(w_032_210, w_024_004, w_029_105);
  not1 I032_211(w_032_211, w_003_046);
  or2  I032_213(w_032_213, w_031_419, w_002_257);
  and2 I032_219(w_032_219, w_020_019, w_005_009);
  or2  I032_221(w_032_221, w_025_093, w_004_265);
  not1 I032_225(w_032_225, w_016_001);
  not1 I032_226(w_032_226, w_021_190);
  or2  I032_228(w_032_228, w_001_007, w_006_222);
  or2  I032_229(w_032_229, w_013_125, w_006_115);
  or2  I032_232(w_032_232, w_028_126, w_025_092);
  nand2 I032_234(w_032_234, w_004_330, w_009_529);
  and2 I032_239(w_032_239, w_004_128, w_000_315);
  not1 I032_240(w_032_240, w_027_082);
  or2  I032_243(w_032_243, w_027_067, w_006_036);
  not1 I032_247(w_032_247, w_004_010);
  not1 I032_249(w_032_249, w_029_032);
  and2 I032_254(w_032_254, w_010_078, w_010_156);
  or2  I032_257(w_032_257, w_026_048, w_001_017);
  nand2 I032_259(w_032_259, w_001_000, w_029_057);
  and2 I032_261(w_032_261, w_005_073, w_010_188);
  and2 I032_264(w_032_264, w_020_433, w_012_086);
  nand2 I032_269(w_032_269, w_009_343, w_026_507);
  nand2 I032_273(w_032_273, w_014_115, w_017_100);
  or2  I032_275(w_032_275, w_027_037, w_029_017);
  and2 I032_279(w_032_279, w_017_373, w_020_320);
  and2 I032_280(w_032_280, w_005_101, w_011_006);
  and2 I032_281(w_032_281, w_027_104, w_013_111);
  and2 I032_283(w_032_283, w_012_013, w_015_430);
  or2  I032_285(w_032_285, w_007_424, w_014_201);
  nand2 I032_287(w_032_287, w_020_381, w_022_129);
  or2  I032_290(w_032_290, w_007_222, w_013_002);
  and2 I032_293(w_032_293, w_013_229, w_009_099);
  not1 I032_294(w_032_294, w_029_079);
  not1 I032_295(w_032_295, w_029_076);
  nand2 I032_297(w_032_297, w_028_141, w_004_414);
  not1 I032_298(w_032_298, w_011_360);
  and2 I032_300(w_032_300, w_021_246, w_001_025);
  nand2 I032_307(w_032_307, w_029_103, w_024_213);
  not1 I032_309(w_032_309, w_026_064);
  or2  I032_310(w_032_310, w_009_081, w_020_476);
  or2  I032_312(w_032_312, w_031_102, w_001_019);
  and2 I032_313(w_032_313, w_031_179, w_028_380);
  not1 I032_321(w_032_321, w_027_153);
  or2  I032_322(w_032_322, w_026_705, w_030_346);
  or2  I032_325(w_032_325, w_000_383, w_017_662);
  or2  I032_328(w_032_328, w_020_609, w_006_239);
  or2  I032_330(w_032_330, w_017_132, w_027_073);
  and2 I032_331(w_032_331, w_025_154, w_026_088);
  or2  I032_342(w_032_342, w_012_237, w_005_025);
  or2  I032_345(w_032_345, w_027_101, w_020_420);
  nand2 I032_346(w_032_346, w_016_005, w_029_100);
  not1 I032_348(w_032_348, w_031_195);
  or2  I032_350(w_032_350, w_031_489, w_011_047);
  and2 I032_352(w_032_352, w_006_221, w_023_099);
  or2  I032_355(w_032_355, w_030_319, w_016_000);
  or2  I032_357(w_032_357, w_006_104, w_031_472);
  not1 I032_359(w_032_359, w_004_319);
  nand2 I032_360(w_032_360, w_006_224, w_004_228);
  not1 I032_363(w_032_363, w_029_029);
  nand2 I032_364(w_032_364, w_003_039, w_018_032);
  or2  I032_368(w_032_368, w_019_006, w_023_113);
  or2  I032_376(w_032_376, w_009_135, w_030_379);
  or2  I032_377(w_032_377, w_027_129, w_018_024);
  nand2 I032_379(w_032_379, w_013_207, w_014_028);
  nand2 I032_389(w_032_389, w_020_605, w_002_552);
  and2 I032_391(w_032_391, w_007_211, w_024_272);
  nand2 I032_395(w_032_395, w_021_164, w_013_211);
  and2 I032_398(w_032_398, w_020_389, w_025_013);
  nand2 I032_399(w_032_399, w_031_012, w_022_087);
  and2 I032_404(w_032_404, w_018_007, w_004_072);
  nand2 I032_409(w_032_409, w_004_245, w_003_072);
  nand2 I032_410(w_032_410, w_019_000, w_015_088);
  and2 I032_411(w_032_411, w_027_073, w_029_107);
  not1 I032_414(w_032_414, w_008_589);
  not1 I032_418(w_032_418, w_002_466);
  not1 I032_425(w_032_425, w_027_031);
  and2 I032_429(w_032_429, w_022_367, w_023_206);
  and2 I032_430(w_032_430, w_021_115, w_018_011);
  nand2 I032_433(w_032_433, w_004_214, w_001_033);
  and2 I032_434(w_032_434, w_017_367, w_003_010);
  and2 I032_437(w_032_437, w_003_073, w_031_499);
  not1 I032_438(w_032_438, w_026_343);
  not1 I032_442(w_032_442, w_029_097);
  not1 I032_443(w_032_443, w_018_004);
  and2 I032_444(w_032_444, w_026_051, w_012_056);
  or2  I032_445(w_032_445, w_031_422, w_003_022);
  not1 I032_446(w_032_446, w_020_564);
  not1 I032_448(w_032_448, w_021_077);
  and2 I032_449(w_032_449, w_016_006, w_018_029);
  nand2 I032_451(w_032_451, w_020_423, w_001_036);
  or2  I032_457(w_032_457, w_005_014, w_017_569);
  nand2 I032_462(w_032_462, w_004_383, w_004_202);
  nand2 I032_464(w_032_464, w_023_153, w_024_108);
  nand2 I032_465(w_032_465, w_008_753, w_031_511);
  nand2 I032_466(w_032_466, w_013_329, w_014_048);
  or2  I032_471(w_032_471, w_031_176, w_022_062);
  nand2 I032_477(w_032_477, w_002_075, w_024_189);
  and2 I032_478(w_032_478, w_014_031, w_013_151);
  nand2 I032_490(w_032_490, w_027_124, w_013_401);
  nand2 I032_491(w_032_491, w_024_082, w_019_013);
  not1 I032_493(w_032_493, w_013_181);
  not1 I032_496(w_032_496, w_026_068);
  not1 I032_497(w_032_497, w_020_551);
  or2  I032_499(w_032_499, w_013_329, w_018_034);
  and2 I032_502(w_032_502, w_014_054, w_026_044);
  and2 I032_504(w_032_504, w_022_231, w_024_478);
  and2 I032_507(w_032_507, w_020_329, w_024_060);
  nand2 I032_508(w_032_508, w_025_173, w_028_156);
  nand2 I032_509(w_032_509, w_022_378, w_001_035);
  nand2 I032_510(w_032_510, w_005_160, w_008_189);
  or2  I032_512(w_032_512, w_015_235, w_031_065);
  or2  I032_514(w_032_514, w_020_380, w_009_080);
  and2 I032_515(w_032_515, w_000_326, w_024_577);
  or2  I032_520(w_032_520, w_019_011, w_009_540);
  nand2 I032_521(w_032_521, w_013_188, w_010_197);
  or2  I032_524(w_032_524, w_027_053, w_029_024);
  and2 I032_525(w_032_525, w_010_597, w_030_033);
  or2  I032_526(w_032_526, w_011_352, w_008_405);
  nand2 I032_533(w_032_533, w_010_627, w_008_511);
  nand2 I032_537(w_032_537, w_029_080, w_027_159);
  or2  I032_540(w_032_540, w_015_258, w_021_093);
  and2 I032_541(w_032_541, w_029_043, w_013_572);
  and2 I032_545(w_032_545, w_014_188, w_031_469);
  or2  I032_546(w_032_546, w_004_325, w_020_025);
  or2  I032_552(w_032_552, w_004_223, w_018_009);
  nand2 I032_553(w_032_553, w_026_304, w_014_231);
  and2 I032_559(w_032_559, w_005_115, w_012_275);
  not1 I032_562(w_032_562, w_026_595);
  not1 I032_568(w_032_568, w_024_088);
  nand2 I032_569(w_032_569, w_027_185, w_014_206);
  and2 I032_570(w_032_570, w_017_286, w_019_000);
  not1 I032_574(w_032_574, w_021_047);
  not1 I032_575(w_032_575, w_019_015);
  or2  I032_579(w_032_579, w_029_069, w_031_518);
  or2  I032_583(w_032_583, w_010_460, w_019_010);
  nand2 I032_588(w_032_588, w_023_147, w_009_621);
  and2 I032_594(w_032_594, w_022_348, w_011_587);
  and2 I032_596(w_032_596, w_023_083, w_017_164);
  not1 I032_597(w_032_597, w_006_078);
  not1 I032_599(w_032_599, w_013_000);
  not1 I032_602(w_032_604, w_032_603);
  or2  I032_603(w_032_605, w_032_604, w_008_588);
  and2 I032_604(w_032_606, w_023_206, w_032_605);
  and2 I032_605(w_032_607, w_032_606, w_021_050);
  and2 I032_606(w_032_603, w_012_001, w_032_607);
  and2 I032_607(w_031_618, w_006_241, w_031_610);
  not1 I033_001(w_033_001, w_016_005);
  not1 I033_002(w_033_002, w_000_599);
  nand2 I033_008(w_033_008, w_005_257, w_028_040);
  nand2 I033_009(w_033_009, w_024_008, w_003_079);
  or2  I033_011(w_033_011, w_002_651, w_002_065);
  nand2 I033_012(w_033_012, w_030_163, w_025_028);
  or2  I033_014(w_033_014, w_012_263, w_019_019);
  not1 I033_015(w_033_015, w_032_376);
  nand2 I033_016(w_033_016, w_000_347, w_006_000);
  or2  I033_017(w_033_017, w_000_141, w_011_147);
  not1 I033_019(w_033_019, w_018_032);
  nand2 I033_021(w_033_021, w_008_312, w_007_149);
  or2  I033_022(w_033_022, w_011_356, w_010_454);
  nand2 I033_024(w_033_024, w_020_088, w_031_265);
  not1 I033_026(w_033_026, w_019_010);
  and2 I033_029(w_033_029, w_004_071, w_005_107);
  or2  I033_053(w_033_053, w_014_120, w_009_080);
  not1 I033_057(w_033_057, w_005_152);
  or2  I033_059(w_033_059, w_002_480, w_028_416);
  nand2 I033_061(w_033_061, w_015_299, w_020_403);
  nand2 I033_062(w_033_062, w_003_054, w_010_680);
  not1 I033_065(w_033_065, w_013_446);
  or2  I033_068(w_033_068, w_026_039, w_008_273);
  nand2 I033_076(w_033_076, w_001_007, w_026_008);
  or2  I033_082(w_033_082, w_005_245, w_022_194);
  or2  I033_084(w_033_084, w_008_414, w_000_405);
  and2 I033_085(w_033_085, w_004_326, w_029_004);
  or2  I033_086(w_033_086, w_001_016, w_020_425);
  not1 I033_087(w_033_087, w_021_226);
  not1 I033_091(w_033_091, w_008_189);
  nand2 I033_094(w_033_094, w_009_342, w_017_096);
  not1 I033_095(w_033_095, w_031_336);
  nand2 I033_100(w_033_100, w_030_408, w_023_054);
  and2 I033_109(w_033_109, w_010_043, w_014_237);
  not1 I033_111(w_033_111, w_009_006);
  and2 I033_114(w_033_114, w_018_040, w_026_317);
  or2  I033_116(w_033_116, w_021_059, w_025_010);
  not1 I033_119(w_033_119, w_006_001);
  nand2 I033_121(w_033_121, w_001_011, w_003_056);
  or2  I033_123(w_033_123, w_027_093, w_015_083);
  or2  I033_127(w_033_127, w_014_003, w_018_003);
  or2  I033_129(w_033_129, w_005_023, w_013_110);
  not1 I033_132(w_033_132, w_017_297);
  or2  I033_142(w_033_142, w_012_126, w_016_008);
  nand2 I033_143(w_033_143, w_028_560, w_011_371);
  not1 I033_148(w_033_148, w_022_322);
  nand2 I033_149(w_033_149, w_001_004, w_013_159);
  and2 I033_157(w_033_157, w_031_483, w_026_687);
  and2 I033_159(w_033_159, w_029_061, w_025_290);
  or2  I033_160(w_033_160, w_023_071, w_003_046);
  and2 I033_161(w_033_161, w_011_632, w_032_060);
  or2  I033_162(w_033_162, w_009_546, w_029_082);
  or2  I033_163(w_033_163, w_019_012, w_019_007);
  and2 I033_171(w_033_171, w_013_370, w_031_068);
  or2  I033_172(w_033_172, w_009_335, w_002_220);
  and2 I033_181(w_033_181, w_027_080, w_015_608);
  or2  I033_182(w_033_182, w_032_090, w_018_022);
  not1 I033_183(w_033_183, w_005_267);
  or2  I033_184(w_033_184, w_003_064, w_012_119);
  and2 I033_191(w_033_191, w_008_751, w_024_040);
  nand2 I033_194(w_033_194, w_003_019, w_019_003);
  not1 I033_197(w_033_197, w_021_099);
  or2  I033_200(w_033_200, w_020_306, w_007_014);
  or2  I033_201(w_033_201, w_009_288, w_025_211);
  nand2 I033_207(w_033_207, w_008_047, w_019_008);
  nand2 I033_208(w_033_208, w_009_143, w_017_174);
  nand2 I033_209(w_033_209, w_013_086, w_031_121);
  or2  I033_216(w_033_216, w_031_581, w_027_125);
  not1 I033_217(w_033_217, w_013_162);
  not1 I033_220(w_033_220, w_007_438);
  not1 I033_224(w_033_224, w_000_706);
  nand2 I033_231(w_033_231, w_007_292, w_020_032);
  not1 I033_235(w_033_235, w_030_300);
  or2  I033_236(w_033_236, w_004_190, w_016_003);
  and2 I033_238(w_033_238, w_015_215, w_012_033);
  or2  I033_241(w_033_241, w_006_009, w_012_262);
  nand2 I033_244(w_033_244, w_030_031, w_000_181);
  or2  I033_249(w_033_249, w_006_236, w_002_534);
  or2  I033_250(w_033_250, w_020_355, w_003_018);
  nand2 I033_251(w_033_251, w_000_014, w_008_031);
  not1 I033_253(w_033_253, w_002_247);
  nand2 I033_256(w_033_256, w_017_482, w_022_114);
  or2  I033_259(w_033_259, w_032_570, w_007_064);
  nand2 I033_263(w_033_263, w_014_019, w_014_168);
  not1 I033_269(w_033_269, w_031_582);
  not1 I033_272(w_033_272, w_017_116);
  nand2 I033_275(w_033_275, w_007_364, w_015_178);
  not1 I033_278(w_033_278, w_016_001);
  and2 I033_282(w_033_282, w_020_205, w_010_385);
  nand2 I033_289(w_033_289, w_008_145, w_015_232);
  and2 I033_291(w_033_291, w_006_235, w_013_321);
  nand2 I033_293(w_033_293, w_001_009, w_000_603);
  not1 I033_297(w_033_297, w_030_348);
  or2  I033_309(w_033_309, w_023_158, w_003_048);
  nand2 I033_310(w_033_310, w_008_037, w_026_042);
  nand2 I033_312(w_033_312, w_014_056, w_015_538);
  nand2 I033_313(w_033_313, w_031_162, w_032_537);
  and2 I033_318(w_033_318, w_010_589, w_001_001);
  nand2 I033_319(w_033_319, w_018_036, w_021_233);
  and2 I033_321(w_033_321, w_016_007, w_013_141);
  and2 I033_322(w_033_322, w_001_010, w_022_333);
  nand2 I033_323(w_033_323, w_002_305, w_016_004);
  not1 I033_328(w_033_328, w_028_184);
  or2  I033_329(w_033_329, w_017_267, w_008_215);
  and2 I033_330(w_033_330, w_022_383, w_031_032);
  not1 I033_331(w_033_331, w_028_025);
  nand2 I033_335(w_033_335, w_001_026, w_001_022);
  nand2 I033_336(w_033_336, w_011_357, w_019_000);
  or2  I033_339(w_033_339, w_010_016, w_026_216);
  and2 I033_340(w_033_340, w_011_635, w_002_623);
  and2 I033_341(w_033_341, w_024_461, w_009_274);
  and2 I033_354(w_033_354, w_002_162, w_032_103);
  and2 I033_355(w_033_355, w_028_559, w_019_016);
  nand2 I033_358(w_033_358, w_019_007, w_030_419);
  or2  I033_363(w_033_363, w_008_218, w_017_513);
  not1 I033_365(w_033_365, w_029_105);
  and2 I033_366(w_033_366, w_023_210, w_015_220);
  not1 I033_369(w_033_369, w_010_400);
  nand2 I033_372(w_033_372, w_004_013, w_016_008);
  or2  I033_377(w_033_377, w_015_449, w_031_498);
  nand2 I033_378(w_033_378, w_022_266, w_015_133);
  and2 I033_379(w_033_379, w_029_055, w_014_089);
  not1 I033_380(w_033_380, w_026_184);
  and2 I033_382(w_033_382, w_020_606, w_016_004);
  nand2 I033_391(w_033_391, w_000_458, w_029_052);
  not1 I033_392(w_033_392, w_017_626);
  not1 I033_396(w_033_396, w_017_373);
  and2 I033_404(w_033_404, w_012_041, w_029_046);
  nand2 I033_406(w_033_406, w_005_143, w_029_051);
  nand2 I033_407(w_033_407, w_009_050, w_031_389);
  nand2 I033_414(w_033_414, w_002_272, w_017_177);
  nand2 I033_419(w_033_419, w_016_008, w_016_007);
  not1 I033_426(w_033_426, w_006_098);
  and2 I033_427(w_033_427, w_032_355, w_008_713);
  nand2 I033_428(w_033_428, w_027_145, w_022_200);
  or2  I033_436(w_033_436, w_023_095, w_008_755);
  or2  I033_437(w_033_437, w_002_406, w_011_020);
  and2 I033_442(w_033_442, w_031_417, w_015_092);
  not1 I033_447(w_033_447, w_001_002);
  nand2 I033_449(w_033_449, w_019_019, w_028_512);
  and2 I033_451(w_033_451, w_011_465, w_005_044);
  nand2 I033_452(w_033_452, w_002_358, w_002_657);
  and2 I033_453(w_033_453, w_001_007, w_024_551);
  not1 I033_462(w_033_462, w_017_070);
  not1 I033_468(w_033_468, w_011_201);
  not1 I033_475(w_033_475, w_029_042);
  and2 I033_486(w_033_486, w_030_208, w_006_026);
  and2 I033_487(w_033_487, w_015_106, w_019_020);
  nand2 I033_488(w_033_488, w_031_163, w_015_113);
  or2  I033_492(w_033_492, w_010_593, w_009_194);
  and2 I033_493(w_033_493, w_015_393, w_003_067);
  and2 I033_494(w_033_494, w_011_471, w_018_043);
  not1 I033_505(w_033_505, w_026_447);
  nand2 I033_506(w_033_506, w_019_001, w_009_182);
  nand2 I033_509(w_033_509, w_012_205, w_029_067);
  and2 I033_510(w_033_510, w_031_618, w_006_184);
  nand2 I033_511(w_033_511, w_014_024, w_014_018);
  and2 I033_512(w_033_512, w_015_598, w_004_374);
  and2 I033_513(w_033_513, w_027_067, w_010_515);
  nand2 I033_515(w_033_515, w_024_172, w_017_603);
  and2 I033_516(w_033_516, w_011_342, w_020_577);
  and2 I033_517(w_033_517, w_026_566, w_023_150);
  and2 I033_522(w_033_522, w_024_559, w_004_091);
  nand2 I033_530(w_033_530, w_016_007, w_012_053);
  and2 I033_534(w_033_534, w_028_145, w_002_496);
  not1 I033_535(w_033_535, w_009_045);
  nand2 I033_537(w_033_537, w_005_050, w_016_003);
  nand2 I033_539(w_033_539, w_015_149, w_017_243);
  not1 I033_541(w_033_541, w_021_118);
  nand2 I033_545(w_033_545, w_005_017, w_018_023);
  or2  I033_546(w_033_546, w_000_268, w_004_445);
  or2  I033_551(w_033_551, w_018_026, w_006_191);
  not1 I033_555(w_033_555, w_002_616);
  not1 I033_557(w_033_557, w_022_177);
  nand2 I033_558(w_033_558, w_013_064, w_016_004);
  not1 I033_560(w_033_560, w_004_071);
  and2 I033_566(w_033_566, w_030_070, w_009_136);
  or2  I033_568(w_033_568, w_001_005, w_017_057);
  not1 I033_569(w_033_569, w_017_407);
  or2  I033_574(w_033_574, w_018_035, w_031_177);
  and2 I033_580(w_033_580, w_012_042, w_004_159);
  nand2 I033_583(w_033_583, w_012_063, w_022_170);
  not1 I033_587(w_033_587, w_018_014);
  or2  I033_590(w_033_590, w_017_193, w_018_029);
  not1 I033_604(w_033_604, w_022_017);
  not1 I033_605(w_033_605, w_027_006);
  nand2 I033_608(w_033_608, w_029_047, w_019_017);
  and2 I033_613(w_033_613, w_026_290, w_001_028);
  or2  I033_614(w_033_614, w_023_156, w_008_351);
  or2  I033_617(w_033_617, w_025_247, w_022_268);
  and2 I033_618(w_033_618, w_008_227, w_003_042);
  and2 I033_619(w_033_619, w_004_050, w_018_037);
  and2 I033_622(w_033_622, w_004_124, w_011_279);
  or2  I033_629(w_033_629, w_012_200, w_015_248);
  not1 I033_630(w_033_630, w_031_476);
  and2 I033_631(w_033_631, w_030_393, w_030_338);
  not1 I033_637(w_033_637, w_005_038);
  nand2 I033_638(w_033_638, w_002_566, w_005_273);
  and2 I033_639(w_033_639, w_031_574, w_013_522);
  and2 I033_646(w_033_646, w_013_353, w_003_076);
  nand2 I033_647(w_033_647, w_019_017, w_019_004);
  nand2 I033_653(w_033_653, w_022_149, w_018_019);
  nand2 I033_656(w_033_656, w_032_273, w_010_076);
  or2  I033_658(w_033_658, w_010_009, w_005_121);
  or2  I033_660(w_033_660, w_022_200, w_008_449);
  and2 I033_670(w_033_670, w_002_311, w_032_051);
  and2 I033_671(w_033_671, w_009_230, w_008_016);
  nand2 I033_675(w_033_675, w_032_446, w_013_011);
  nand2 I033_685(w_033_685, w_023_082, w_019_008);
  not1 I033_689(w_033_689, w_010_417);
  and2 I033_692(w_033_692, w_028_034, w_003_027);
  or2  I033_695(w_033_695, w_003_081, w_012_177);
  nand2 I033_698(w_033_698, w_012_293, w_010_328);
  or2  I033_703(w_033_703, w_017_234, w_026_000);
  not1 I033_705(w_033_705, w_013_016);
  and2 I033_710(w_033_710, w_024_051, w_010_499);
  or2  I033_711(w_033_711, w_011_187, w_019_019);
  or2  I033_715(w_033_715, w_010_415, w_019_009);
  nand2 I033_718(w_033_718, w_006_003, w_008_024);
  and2 I033_719(w_033_719, w_002_500, w_009_594);
  or2  I033_722(w_033_722, w_032_552, w_020_065);
  nand2 I033_724(w_033_724, w_031_501, w_018_024);
  and2 I033_725(w_033_725, w_011_017, w_027_184);
  not1 I033_726(w_033_726, w_022_315);
  not1 I033_727(w_033_727, w_000_564);
  nand2 I033_730(w_033_730, w_026_534, w_005_104);
  or2  I033_735(w_033_735, w_008_504, w_000_259);
  not1 I033_740(w_033_740, w_031_482);
  nand2 I033_745(w_033_745, w_005_164, w_007_042);
  not1 I033_748(w_033_748, w_016_003);
  or2  I033_751(w_033_751, w_003_039, w_007_029);
  not1 I033_753(w_033_753, w_002_711);
  not1 I033_756(w_033_756, w_004_269);
  nand2 I033_762(w_033_762, w_022_128, w_005_146);
  not1 I033_766(w_033_766, w_017_280);
  nand2 I033_769(w_033_769, w_017_562, w_031_081);
  not1 I033_770(w_033_770, w_028_436);
  not1 I033_771(w_033_771, w_020_445);
  not1 I033_775(w_033_775, w_020_490);
  nand2 I033_779(w_033_779, w_012_257, w_014_099);
  not1 I033_783(w_033_783, w_006_068);
  and2 I033_784(w_032_609, w_001_027, w_032_603);
  or2  I034_000(w_034_000, w_016_003, w_023_158);
  and2 I034_001(w_034_001, w_022_136, w_010_177);
  and2 I034_002(w_034_002, w_023_216, w_026_257);
  not1 I034_003(w_034_003, w_009_193);
  nand2 I034_004(w_034_004, w_030_088, w_004_035);
  nand2 I034_005(w_034_005, w_002_495, w_015_142);
  not1 I034_006(w_034_006, w_020_416);
  nand2 I034_007(w_034_007, w_003_081, w_024_557);
  or2  I034_008(w_034_008, w_012_304, w_025_113);
  nand2 I034_009(w_034_009, w_022_408, w_023_073);
  not1 I034_010(w_034_010, w_007_220);
  not1 I034_011(w_034_011, w_003_004);
  and2 I034_012(w_034_012, w_008_568, w_004_199);
  not1 I034_013(w_034_013, w_005_015);
  and2 I034_015(w_034_015, w_020_126, w_010_099);
  not1 I034_016(w_034_016, w_030_359);
  not1 I034_017(w_034_017, w_000_032);
  and2 I034_018(w_034_018, w_025_304, w_000_659);
  and2 I034_019(w_034_019, w_028_200, w_013_372);
  nand2 I034_020(w_034_020, w_004_182, w_000_714);
  nand2 I034_021(w_034_021, w_014_142, w_022_247);
  and2 I034_022(w_034_022, w_017_054, w_000_386);
  nand2 I034_023(w_034_023, w_031_297, w_006_177);
  not1 I034_024(w_034_024, w_014_004);
  nand2 I034_025(w_034_025, w_014_009, w_006_174);
  and2 I034_026(w_034_026, w_027_048, w_032_477);
  nand2 I034_027(w_034_027, w_006_238, w_002_092);
  and2 I034_028(w_034_028, w_033_339, w_006_166);
  or2  I034_029(w_034_029, w_014_016, w_024_499);
  and2 I034_030(w_034_030, w_004_167, w_004_264);
  nand2 I034_031(w_034_031, w_005_022, w_015_209);
  or2  I034_032(w_034_032, w_025_210, w_012_277);
  and2 I034_033(w_034_033, w_018_032, w_016_005);
  and2 I034_034(w_034_034, w_032_293, w_032_132);
  or2  I034_035(w_034_035, w_011_180, w_016_002);
  and2 I034_036(w_034_036, w_028_196, w_019_001);
  and2 I034_037(w_034_037, w_014_070, w_013_077);
  or2  I034_038(w_034_038, w_003_015, w_033_249);
  and2 I034_039(w_034_039, w_025_263, w_020_147);
  and2 I034_040(w_034_040, w_032_609, w_011_461);
  nand2 I034_041(w_034_041, w_003_026, w_018_016);
  nand2 I034_042(w_034_042, w_004_147, w_023_149);
  or2  I034_043(w_034_043, w_030_198, w_028_078);
  nand2 I034_044(w_034_044, w_007_440, w_018_020);
  not1 I034_045(w_034_045, w_026_196);
  or2  I034_046(w_034_046, w_021_160, w_001_010);
  nand2 I034_047(w_034_047, w_021_097, w_019_010);
  nand2 I034_048(w_034_048, w_003_056, w_004_109);
  and2 I034_049(w_034_049, w_002_044, w_021_211);
  or2  I034_050(w_034_050, w_015_351, w_012_089);
  and2 I034_051(w_034_051, w_004_408, w_020_069);
  and2 I034_052(w_034_052, w_011_592, w_024_073);
  and2 I034_053(w_034_053, w_018_042, w_025_137);
  not1 I034_054(w_034_054, w_020_450);
  nand2 I034_055(w_034_055, w_024_041, w_017_048);
  or2  I034_056(w_034_056, w_004_024, w_004_321);
  not1 I034_057(w_034_057, w_017_664);
  not1 I034_058(w_034_058, w_021_272);
  and2 I034_059(w_034_059, w_026_077, w_001_003);
  or2  I034_060(w_034_060, w_022_342, w_021_081);
  nand2 I034_061(w_034_061, w_032_210, w_025_097);
  or2  I034_062(w_034_062, w_024_227, w_006_084);
  and2 I034_063(w_034_063, w_010_677, w_009_322);
  nand2 I034_064(w_034_064, w_000_186, w_005_244);
  nand2 I034_065(w_034_065, w_021_163, w_004_028);
  and2 I034_066(w_034_066, w_007_031, w_021_208);
  or2  I034_067(w_034_067, w_026_439, w_016_003);
  not1 I034_068(w_034_068, w_031_276);
  or2  I034_069(w_034_069, w_004_066, w_008_686);
  nand2 I034_070(w_034_070, w_017_560, w_028_076);
  nand2 I034_071(w_034_071, w_033_426, w_020_428);
  and2 I034_072(w_034_072, w_032_457, w_023_129);
  not1 I034_073(w_034_073, w_010_466);
  nand2 I034_074(w_034_074, w_010_106, w_007_120);
  and2 I034_075(w_034_075, w_013_396, w_019_003);
  nand2 I035_000(w_035_000, w_023_008, w_023_154);
  or2  I035_001(w_035_001, w_031_453, w_008_610);
  nand2 I035_002(w_035_002, w_017_226, w_025_026);
  nand2 I035_003(w_035_003, w_023_100, w_002_267);
  nand2 I035_004(w_035_004, w_014_131, w_002_526);
  or2  I035_005(w_035_005, w_023_039, w_009_077);
  not1 I035_006(w_035_006, w_034_072);
  and2 I035_007(w_035_007, w_022_006, w_004_176);
  nand2 I035_008(w_035_008, w_013_048, w_016_003);
  not1 I035_009(w_035_009, w_018_040);
  not1 I035_010(w_035_010, w_007_235);
  nand2 I035_012(w_035_012, w_023_117, w_031_144);
  nand2 I035_013(w_035_013, w_033_011, w_017_051);
  nand2 I035_014(w_035_014, w_017_409, w_034_026);
  or2  I035_015(w_035_015, w_024_178, w_004_386);
  and2 I035_016(w_035_016, w_023_203, w_020_387);
  and2 I035_017(w_035_017, w_006_092, w_034_075);
  not1 I035_018(w_035_018, w_008_085);
  nand2 I035_019(w_035_019, w_004_390, w_013_318);
  or2  I035_020(w_035_020, w_031_112, w_025_280);
  not1 I035_021(w_035_021, w_024_190);
  nand2 I035_022(w_035_022, w_013_148, w_013_551);
  and2 I035_023(w_035_023, w_013_306, w_005_218);
  not1 I035_024(w_035_024, w_011_044);
  not1 I035_025(w_035_025, w_005_173);
  not1 I035_027(w_035_027, w_033_766);
  and2 I035_028(w_035_028, w_029_104, w_011_309);
  not1 I035_029(w_035_029, w_008_009);
  and2 I035_030(w_035_030, w_017_140, w_017_019);
  nand2 I035_031(w_035_031, w_002_040, w_029_072);
  or2  I035_032(w_035_032, w_032_073, w_011_046);
  not1 I035_034(w_035_034, w_034_027);
  not1 I035_035(w_035_035, w_005_091);
  nand2 I035_036(w_035_036, w_024_464, w_005_184);
  or2  I035_037(w_035_037, w_022_266, w_001_017);
  and2 I035_039(w_035_039, w_030_050, w_019_011);
  nand2 I035_040(w_035_040, w_010_516, w_030_055);
  and2 I035_042(w_035_042, w_011_280, w_024_537);
  and2 I035_043(w_035_043, w_030_273, w_033_319);
  or2  I035_044(w_035_044, w_000_559, w_033_685);
  not1 I035_045(w_035_045, w_031_488);
  nand2 I035_046(w_035_046, w_003_007, w_032_118);
  and2 I035_047(w_035_047, w_008_436, w_012_176);
  nand2 I035_048(w_035_048, w_018_037, w_014_245);
  or2  I035_049(w_035_049, w_004_279, w_007_361);
  or2  I035_050(w_035_050, w_005_042, w_012_182);
  nand2 I035_051(w_035_051, w_011_420, w_022_249);
  and2 I035_052(w_035_052, w_000_295, w_022_202);
  nand2 I035_053(w_035_053, w_027_042, w_001_033);
  or2  I035_054(w_035_054, w_023_112, w_009_048);
  not1 I035_055(w_035_055, w_014_269);
  not1 I035_056(w_035_056, w_033_182);
  nand2 I035_057(w_035_057, w_015_062, w_033_148);
  and2 I035_059(w_035_059, w_018_003, w_032_437);
  not1 I035_060(w_035_060, w_024_295);
  or2  I035_061(w_035_061, w_028_232, w_030_083);
  not1 I035_062(w_035_062, w_010_641);
  not1 I035_063(w_035_063, w_029_091);
  and2 I035_064(w_035_064, w_001_007, w_026_535);
  and2 I035_065(w_035_065, w_001_030, w_020_406);
  or2  I035_066(w_035_066, w_015_186, w_034_055);
  nand2 I035_067(w_035_067, w_027_011, w_018_014);
  nand2 I035_068(w_035_068, w_023_023, w_028_268);
  or2  I035_069(w_035_069, w_015_110, w_014_164);
  or2  I035_070(w_035_070, w_024_057, w_008_016);
  not1 I035_072(w_035_072, w_027_117);
  and2 I035_073(w_035_073, w_027_195, w_016_005);
  not1 I035_074(w_035_074, w_011_042);
  or2  I035_076(w_035_076, w_017_087, w_005_033);
  and2 I035_077(w_035_077, w_007_222, w_026_604);
  not1 I035_078(w_035_078, w_010_425);
  and2 I035_080(w_035_080, w_034_034, w_012_109);
  and2 I035_081(w_035_081, w_000_697, w_004_051);
  or2  I035_082(w_035_082, w_018_026, w_021_212);
  nand2 I035_083(w_035_083, w_027_142, w_022_044);
  or2  I035_084(w_035_084, w_013_026, w_033_289);
  nand2 I035_085(w_035_085, w_024_178, w_024_116);
  not1 I035_087(w_035_087, w_033_522);
  nand2 I035_088(w_035_088, w_014_125, w_003_065);
  or2  I035_090(w_035_090, w_029_000, w_016_005);
  or2  I035_091(w_035_091, w_030_108, w_031_231);
  nand2 I035_092(w_035_092, w_021_189, w_032_574);
  or2  I035_093(w_035_093, w_029_037, w_020_396);
  nand2 I035_094(w_035_094, w_018_020, w_025_037);
  nand2 I035_095(w_035_095, w_028_345, w_034_070);
  or2  I035_096(w_035_096, w_029_013, w_034_004);
  not1 I035_097(w_035_097, w_033_622);
  not1 I035_098(w_035_098, w_006_152);
  or2  I035_099(w_035_099, w_004_084, w_016_004);
  nand2 I035_100(w_035_100, w_010_006, w_030_288);
  or2  I035_101(w_035_101, w_025_001, w_019_004);
  or2  I035_102(w_035_102, w_025_039, w_034_042);
  nand2 I035_103(w_035_103, w_005_225, w_028_175);
  not1 I035_104(w_035_104, w_026_585);
  and2 I035_105(w_035_105, w_010_542, w_023_194);
  or2  I035_106(w_035_106, w_016_001, w_001_000);
  or2  I035_107(w_035_107, w_008_022, w_033_369);
  not1 I035_108(w_035_108, w_017_010);
  not1 I035_110(w_035_110, w_022_386);
  not1 I035_111(w_035_111, w_014_182);
  not1 I035_112(w_035_112, w_001_024);
  and2 I035_114(w_035_114, w_018_012, w_026_144);
  nand2 I035_115(w_035_115, w_029_052, w_006_112);
  or2  I035_116(w_035_116, w_024_312, w_015_442);
  nand2 I035_117(w_035_117, w_001_006, w_023_029);
  not1 I035_118(w_035_118, w_016_005);
  not1 I035_119(w_035_119, w_015_392);
  not1 I035_120(w_035_120, w_018_040);
  or2  I035_121(w_035_121, w_033_414, w_013_098);
  not1 I035_122(w_035_122, w_033_530);
  and2 I035_124(w_035_124, w_011_138, w_000_540);
  nand2 I035_125(w_035_125, w_024_265, w_017_663);
  or2  I035_126(w_035_126, w_006_081, w_027_123);
  nand2 I035_127(w_035_127, w_022_048, w_028_397);
  and2 I036_002(w_036_002, w_009_428, w_020_259);
  and2 I036_004(w_036_004, w_015_081, w_013_376);
  and2 I036_006(w_036_006, w_007_077, w_027_067);
  not1 I036_009(w_036_009, w_013_209);
  and2 I036_010(w_036_010, w_017_375, w_021_209);
  not1 I036_011(w_036_011, w_034_032);
  not1 I036_012(w_036_012, w_035_032);
  nand2 I036_014(w_036_014, w_035_017, w_003_008);
  nand2 I036_018(w_036_018, w_010_628, w_001_002);
  and2 I036_019(w_036_019, w_029_033, w_004_015);
  not1 I036_020(w_036_020, w_028_336);
  not1 I036_022(w_036_022, w_025_018);
  not1 I036_023(w_036_023, w_030_247);
  and2 I036_024(w_036_024, w_017_579, w_011_630);
  nand2 I036_026(w_036_026, w_028_038, w_005_242);
  not1 I036_028(w_036_028, w_010_606);
  not1 I036_029(w_036_029, w_014_277);
  and2 I036_032(w_036_032, w_017_315, w_034_075);
  nand2 I036_033(w_036_033, w_006_198, w_028_300);
  or2  I036_034(w_036_034, w_022_345, w_028_209);
  not1 I036_035(w_036_035, w_002_602);
  nand2 I036_037(w_036_037, w_026_070, w_026_105);
  not1 I036_039(w_036_039, w_020_157);
  and2 I036_042(w_036_042, w_010_121, w_013_134);
  or2  I036_043(w_036_043, w_029_093, w_004_115);
  or2  I036_044(w_036_044, w_030_145, w_011_175);
  and2 I036_046(w_036_046, w_017_667, w_017_168);
  not1 I036_047(w_036_047, w_014_286);
  not1 I036_049(w_036_049, w_018_020);
  nand2 I036_050(w_036_050, w_004_043, w_012_109);
  not1 I036_052(w_036_052, w_021_218);
  nand2 I036_053(w_036_053, w_030_123, w_000_141);
  or2  I036_058(w_036_058, w_026_708, w_031_143);
  not1 I036_059(w_036_059, w_014_120);
  and2 I036_060(w_036_060, w_031_111, w_012_116);
  nand2 I036_062(w_036_062, w_008_659, w_012_213);
  not1 I036_063(w_036_063, w_008_246);
  nand2 I036_064(w_036_064, w_017_069, w_020_586);
  or2  I036_066(w_036_066, w_017_524, w_032_144);
  and2 I036_068(w_036_068, w_016_000, w_022_395);
  nand2 I036_071(w_036_071, w_022_088, w_032_342);
  and2 I036_072(w_036_072, w_034_032, w_030_145);
  not1 I036_073(w_036_073, w_027_091);
  not1 I036_074(w_036_074, w_009_601);
  or2  I036_075(w_036_075, w_003_054, w_000_035);
  not1 I036_076(w_036_076, w_035_050);
  or2  I036_078(w_036_078, w_032_279, w_015_516);
  and2 I036_079(w_036_079, w_017_005, w_014_017);
  not1 I036_080(w_036_080, w_003_056);
  nand2 I036_082(w_036_082, w_017_222, w_023_101);
  and2 I036_083(w_036_083, w_002_299, w_033_160);
  and2 I036_084(w_036_084, w_021_205, w_017_042);
  and2 I036_085(w_036_085, w_012_078, w_024_221);
  nand2 I036_087(w_036_087, w_024_157, w_009_350);
  not1 I036_088(w_036_088, w_032_052);
  and2 I036_090(w_036_090, w_022_386, w_012_120);
  nand2 I036_091(w_036_091, w_009_384, w_028_277);
  not1 I036_093(w_036_093, w_033_209);
  or2  I036_094(w_036_094, w_021_224, w_031_027);
  or2  I036_096(w_036_096, w_034_073, w_029_085);
  nand2 I036_097(w_036_097, w_005_108, w_027_063);
  or2  I036_099(w_036_099, w_001_019, w_003_061);
  and2 I036_101(w_036_101, w_008_511, w_012_323);
  nand2 I036_103(w_036_103, w_026_657, w_007_049);
  and2 I036_109(w_036_109, w_014_136, w_011_072);
  and2 I036_110(w_036_110, w_034_071, w_034_036);
  not1 I036_112(w_036_112, w_013_153);
  nand2 I036_114(w_036_114, w_017_186, w_000_265);
  not1 I036_117(w_036_117, w_019_018);
  not1 I036_118(w_036_118, w_000_308);
  nand2 I036_120(w_036_120, w_012_187, w_010_222);
  or2  I036_121(w_036_121, w_022_331, w_026_321);
  or2  I036_123(w_036_123, w_021_097, w_020_068);
  and2 I036_125(w_036_125, w_029_035, w_026_288);
  nand2 I036_126(w_036_126, w_025_160, w_034_059);
  nand2 I036_128(w_036_128, w_013_067, w_020_536);
  and2 I036_129(w_036_129, w_030_051, w_029_035);
  nand2 I036_131(w_036_131, w_008_541, w_023_141);
  or2  I036_132(w_036_132, w_016_003, w_019_014);
  not1 I036_134(w_036_134, w_007_128);
  or2  I036_136(w_036_136, w_027_011, w_030_178);
  not1 I036_138(w_036_138, w_000_316);
  nand2 I036_139(w_036_139, w_016_006, w_014_140);
  nand2 I036_140(w_036_140, w_003_033, w_027_151);
  and2 I036_141(w_036_141, w_034_001, w_009_446);
  and2 I036_144(w_036_144, w_028_127, w_025_120);
  nand2 I036_146(w_036_146, w_019_001, w_034_070);
  not1 I036_148(w_036_148, w_001_010);
  not1 I036_151(w_036_151, w_030_149);
  and2 I036_153(w_036_153, w_007_439, w_026_489);
  nand2 I036_154(w_036_154, w_032_442, w_019_001);
  nand2 I036_156(w_036_156, w_015_428, w_011_195);
  and2 I036_157(w_036_157, w_016_002, w_030_163);
  and2 I036_158(w_036_158, w_030_117, w_005_095);
  or2  I036_160(w_036_160, w_003_025, w_008_207);
  and2 I036_161(w_036_161, w_027_002, w_028_279);
  and2 I036_162(w_036_162, w_008_708, w_007_195);
  and2 I036_163(w_036_163, w_035_102, w_028_171);
  or2  I036_164(w_036_164, w_003_082, w_025_288);
  nand2 I036_165(w_036_165, w_010_563, w_001_003);
  and2 I036_166(w_036_166, w_018_003, w_030_319);
  nand2 I036_170(w_036_170, w_014_024, w_020_529);
  or2  I036_173(w_036_173, w_033_647, w_015_464);
  not1 I036_175(w_036_175, w_033_745);
  or2  I036_177(w_036_177, w_008_367, w_030_070);
  or2  I036_178(w_036_178, w_020_132, w_022_384);
  not1 I036_179(w_036_179, w_001_012);
  nand2 I036_180(w_036_180, w_035_027, w_023_073);
  nand2 I036_182(w_036_182, w_005_254, w_035_003);
  and2 I036_186(w_036_186, w_033_653, w_020_320);
  or2  I036_188(w_036_188, w_008_202, w_014_083);
  or2  I036_190(w_036_190, w_001_013, w_017_572);
  nand2 I036_191(w_036_191, w_001_004, w_027_008);
  nand2 I036_192(w_036_192, w_003_054, w_029_069);
  or2  I036_194(w_036_194, w_031_174, w_015_629);
  not1 I036_197(w_036_197, w_026_441);
  or2  I036_200(w_036_200, w_011_176, w_026_366);
  not1 I036_201(w_036_201, w_006_196);
  or2  I036_206(w_036_206, w_007_037, w_030_291);
  or2  I036_207(w_036_207, w_000_657, w_031_105);
  nand2 I036_211(w_036_211, w_005_311, w_025_204);
  not1 I036_215(w_036_215, w_030_222);
  not1 I036_217(w_036_217, w_033_511);
  and2 I036_221(w_036_221, w_006_020, w_033_779);
  and2 I036_224(w_036_224, w_030_302, w_021_166);
  nand2 I036_227(w_036_227, w_033_555, w_035_027);
  or2  I036_229(w_036_229, w_011_618, w_031_380);
  nand2 I036_231(w_036_231, w_000_596, w_015_469);
  not1 I036_232(w_036_232, w_019_015);
  and2 I036_235(w_036_235, w_008_214, w_025_056);
  nand2 I036_237(w_036_237, w_004_340, w_022_012);
  not1 I036_239(w_036_239, w_006_215);
  nand2 I036_240(w_036_240, w_004_082, w_032_030);
  and2 I036_241(w_036_241, w_034_017, w_032_298);
  nand2 I036_242(w_036_242, w_022_296, w_027_115);
  nand2 I036_243(w_036_243, w_028_542, w_002_520);
  not1 I036_244(w_036_244, w_004_085);
  not1 I036_245(w_036_245, w_021_119);
  and2 I036_247(w_036_247, w_031_136, w_004_222);
  and2 I036_251(w_036_251, w_009_553, w_024_026);
  and2 I036_255(w_036_255, w_030_213, w_024_123);
  not1 I036_256(w_036_256, w_015_170);
  nand2 I036_257(w_036_257, w_008_561, w_016_001);
  or2  I036_258(w_036_258, w_025_204, w_034_016);
  nand2 I036_259(w_036_259, w_023_169, w_028_446);
  not1 I036_261(w_036_261, w_018_028);
  not1 I036_262(w_036_262, w_012_095);
  and2 I036_265(w_036_265, w_008_022, w_026_620);
  not1 I036_266(w_036_266, w_034_016);
  not1 I036_267(w_036_267, w_035_124);
  not1 I036_269(w_036_269, w_008_241);
  or2  I036_271(w_036_271, w_010_750, w_023_117);
  nand2 I036_272(w_036_272, w_010_027, w_012_238);
  or2  I036_273(w_036_273, w_008_061, w_003_064);
  nand2 I036_274(w_036_274, w_003_061, w_007_438);
  not1 I036_276(w_036_276, w_003_000);
  nand2 I036_277(w_036_277, w_008_571, w_024_079);
  or2  I036_278(w_036_278, w_027_182, w_017_094);
  not1 I036_281(w_036_281, w_023_092);
  not1 I036_282(w_036_282, w_008_137);
  and2 I036_283(w_036_283, w_017_435, w_024_268);
  not1 I036_284(w_036_284, w_032_391);
  not1 I036_286(w_036_286, w_020_363);
  and2 I036_289(w_036_289, w_022_259, w_020_099);
  and2 I036_291(w_036_291, w_028_088, w_019_005);
  nand2 I036_294(w_036_294, w_035_037, w_008_019);
  not1 I036_295(w_036_295, w_004_237);
  not1 I036_296(w_036_296, w_004_398);
  not1 I036_297(w_036_297, w_005_165);
  not1 I036_298(w_036_298, w_034_072);
  not1 I036_299(w_036_299, w_014_291);
  not1 I036_302(w_036_302, w_023_017);
  or2  I036_304(w_036_304, w_001_018, w_011_489);
  and2 I036_305(w_036_305, w_009_490, w_028_208);
  and2 I036_307(w_036_307, w_018_037, w_004_160);
  and2 I036_309(w_036_309, w_011_169, w_009_131);
  nand2 I036_310(w_036_310, w_026_050, w_032_575);
  not1 I036_311(w_036_311, w_007_264);
  not1 I036_312(w_036_312, w_016_000);
  not1 I036_313(w_036_313, w_019_020);
  nand2 I036_314(w_036_314, w_025_277, w_003_071);
  or2  I036_318(w_036_318, w_019_019, w_000_045);
  not1 I036_319(w_036_319, w_009_600);
  nand2 I036_322(w_036_322, w_023_031, w_008_082);
  nand2 I036_323(w_036_323, w_029_114, w_019_000);
  or2  I036_324(w_036_324, w_032_559, w_032_259);
  or2  I036_327(w_036_327, w_034_049, w_025_145);
  nand2 I036_328(w_036_328, w_011_550, w_018_003);
  and2 I036_330(w_036_330, w_034_033, w_030_163);
  and2 I036_335(w_036_335, w_017_649, w_032_109);
  not1 I036_336(w_036_336, w_010_686);
  or2  I036_348(w_036_348, w_007_060, w_021_100);
  nand2 I036_349(w_036_349, w_025_076, w_013_050);
  nand2 I036_350(w_036_350, w_034_021, w_023_031);
  nand2 I036_354(w_036_354, w_007_084, w_008_490);
  not1 I036_357(w_036_357, w_013_031);
  or2  I036_359(w_036_359, w_034_051, w_010_005);
  not1 I036_368(w_036_368, w_004_243);
  not1 I036_376(w_036_376, w_010_540);
  nand2 I036_386(w_036_386, w_010_006, w_017_463);
  and2 I036_393(w_036_393, w_017_458, w_004_066);
  not1 I036_395(w_036_395, w_013_069);
  not1 I036_400(w_036_400, w_033_201);
  and2 I036_404(w_036_404, w_017_116, w_029_008);
  or2  I036_408(w_036_408, w_008_261, w_005_041);
  or2  I036_412(w_036_412, w_027_134, w_000_184);
  and2 I036_430(w_036_430, w_023_159, w_003_005);
  nand2 I036_432(w_036_432, w_010_633, w_006_120);
  or2  I036_440(w_036_440, w_024_478, w_010_735);
  and2 I036_444(w_036_444, w_031_295, w_019_019);
  and2 I036_447(w_036_447, w_008_541, w_015_577);
  nand2 I036_449(w_036_449, w_024_166, w_030_312);
  not1 I036_455(w_036_455, w_033_087);
  nand2 I036_459(w_036_459, w_024_095, w_026_128);
  or2  I036_461(w_036_461, w_009_443, w_005_063);
  or2  I037_001(w_037_001, w_015_390, w_014_258);
  not1 I037_002(w_037_002, w_009_001);
  or2  I037_003(w_037_003, w_030_300, w_007_159);
  not1 I037_008(w_037_008, w_012_342);
  and2 I037_010(w_037_010, w_014_250, w_004_011);
  and2 I037_011(w_037_011, w_012_019, w_000_061);
  nand2 I037_013(w_037_013, w_024_018, w_031_129);
  nand2 I037_015(w_037_015, w_034_047, w_030_011);
  not1 I037_017(w_037_017, w_024_180);
  and2 I037_020(w_037_020, w_034_002, w_030_024);
  nand2 I037_021(w_037_021, w_031_460, w_009_020);
  nand2 I037_022(w_037_022, w_002_214, w_011_024);
  or2  I037_023(w_037_023, w_031_193, w_027_049);
  or2  I037_024(w_037_024, w_005_245, w_021_048);
  and2 I037_026(w_037_026, w_036_395, w_005_056);
  not1 I037_028(w_037_028, w_016_000);
  and2 I037_030(w_037_030, w_014_048, w_013_404);
  and2 I037_031(w_037_031, w_009_329, w_028_107);
  or2  I037_032(w_037_032, w_011_156, w_010_768);
  or2  I037_033(w_037_033, w_010_036, w_026_130);
  not1 I037_034(w_037_034, w_012_177);
  or2  I037_036(w_037_036, w_029_038, w_030_036);
  or2  I037_041(w_037_041, w_015_052, w_006_162);
  nand2 I037_042(w_037_042, w_024_214, w_025_152);
  and2 I037_044(w_037_044, w_032_364, w_003_084);
  not1 I037_045(w_037_045, w_033_566);
  not1 I037_047(w_037_047, w_034_048);
  and2 I037_048(w_037_048, w_012_076, w_023_131);
  not1 I037_049(w_037_049, w_010_551);
  or2  I037_050(w_037_050, w_009_384, w_031_014);
  not1 I037_051(w_037_051, w_017_531);
  or2  I037_055(w_037_055, w_016_006, w_020_225);
  not1 I037_059(w_037_059, w_030_320);
  or2  I037_060(w_037_060, w_015_007, w_025_294);
  and2 I037_062(w_037_062, w_024_473, w_025_069);
  not1 I037_063(w_037_063, w_018_016);
  and2 I037_064(w_037_064, w_012_026, w_000_497);
  and2 I037_066(w_037_066, w_013_160, w_009_515);
  nand2 I037_068(w_037_068, w_010_118, w_035_053);
  or2  I037_070(w_037_070, w_028_133, w_016_005);
  or2  I037_071(w_037_071, w_006_158, w_024_224);
  nand2 I037_073(w_037_073, w_003_042, w_017_132);
  nand2 I037_074(w_037_074, w_015_036, w_009_161);
  nand2 I037_075(w_037_075, w_013_249, w_013_080);
  and2 I037_076(w_037_076, w_011_545, w_025_037);
  nand2 I037_077(w_037_077, w_012_031, w_024_510);
  or2  I037_081(w_037_081, w_013_183, w_032_514);
  and2 I037_082(w_037_082, w_023_160, w_026_635);
  and2 I037_083(w_037_083, w_014_042, w_034_067);
  nand2 I037_085(w_037_085, w_000_129, w_014_218);
  and2 I037_086(w_037_086, w_017_189, w_018_040);
  or2  I037_087(w_037_087, w_009_329, w_005_157);
  nand2 I037_088(w_037_088, w_003_006, w_001_009);
  not1 I037_089(w_037_089, w_026_645);
  or2  I037_093(w_037_093, w_028_190, w_010_219);
  and2 I037_095(w_037_095, w_006_142, w_031_186);
  nand2 I037_096(w_037_096, w_031_253, w_027_061);
  or2  I037_097(w_037_097, w_026_649, w_000_165);
  not1 I037_100(w_037_100, w_026_152);
  nand2 I037_101(w_037_101, w_017_030, w_022_137);
  and2 I037_103(w_037_103, w_007_248, w_008_094);
  or2  I037_104(w_037_104, w_008_611, w_006_018);
  or2  I037_105(w_037_105, w_008_669, w_004_451);
  not1 I037_110(w_037_110, w_031_133);
  and2 I037_115(w_037_115, w_034_012, w_034_048);
  not1 I037_117(w_037_117, w_017_371);
  and2 I037_119(w_037_119, w_003_054, w_011_083);
  not1 I037_120(w_037_120, w_021_226);
  or2  I037_122(w_037_122, w_024_005, w_010_357);
  and2 I037_123(w_037_123, w_032_588, w_009_097);
  not1 I037_124(w_037_124, w_023_013);
  nand2 I037_129(w_037_129, w_014_220, w_011_087);
  not1 I037_130(w_037_130, w_021_243);
  and2 I037_131(w_037_131, w_011_472, w_034_041);
  and2 I037_132(w_037_132, w_003_037, w_013_105);
  or2  I037_133(w_037_133, w_035_101, w_007_017);
  and2 I037_140(w_037_140, w_015_433, w_025_095);
  not1 I037_141(w_037_141, w_012_130);
  or2  I037_146(w_037_146, w_021_097, w_016_006);
  nand2 I037_147(w_037_147, w_009_152, w_003_040);
  and2 I037_149(w_037_149, w_018_027, w_022_206);
  nand2 I037_150(w_037_150, w_022_271, w_019_010);
  or2  I037_152(w_037_152, w_012_171, w_017_086);
  nand2 I037_153(w_037_153, w_010_018, w_010_679);
  and2 I037_154(w_037_154, w_009_295, w_012_042);
  not1 I037_155(w_037_155, w_020_183);
  or2  I037_157(w_037_157, w_035_124, w_027_168);
  or2  I037_158(w_037_158, w_014_145, w_019_015);
  or2  I037_162(w_037_162, w_003_050, w_023_086);
  nand2 I037_164(w_037_164, w_012_120, w_000_576);
  or2  I037_166(w_037_166, w_029_046, w_028_575);
  nand2 I037_168(w_037_168, w_013_370, w_014_075);
  nand2 I037_169(w_037_169, w_018_010, w_015_113);
  and2 I037_172(w_037_172, w_019_008, w_026_490);
  and2 I037_173(w_037_173, w_018_032, w_013_186);
  nand2 I037_177(w_037_177, w_033_380, w_025_297);
  nand2 I037_185(w_037_185, w_027_182, w_023_143);
  and2 I037_186(w_037_186, w_025_060, w_033_015);
  or2  I037_188(w_037_188, w_036_232, w_002_414);
  or2  I037_189(w_037_189, w_016_002, w_033_725);
  not1 I037_195(w_037_195, w_022_115);
  and2 I037_198(w_037_198, w_000_641, w_008_077);
  nand2 I037_200(w_037_200, w_028_139, w_010_087);
  or2  I037_201(w_037_201, w_021_051, w_028_517);
  nand2 I037_203(w_037_203, w_012_049, w_002_048);
  not1 I037_206(w_037_206, w_034_074);
  or2  I037_207(w_037_207, w_029_007, w_030_196);
  or2  I037_208(w_037_208, w_011_514, w_006_221);
  or2  I037_210(w_037_210, w_024_107, w_034_008);
  not1 I037_211(w_037_211, w_032_057);
  and2 I037_212(w_037_212, w_017_019, w_001_010);
  and2 I037_217(w_037_217, w_021_095, w_018_043);
  nand2 I037_218(w_037_218, w_035_063, w_033_331);
  not1 I037_221(w_037_221, w_025_072);
  not1 I037_223(w_037_223, w_025_131);
  or2  I037_225(w_037_225, w_033_583, w_014_203);
  not1 I037_228(w_037_228, w_006_226);
  not1 I037_229(w_037_229, w_000_763);
  and2 I037_231(w_037_231, w_024_089, w_009_297);
  nand2 I037_232(w_037_232, w_006_080, w_012_048);
  or2  I037_233(w_037_233, w_019_008, w_002_076);
  nand2 I037_234(w_037_234, w_021_241, w_022_262);
  or2  I037_235(w_037_235, w_007_040, w_030_305);
  nand2 I037_236(w_037_236, w_026_118, w_028_224);
  or2  I037_242(w_037_242, w_015_260, w_001_006);
  or2  I037_245(w_037_245, w_011_490, w_017_543);
  or2  I037_246(w_037_246, w_000_159, w_021_241);
  and2 I037_248(w_037_248, w_001_019, w_005_239);
  and2 I037_249(w_037_249, w_022_131, w_016_008);
  nand2 I037_251(w_037_251, w_013_295, w_020_307);
  not1 I037_253(w_037_253, w_004_162);
  not1 I037_257(w_037_257, w_020_450);
  not1 I037_258(w_037_258, w_011_502);
  or2  I037_261(w_037_261, w_027_036, w_002_624);
  or2  I037_262(w_037_262, w_012_015, w_009_265);
  nand2 I037_263(w_037_263, w_030_168, w_006_135);
  not1 I037_266(w_037_266, w_001_011);
  nand2 I037_267(w_037_267, w_019_006, w_027_082);
  or2  I037_268(w_037_268, w_032_138, w_018_017);
  and2 I037_273(w_037_273, w_023_073, w_023_019);
  nand2 I037_277(w_037_277, w_023_017, w_029_096);
  and2 I037_278(w_037_278, w_031_548, w_032_163);
  and2 I037_279(w_037_279, w_026_585, w_009_101);
  or2  I037_280(w_037_280, w_033_658, w_035_044);
  or2  I037_285(w_037_285, w_004_464, w_016_002);
  or2  I037_286(w_037_286, w_026_491, w_024_142);
  or2  I037_287(w_037_287, w_000_574, w_034_012);
  and2 I037_293(w_037_293, w_029_062, w_003_069);
  not1 I037_295(w_037_295, w_021_042);
  or2  I037_300(w_037_300, w_019_003, w_022_214);
  nand2 I037_301(w_037_301, w_029_021, w_007_134);
  or2  I037_302(w_037_302, w_015_190, w_033_365);
  not1 I037_303(w_037_303, w_001_017);
  not1 I037_305(w_037_305, w_031_366);
  nand2 I037_308(w_037_308, w_008_172, w_029_064);
  not1 I037_309(w_037_309, w_008_479);
  not1 I037_310(w_037_310, w_017_016);
  nand2 I037_312(w_037_312, w_016_007, w_005_099);
  and2 I037_313(w_037_313, w_016_002, w_008_020);
  or2  I037_314(w_037_314, w_021_081, w_017_033);
  and2 I037_315(w_037_315, w_025_119, w_022_362);
  not1 I037_316(w_037_316, w_008_041);
  not1 I037_318(w_037_318, w_001_009);
  or2  I037_319(w_037_319, w_032_583, w_020_269);
  nand2 I037_320(w_037_320, w_036_310, w_021_219);
  nand2 I037_323(w_037_323, w_034_033, w_027_131);
  nand2 I037_330(w_037_330, w_025_035, w_028_132);
  nand2 I037_332(w_037_332, w_004_175, w_003_079);
  nand2 I037_333(w_037_333, w_032_546, w_029_072);
  nand2 I037_336(w_037_336, w_029_102, w_013_445);
  nand2 I037_338(w_037_338, w_027_178, w_022_399);
  not1 I037_339(w_037_339, w_009_572);
  and2 I037_343(w_037_343, w_006_202, w_030_231);
  nand2 I037_345(w_037_345, w_005_141, w_003_019);
  nand2 I037_346(w_037_346, w_029_067, w_019_009);
  and2 I037_348(w_037_350, w_024_086, w_037_349);
  and2 I037_349(w_037_351, w_028_433, w_037_350);
  or2  I037_350(w_037_349, w_022_132, w_037_351);
  and2 I038_000(w_038_000, w_027_073, w_034_065);
  not1 I038_002(w_038_002, w_004_056);
  not1 I038_005(w_038_005, w_006_016);
  nand2 I038_011(w_038_011, w_011_022, w_035_042);
  not1 I038_012(w_038_012, w_012_062);
  or2  I038_016(w_038_016, w_033_379, w_002_419);
  or2  I038_018(w_038_018, w_037_185, w_018_007);
  and2 I038_019(w_038_019, w_030_264, w_015_265);
  and2 I038_020(w_038_020, w_032_434, w_029_060);
  not1 I038_021(w_038_021, w_008_298);
  nand2 I038_022(w_038_022, w_028_039, w_024_445);
  not1 I038_024(w_038_024, w_026_286);
  nand2 I038_025(w_038_025, w_003_020, w_007_285);
  and2 I038_032(w_038_032, w_019_015, w_032_175);
  nand2 I038_033(w_038_033, w_025_217, w_020_407);
  and2 I038_043(w_038_043, w_032_596, w_028_121);
  and2 I038_044(w_038_044, w_026_174, w_001_010);
  or2  I038_047(w_038_047, w_032_114, w_007_275);
  not1 I038_051(w_038_051, w_021_006);
  nand2 I038_052(w_038_052, w_005_107, w_010_479);
  or2  I038_053(w_038_053, w_007_261, w_024_387);
  and2 I038_054(w_038_054, w_018_025, w_026_033);
  or2  I038_055(w_038_055, w_032_249, w_037_089);
  or2  I038_059(w_038_059, w_011_139, w_025_160);
  not1 I038_061(w_038_061, w_000_605);
  or2  I038_064(w_038_064, w_006_189, w_036_042);
  and2 I038_065(w_038_065, w_037_345, w_015_024);
  and2 I038_066(w_038_066, w_002_414, w_035_096);
  or2  I038_067(w_038_067, w_031_508, w_012_036);
  or2  I038_068(w_038_068, w_017_482, w_008_292);
  or2  I038_070(w_038_070, w_030_417, w_028_118);
  not1 I038_074(w_038_074, w_032_257);
  or2  I038_076(w_038_076, w_004_128, w_027_083);
  or2  I038_077(w_038_077, w_013_011, w_036_099);
  and2 I038_079(w_038_079, w_016_006, w_001_004);
  and2 I038_082(w_038_082, w_004_231, w_004_184);
  and2 I038_085(w_038_085, w_012_012, w_003_081);
  or2  I038_087(w_038_087, w_017_416, w_010_742);
  not1 I038_090(w_038_090, w_014_122);
  nand2 I038_093(w_038_093, w_017_020, w_012_029);
  not1 I038_095(w_038_095, w_001_025);
  not1 I038_096(w_038_096, w_030_208);
  not1 I038_097(w_038_097, w_033_568);
  and2 I038_099(w_038_099, w_009_041, w_003_014);
  and2 I038_100(w_038_100, w_008_061, w_030_302);
  or2  I038_103(w_038_103, w_026_665, w_016_007);
  or2  I038_106(w_038_106, w_015_057, w_012_137);
  not1 I038_108(w_038_108, w_036_197);
  not1 I038_111(w_038_111, w_006_174);
  not1 I038_115(w_038_115, w_018_036);
  not1 I038_116(w_038_116, w_025_186);
  or2  I038_117(w_038_117, w_011_134, w_037_278);
  or2  I038_120(w_038_120, w_032_041, w_030_242);
  or2  I038_121(w_038_121, w_029_049, w_007_055);
  not1 I038_123(w_038_123, w_005_052);
  nand2 I038_132(w_038_132, w_029_072, w_023_025);
  and2 I038_134(w_038_134, w_021_259, w_015_277);
  or2  I038_135(w_038_135, w_006_032, w_008_225);
  and2 I038_138(w_038_138, w_018_025, w_022_129);
  nand2 I038_140(w_038_140, w_019_018, w_027_163);
  nand2 I038_142(w_038_142, w_001_020, w_018_024);
  not1 I038_143(w_038_143, w_030_071);
  or2  I038_144(w_038_144, w_029_038, w_023_087);
  nand2 I038_146(w_038_146, w_012_305, w_006_244);
  not1 I038_147(w_038_147, w_012_310);
  and2 I038_148(w_038_148, w_001_000, w_033_163);
  not1 I038_149(w_038_149, w_012_032);
  not1 I038_150(w_038_150, w_017_286);
  and2 I038_151(w_038_151, w_028_035, w_016_001);
  and2 I038_152(w_038_152, w_025_291, w_002_686);
  nand2 I038_157(w_038_157, w_030_161, w_017_031);
  or2  I038_160(w_038_160, w_020_251, w_023_142);
  or2  I038_162(w_038_162, w_037_026, w_032_525);
  or2  I038_163(w_038_163, w_025_131, w_032_134);
  nand2 I038_164(w_038_164, w_004_282, w_034_075);
  or2  I038_169(w_038_169, w_025_219, w_035_039);
  and2 I038_173(w_038_173, w_030_354, w_002_464);
  nand2 I038_176(w_038_176, w_002_068, w_029_039);
  and2 I038_178(w_038_178, w_034_020, w_032_092);
  nand2 I038_182(w_038_182, w_019_019, w_035_034);
  not1 I038_185(w_038_185, w_021_078);
  or2  I038_188(w_038_188, w_032_346, w_006_167);
  nand2 I038_193(w_038_193, w_015_281, w_034_007);
  not1 I038_196(w_038_196, w_011_060);
  not1 I038_200(w_038_200, w_017_179);
  not1 I038_203(w_038_203, w_029_045);
  or2  I038_211(w_038_211, w_022_145, w_033_447);
  or2  I038_225(w_038_225, w_011_491, w_030_385);
  nand2 I038_234(w_038_234, w_037_262, w_015_399);
  nand2 I038_240(w_038_240, w_004_290, w_004_039);
  and2 I038_247(w_038_247, w_015_224, w_022_296);
  nand2 I038_255(w_038_255, w_001_002, w_003_042);
  nand2 I038_256(w_038_256, w_034_065, w_017_247);
  and2 I038_260(w_038_260, w_033_436, w_010_678);
  or2  I038_265(w_038_265, w_007_289, w_024_311);
  nand2 I038_268(w_038_268, w_016_001, w_017_270);
  nand2 I038_275(w_038_275, w_034_044, w_004_196);
  not1 I038_285(w_038_285, w_037_081);
  nand2 I038_288(w_038_288, w_006_098, w_001_034);
  not1 I038_290(w_038_290, w_003_036);
  and2 I038_297(w_038_297, w_019_001, w_027_111);
  or2  I038_298(w_038_298, w_037_285, w_028_026);
  and2 I038_299(w_038_299, w_014_009, w_024_358);
  and2 I038_302(w_038_302, w_024_342, w_017_002);
  nand2 I038_303(w_038_303, w_021_249, w_033_002);
  not1 I038_304(w_038_304, w_004_405);
  or2  I038_308(w_038_308, w_037_198, w_003_061);
  nand2 I038_311(w_038_311, w_037_030, w_009_048);
  or2  I038_315(w_038_315, w_033_269, w_000_531);
  not1 I038_317(w_038_317, w_028_099);
  not1 I038_321(w_038_321, w_019_010);
  and2 I038_322(w_038_322, w_036_235, w_034_049);
  and2 I038_325(w_038_325, w_009_078, w_004_456);
  nand2 I038_331(w_038_331, w_036_207, w_031_127);
  or2  I038_333(w_038_333, w_000_553, w_010_122);
  and2 I038_337(w_038_337, w_018_040, w_005_018);
  nand2 I038_340(w_038_340, w_004_092, w_013_046);
  not1 I038_358(w_038_358, w_023_011);
  nand2 I038_359(w_038_359, w_023_096, w_005_191);
  nand2 I038_365(w_038_365, w_032_429, w_014_145);
  or2  I038_368(w_038_368, w_022_158, w_020_077);
  nand2 I038_370(w_038_370, w_015_172, w_001_009);
  not1 I038_377(w_038_377, w_034_017);
  and2 I038_383(w_038_383, w_010_556, w_015_447);
  and2 I038_385(w_038_385, w_025_221, w_003_009);
  or2  I038_386(w_038_386, w_000_133, w_031_034);
  or2  I038_396(w_038_396, w_037_087, w_012_325);
  nand2 I038_397(w_038_397, w_011_620, w_003_083);
  nand2 I038_402(w_038_402, w_033_715, w_011_095);
  or2  I038_405(w_038_405, w_012_187, w_019_002);
  and2 I038_415(w_038_415, w_031_548, w_014_135);
  nand2 I038_418(w_038_418, w_024_444, w_012_271);
  and2 I038_423(w_038_423, w_008_170, w_012_201);
  not1 I038_429(w_038_429, w_017_012);
  not1 I038_431(w_038_431, w_009_036);
  and2 I038_434(w_038_434, w_025_072, w_005_057);
  or2  I038_435(w_038_435, w_028_244, w_016_002);
  and2 I038_447(w_038_447, w_009_272, w_030_290);
  nand2 I038_454(w_038_454, w_028_402, w_020_216);
  and2 I038_455(w_038_455, w_002_706, w_016_003);
  nand2 I038_456(w_038_456, w_018_031, w_028_325);
  nand2 I038_457(w_038_457, w_007_025, w_027_155);
  or2  I038_458(w_038_458, w_008_711, w_005_313);
  and2 I038_462(w_038_462, w_005_083, w_024_435);
  or2  I038_465(w_038_465, w_000_196, w_029_075);
  or2  I038_467(w_038_467, w_000_393, w_007_107);
  not1 I038_468(w_038_468, w_001_001);
  nand2 I038_469(w_038_469, w_006_239, w_023_217);
  not1 I038_471(w_038_471, w_036_139);
  and2 I038_472(w_038_472, w_036_349, w_025_088);
  and2 I038_484(w_038_484, w_024_175, w_037_119);
  nand2 I038_486(w_038_486, w_013_133, w_004_025);
  or2  I038_489(w_038_489, w_020_511, w_000_520);
  not1 I038_491(w_038_491, w_020_132);
  or2  I038_495(w_038_495, w_021_209, w_037_201);
  and2 I038_496(w_038_496, w_018_037, w_023_193);
  and2 I038_498(w_038_498, w_004_450, w_016_002);
  not1 I038_499(w_038_499, w_018_026);
  not1 I038_501(w_038_501, w_016_003);
  or2  I038_503(w_038_503, w_011_276, w_026_451);
  nand2 I038_504(w_038_504, w_036_291, w_005_256);
  not1 I038_505(w_038_505, w_025_088);
  not1 I038_508(w_038_508, w_021_213);
  not1 I038_512(w_038_512, w_002_446);
  not1 I038_515(w_038_515, w_026_380);
  not1 I038_516(w_038_516, w_034_053);
  not1 I038_521(w_038_521, w_017_111);
  nand2 I038_526(w_038_526, w_007_166, w_016_006);
  or2  I038_531(w_038_531, w_002_193, w_006_095);
  nand2 I038_532(w_038_532, w_001_033, w_012_294);
  nand2 I038_538(w_038_538, w_012_344, w_024_230);
  not1 I038_542(w_038_542, w_031_462);
  or2  I038_546(w_038_546, w_013_100, w_030_004);
  not1 I038_548(w_038_548, w_007_092);
  and2 I038_549(w_038_549, w_001_011, w_025_174);
  not1 I038_550(w_038_550, w_008_145);
  not1 I038_551(w_038_551, w_023_115);
  nand2 I038_559(w_038_559, w_001_010, w_032_083);
  not1 I038_565(w_038_565, w_005_053);
  not1 I038_567(w_038_567, w_029_109);
  or2  I038_575(w_038_575, w_030_295, w_018_036);
  not1 I038_588(w_038_588, w_022_310);
  not1 I038_589(w_038_589, w_010_570);
  nand2 I038_590(w_038_590, w_028_096, w_009_597);
  and2 I038_591(w_038_591, w_010_084, w_013_265);
  nand2 I038_597(w_038_597, w_037_185, w_010_400);
  not1 I038_598(w_038_598, w_001_036);
  not1 I038_600(w_038_600, w_027_066);
  or2  I038_601(w_038_601, w_006_189, w_033_726);
  and2 I038_602(w_038_602, w_012_104, w_031_483);
  and2 I038_604(w_038_604, w_028_409, w_028_248);
  or2  I038_606(w_038_606, w_021_117, w_008_117);
  or2  I038_610(w_038_610, w_017_437, w_036_239);
  nand2 I038_618(w_038_618, w_008_367, w_030_202);
  nand2 I038_623(w_038_625, w_038_624, w_025_191);
  or2  I038_624(w_038_626, w_005_216, w_038_625);
  not1 I038_625(w_038_627, w_038_626);
  not1 I038_626(w_038_628, w_038_627);
  and2 I038_627(w_038_629, w_038_628, w_011_438);
  or2  I038_628(w_038_630, w_001_026, w_038_629);
  and2 I038_629(w_038_631, w_026_201, w_038_630);
  and2 I038_630(w_038_632, w_023_217, w_038_631);
  or2  I038_631(w_038_624, w_018_038, w_038_632);
  nand2 I039_003(w_039_003, w_002_233, w_038_051);
  and2 I039_005(w_039_005, w_005_027, w_026_519);
  not1 I039_007(w_039_007, w_037_049);
  or2  I039_010(w_039_010, w_031_528, w_035_066);
  nand2 I039_014(w_039_014, w_024_496, w_023_078);
  and2 I039_016(w_039_016, w_023_166, w_026_514);
  not1 I039_024(w_039_024, w_000_283);
  not1 I039_029(w_039_029, w_025_072);
  or2  I039_030(w_039_030, w_011_062, w_034_025);
  nand2 I039_032(w_039_032, w_002_661, w_024_026);
  not1 I039_033(w_039_033, w_038_096);
  nand2 I039_035(w_039_035, w_017_004, w_003_063);
  nand2 I039_037(w_039_037, w_019_002, w_032_398);
  nand2 I039_039(w_039_039, w_017_371, w_016_007);
  not1 I039_040(w_039_040, w_034_023);
  or2  I039_043(w_039_043, w_030_201, w_034_070);
  or2  I039_046(w_039_046, w_008_072, w_024_210);
  and2 I039_050(w_039_050, w_004_023, w_013_263);
  not1 I039_051(w_039_051, w_016_002);
  not1 I039_052(w_039_052, w_000_573);
  nand2 I039_054(w_039_054, w_023_099, w_034_066);
  not1 I039_055(w_039_055, w_017_552);
  not1 I039_057(w_039_057, w_002_268);
  not1 I039_061(w_039_061, w_034_071);
  not1 I039_063(w_039_063, w_036_166);
  not1 I039_064(w_039_064, w_036_063);
  not1 I039_066(w_039_066, w_029_014);
  and2 I039_068(w_039_068, w_032_520, w_017_453);
  or2  I039_069(w_039_069, w_003_017, w_002_620);
  or2  I039_072(w_039_072, w_018_030, w_036_412);
  or2  I039_073(w_039_073, w_026_217, w_010_499);
  or2  I039_076(w_039_076, w_016_001, w_036_163);
  or2  I039_078(w_039_078, w_032_254, w_009_492);
  not1 I039_079(w_039_079, w_034_029);
  not1 I039_082(w_039_082, w_034_043);
  or2  I039_085(w_039_085, w_007_141, w_012_275);
  not1 I039_088(w_039_088, w_026_028);
  and2 I039_089(w_039_089, w_010_500, w_023_025);
  or2  I039_092(w_039_092, w_010_414, w_002_118);
  nand2 I039_093(w_039_093, w_033_021, w_018_016);
  or2  I039_095(w_039_095, w_021_201, w_010_224);
  nand2 I039_099(w_039_099, w_020_196, w_025_165);
  not1 I039_103(w_039_103, w_016_004);
  not1 I039_104(w_039_104, w_009_502);
  nand2 I039_108(w_039_108, w_011_120, w_003_022);
  not1 I039_111(w_039_111, w_010_008);
  and2 I039_117(w_039_117, w_002_552, w_014_191);
  and2 I039_119(w_039_119, w_002_520, w_030_360);
  not1 I039_121(w_039_121, w_009_448);
  or2  I039_127(w_039_127, w_020_011, w_007_179);
  nand2 I039_141(w_039_141, w_036_256, w_031_330);
  and2 I039_143(w_039_143, w_004_373, w_013_527);
  nand2 I039_145(w_039_145, w_028_034, w_037_041);
  not1 I039_148(w_039_148, w_011_011);
  or2  I039_152(w_039_152, w_024_139, w_021_233);
  nand2 I039_155(w_039_155, w_027_173, w_025_201);
  not1 I039_158(w_039_158, w_035_006);
  nand2 I039_160(w_039_160, w_017_066, w_036_138);
  nand2 I039_161(w_039_161, w_024_262, w_025_040);
  not1 I039_167(w_039_167, w_024_003);
  nand2 I039_170(w_039_170, w_003_033, w_020_067);
  not1 I039_173(w_039_173, w_032_052);
  and2 I039_175(w_039_175, w_024_129, w_034_050);
  and2 I039_182(w_039_182, w_022_307, w_026_394);
  and2 I039_185(w_039_185, w_017_322, w_003_032);
  nand2 I039_187(w_039_187, w_015_128, w_035_090);
  or2  I039_197(w_039_197, w_035_018, w_019_020);
  not1 I039_203(w_039_203, w_035_016);
  nand2 I039_206(w_039_206, w_009_571, w_036_062);
  and2 I039_208(w_039_208, w_004_059, w_007_157);
  or2  I039_213(w_039_213, w_006_146, w_008_726);
  and2 I039_214(w_039_214, w_036_047, w_034_041);
  nand2 I039_218(w_039_218, w_033_535, w_035_087);
  not1 I039_219(w_039_219, w_005_236);
  not1 I039_221(w_039_221, w_018_013);
  and2 I039_228(w_039_228, w_012_034, w_011_515);
  and2 I039_231(w_039_231, w_008_408, w_038_163);
  nand2 I039_240(w_039_240, w_017_184, w_033_745);
  or2  I039_242(w_039_242, w_026_216, w_013_363);
  or2  I039_256(w_039_256, w_005_174, w_004_210);
  nand2 I039_258(w_039_258, w_015_086, w_013_075);
  or2  I039_260(w_039_260, w_016_006, w_033_021);
  or2  I039_263(w_039_263, w_011_430, w_038_044);
  nand2 I039_264(w_039_264, w_007_332, w_005_270);
  and2 I039_267(w_039_267, w_038_169, w_016_003);
  or2  I039_278(w_039_278, w_024_157, w_010_191);
  and2 I039_280(w_039_280, w_036_276, w_022_205);
  nand2 I039_289(w_039_289, w_023_005, w_036_286);
  and2 I039_295(w_039_295, w_017_424, w_027_159);
  nand2 I039_300(w_039_300, w_030_057, w_014_045);
  and2 I039_301(w_039_301, w_025_057, w_005_238);
  not1 I039_302(w_039_302, w_017_146);
  nand2 I039_306(w_039_306, w_025_236, w_028_181);
  not1 I039_309(w_039_309, w_028_045);
  or2  I039_317(w_039_317, w_037_146, w_037_318);
  nand2 I039_318(w_039_318, w_006_184, w_009_125);
  or2  I039_324(w_039_324, w_008_126, w_001_030);
  or2  I039_327(w_039_327, w_007_307, w_015_126);
  not1 I039_329(w_039_329, w_005_181);
  or2  I039_348(w_039_348, w_012_061, w_002_531);
  nand2 I039_351(w_039_351, w_012_201, w_018_011);
  nand2 I039_352(w_039_352, w_003_050, w_032_243);
  nand2 I039_360(w_039_360, w_036_059, w_010_341);
  or2  I039_361(w_039_361, w_020_599, w_014_062);
  nand2 I039_367(w_039_367, w_031_058, w_012_260);
  nand2 I039_368(w_039_368, w_021_059, w_012_276);
  and2 I039_370(w_039_370, w_033_653, w_014_185);
  or2  I039_371(w_039_371, w_025_051, w_031_074);
  not1 I039_372(w_039_372, w_015_234);
  nand2 I039_373(w_039_373, w_003_050, w_017_374);
  not1 I039_374(w_039_374, w_037_085);
  nand2 I039_377(w_039_377, w_006_180, w_022_369);
  not1 I039_380(w_039_380, w_034_057);
  nand2 I039_383(w_039_383, w_020_142, w_006_070);
  nand2 I039_395(w_039_395, w_033_289, w_036_072);
  or2  I039_396(w_039_396, w_030_311, w_038_117);
  nand2 I039_401(w_039_401, w_000_211, w_016_007);
  nand2 I039_404(w_039_404, w_008_489, w_013_186);
  nand2 I039_406(w_039_406, w_014_153, w_014_197);
  not1 I039_413(w_039_413, w_005_295);
  nand2 I039_415(w_039_415, w_015_524, w_036_259);
  or2  I039_421(w_039_421, w_015_118, w_004_096);
  not1 I039_422(w_039_422, w_008_620);
  not1 I039_424(w_039_424, w_027_004);
  not1 I039_425(w_039_425, w_027_187);
  and2 I039_427(w_039_427, w_010_454, w_013_032);
  not1 I039_428(w_039_428, w_033_769);
  not1 I039_429(w_039_429, w_008_403);
  not1 I039_432(w_039_432, w_034_040);
  not1 I039_440(w_039_440, w_014_067);
  not1 I039_446(w_039_446, w_036_444);
  or2  I039_448(w_039_448, w_031_362, w_032_466);
  and2 I039_459(w_039_459, w_026_201, w_023_105);
  nand2 I039_466(w_039_466, w_032_504, w_009_027);
  or2  I039_470(w_039_470, w_018_032, w_000_155);
  and2 I039_471(w_039_471, w_019_017, w_023_143);
  or2  I039_478(w_039_478, w_009_198, w_004_418);
  not1 I039_492(w_039_492, w_000_653);
  nand2 I039_493(w_039_493, w_013_123, w_031_151);
  not1 I039_495(w_039_495, w_025_281);
  nand2 I039_505(w_039_505, w_035_115, w_022_293);
  not1 I039_506(w_039_506, w_010_397);
  nand2 I039_510(w_039_510, w_013_128, w_036_242);
  nand2 I039_513(w_039_513, w_024_044, w_010_698);
  or2  I039_515(w_039_515, w_036_044, w_007_387);
  nand2 I039_518(w_039_518, w_014_212, w_009_318);
  or2  I039_519(w_039_519, w_032_348, w_000_709);
  or2  I039_522(w_039_522, w_026_026, w_019_006);
  nand2 I039_524(w_039_524, w_017_374, w_038_085);
  not1 I039_527(w_039_527, w_033_751);
  or2  I039_528(w_039_528, w_023_172, w_001_028);
  not1 I039_530(w_039_530, w_010_232);
  nand2 I039_534(w_039_534, w_029_047, w_006_249);
  and2 I039_536(w_039_536, w_029_017, w_006_027);
  not1 I039_537(w_039_537, w_032_411);
  or2  I039_538(w_039_538, w_026_149, w_024_347);
  not1 I039_539(w_039_539, w_022_237);
  and2 I039_543(w_039_543, w_028_536, w_013_222);
  nand2 I039_544(w_039_544, w_010_484, w_038_565);
  nand2 I039_550(w_039_550, w_007_118, w_014_071);
  not1 I039_552(w_039_552, w_010_012);
  nand2 I039_553(w_039_553, w_013_200, w_014_096);
  nand2 I039_559(w_039_559, w_022_348, w_015_003);
  and2 I039_561(w_039_561, w_005_010, w_014_149);
  not1 I039_567(w_039_567, w_023_103);
  and2 I039_569(w_039_569, w_013_220, w_031_012);
  not1 I039_571(w_039_571, w_035_046);
  nand2 I039_578(w_039_578, w_025_054, w_005_227);
  nand2 I039_580(w_039_580, w_022_082, w_031_467);
  not1 I039_581(w_039_581, w_038_090);
  nand2 I039_586(w_039_586, w_014_146, w_025_140);
  or2  I039_588(w_039_588, w_008_466, w_002_518);
  or2  I039_598(w_039_598, w_002_450, w_015_600);
  and2 I039_599(w_039_599, w_038_275, w_038_016);
  and2 I039_600(w_039_600, w_025_269, w_028_003);
  or2  I039_602(w_039_602, w_038_546, w_005_286);
  or2  I039_604(w_039_604, w_031_290, w_016_005);
  or2  I039_606(w_039_606, w_009_328, w_025_204);
  nand2 I039_609(w_039_609, w_011_214, w_035_020);
  and2 I039_612(w_039_612, w_027_140, w_023_178);
  or2  I039_616(w_039_616, w_006_081, w_032_049);
  not1 I039_620(w_039_620, w_001_005);
  not1 I039_621(w_039_621, w_031_439);
  not1 I039_625(w_039_625, w_021_043);
  or2  I039_634(w_039_634, w_012_333, w_037_129);
  and2 I039_646(w_039_646, w_032_154, w_025_124);
  not1 I039_648(w_039_648, w_024_284);
  nand2 I039_650(w_039_650, w_010_556, w_033_366);
  not1 I039_652(w_039_652, w_029_028);
  nand2 I039_656(w_039_656, w_024_097, w_013_323);
  and2 I039_657(w_039_657, w_023_213, w_035_106);
  or2  I039_658(w_039_658, w_017_030, w_035_078);
  or2  I039_667(w_039_667, w_001_011, w_009_230);
  not1 I039_668(w_039_668, w_006_082);
  and2 I039_676(w_039_676, w_019_004, w_030_040);
  not1 I039_680(w_039_680, w_013_201);
  nand2 I039_681(w_039_681, w_010_414, w_003_066);
  not1 I039_697(w_039_697, w_016_002);
  or2  I039_699(w_039_699, w_027_009, w_027_116);
  nand2 I039_706(w_039_706, w_037_280, w_002_191);
  or2  I039_708(w_039_708, w_011_350, w_004_158);
  nand2 I039_710(w_039_710, w_013_029, w_025_155);
  or2  I039_713(w_039_713, w_014_175, w_012_142);
  nand2 I039_714(w_039_714, w_026_152, w_027_093);
  or2  I039_718(w_039_718, w_023_075, w_003_045);
  or2  I039_719(w_039_719, w_004_192, w_012_277);
  and2 I040_000(w_040_000, w_030_100, w_006_071);
  or2  I040_004(w_040_004, w_015_402, w_005_029);
  nand2 I040_005(w_040_005, w_026_004, w_019_011);
  nand2 I040_008(w_040_008, w_020_021, w_014_076);
  or2  I040_012(w_040_012, w_013_151, w_035_054);
  or2  I040_013(w_040_013, w_002_580, w_014_071);
  nand2 I040_014(w_040_014, w_033_220, w_012_058);
  or2  I040_015(w_040_015, w_027_148, w_029_060);
  nand2 I040_017(w_040_017, w_019_006, w_002_083);
  and2 I040_019(w_040_019, w_009_512, w_013_124);
  and2 I040_021(w_040_021, w_024_193, w_001_024);
  nand2 I040_027(w_040_027, w_032_149, w_007_194);
  and2 I040_031(w_040_031, w_013_024, w_012_011);
  or2  I040_032(w_040_032, w_009_070, w_015_480);
  and2 I040_039(w_040_039, w_001_022, w_001_013);
  nand2 I040_040(w_040_040, w_038_000, w_002_005);
  and2 I040_043(w_040_043, w_021_202, w_027_059);
  or2  I040_044(w_040_044, w_018_012, w_025_114);
  or2  I040_045(w_040_045, w_001_006, w_021_074);
  nand2 I040_047(w_040_047, w_034_038, w_014_159);
  nand2 I040_049(w_040_049, w_022_001, w_001_024);
  or2  I040_050(w_040_050, w_023_189, w_036_262);
  and2 I040_051(w_040_051, w_015_103, w_001_004);
  not1 I040_053(w_040_053, w_008_342);
  or2  I040_054(w_040_054, w_002_692, w_011_088);
  or2  I040_063(w_040_063, w_038_542, w_033_161);
  or2  I040_065(w_040_065, w_001_022, w_029_070);
  or2  I040_067(w_040_067, w_020_160, w_032_174);
  and2 I040_068(w_040_068, w_017_612, w_004_191);
  and2 I040_070(w_040_070, w_039_372, w_017_186);
  or2  I040_071(w_040_071, w_030_312, w_026_371);
  and2 I040_072(w_040_072, w_011_027, w_003_079);
  or2  I040_077(w_040_077, w_010_322, w_031_273);
  not1 I040_080(w_040_080, w_001_019);
  nand2 I040_083(w_040_083, w_032_229, w_009_035);
  and2 I040_086(w_040_086, w_021_220, w_002_214);
  nand2 I040_088(w_040_088, w_009_230, w_002_000);
  and2 I040_090(w_040_090, w_008_202, w_032_124);
  nand2 I040_091(w_040_091, w_008_334, w_008_156);
  and2 I040_096(w_040_096, w_000_016, w_027_107);
  or2  I040_098(w_040_098, w_004_005, w_030_236);
  not1 I040_099(w_040_099, w_014_029);
  not1 I040_101(w_040_101, w_005_313);
  not1 I040_102(w_040_102, w_028_147);
  nand2 I040_106(w_040_106, w_035_112, w_020_029);
  and2 I040_119(w_040_119, w_001_020, w_009_344);
  nand2 I040_120(w_040_120, w_030_049, w_030_370);
  or2  I040_123(w_040_123, w_020_108, w_020_136);
  not1 I040_129(w_040_129, w_026_493);
  nand2 I040_132(w_040_132, w_030_276, w_032_175);
  not1 I040_133(w_040_133, w_018_037);
  and2 I040_139(w_040_139, w_022_309, w_014_108);
  nand2 I040_146(w_040_146, w_019_002, w_034_048);
  or2  I040_147(w_040_147, w_001_034, w_032_240);
  and2 I040_149(w_040_149, w_000_246, w_034_022);
  or2  I040_163(w_040_163, w_027_167, w_014_150);
  nand2 I040_164(w_040_164, w_018_019, w_038_157);
  or2  I040_166(w_040_166, w_002_030, w_002_006);
  not1 I040_174(w_040_174, w_036_232);
  not1 I040_180(w_040_180, w_033_330);
  and2 I040_184(w_040_184, w_037_249, w_034_068);
  and2 I040_193(w_040_193, w_034_009, w_037_060);
  not1 I040_196(w_040_196, w_036_131);
  not1 I040_210(w_040_210, w_027_044);
  and2 I040_219(w_040_219, w_016_001, w_019_015);
  or2  I040_221(w_040_221, w_004_257, w_010_441);
  or2  I040_225(w_040_225, w_039_141, w_033_123);
  or2  I040_228(w_040_228, w_020_475, w_039_373);
  or2  I040_234(w_040_234, w_024_034, w_013_412);
  and2 I040_235(w_040_235, w_025_130, w_015_119);
  or2  I040_238(w_040_238, w_024_017, w_002_655);
  or2  I040_241(w_040_241, w_034_040, w_005_133);
  or2  I040_243(w_040_243, w_030_278, w_010_736);
  and2 I040_246(w_040_246, w_007_053, w_015_348);
  and2 I040_252(w_040_252, w_005_025, w_023_101);
  and2 I040_254(w_040_254, w_019_011, w_004_047);
  or2  I040_257(w_040_257, w_014_202, w_010_191);
  not1 I040_268(w_040_268, w_029_027);
  not1 I040_278(w_040_278, w_017_056);
  and2 I040_281(w_040_281, w_000_624, w_017_017);
  or2  I040_283(w_040_283, w_034_065, w_030_228);
  not1 I040_286(w_040_286, w_033_510);
  not1 I040_288(w_040_288, w_003_034);
  and2 I040_294(w_040_294, w_032_294, w_027_064);
  and2 I040_295(w_040_295, w_030_099, w_036_393);
  and2 I040_298(w_040_298, w_025_048, w_021_168);
  and2 I040_299(w_040_299, w_024_059, w_032_414);
  or2  I040_304(w_040_304, w_037_001, w_009_032);
  or2  I040_309(w_040_309, w_002_576, w_019_018);
  nand2 I040_311(w_040_311, w_017_012, w_007_422);
  and2 I040_312(w_040_312, w_016_000, w_006_013);
  nand2 I040_316(w_040_316, w_016_004, w_003_073);
  nand2 I040_317(w_040_317, w_034_034, w_026_123);
  or2  I040_318(w_040_318, w_025_098, w_021_034);
  nand2 I040_322(w_040_322, w_039_278, w_028_162);
  and2 I040_324(w_040_324, w_005_193, w_033_551);
  not1 I040_325(w_040_325, w_006_079);
  not1 I040_327(w_040_327, w_023_084);
  not1 I040_328(w_040_328, w_022_297);
  or2  I040_340(w_040_340, w_028_361, w_017_343);
  or2  I040_343(w_040_343, w_010_242, w_030_083);
  and2 I040_346(w_040_346, w_023_092, w_037_120);
  and2 I040_348(w_040_348, w_020_297, w_017_426);
  and2 I040_353(w_040_353, w_007_428, w_030_080);
  not1 I040_356(w_040_356, w_028_499);
  not1 I040_357(w_040_357, w_017_403);
  not1 I040_358(w_040_358, w_037_169);
  or2  I040_360(w_040_360, w_025_054, w_005_178);
  not1 I040_361(w_040_361, w_033_015);
  or2  I040_366(w_040_366, w_013_104, w_010_155);
  or2  I040_367(w_040_367, w_035_082, w_010_164);
  or2  I040_371(w_040_371, w_027_146, w_033_391);
  not1 I040_373(w_040_373, w_025_101);
  nand2 I040_382(w_040_382, w_039_228, w_003_005);
  nand2 I040_386(w_040_386, w_005_226, w_014_105);
  or2  I040_393(w_040_393, w_024_010, w_016_002);
  or2  I040_395(w_040_395, w_036_011, w_017_495);
  not1 I040_404(w_040_404, w_007_428);
  and2 I040_405(w_040_405, w_013_357, w_034_053);
  not1 I040_409(w_040_409, w_018_004);
  or2  I040_415(w_040_415, w_034_059, w_038_103);
  nand2 I040_423(w_040_423, w_038_600, w_004_132);
  not1 I040_425(w_040_425, w_005_094);
  and2 I040_427(w_040_427, w_011_290, w_029_082);
  or2  I040_428(w_040_428, w_016_000, w_019_018);
  or2  I040_430(w_040_430, w_004_030, w_007_202);
  or2  I040_432(w_040_432, w_026_076, w_015_046);
  or2  I040_433(w_040_433, w_011_057, w_004_000);
  nand2 I040_439(w_040_439, w_021_083, w_024_184);
  and2 I040_440(w_040_440, w_028_184, w_027_078);
  and2 I040_441(w_040_441, w_020_010, w_035_064);
  or2  I040_442(w_040_442, w_033_698, w_029_008);
  or2  I040_449(w_040_449, w_013_140, w_020_615);
  and2 I040_462(w_040_462, w_036_447, w_028_057);
  not1 I040_463(w_040_463, w_015_548);
  or2  I040_464(w_040_464, w_031_065, w_001_012);
  not1 I040_468(w_040_468, w_028_512);
  nand2 I040_469(w_040_469, w_028_205, w_007_113);
  and2 I040_475(w_040_475, w_037_047, w_001_019);
  or2  I040_478(w_040_478, w_024_225, w_010_295);
  and2 I040_479(w_040_479, w_030_177, w_036_083);
  or2  I040_480(w_040_480, w_037_001, w_020_283);
  and2 I040_481(w_040_481, w_037_082, w_016_000);
  or2  I040_482(w_040_482, w_017_120, w_007_241);
  and2 I040_484(w_040_484, w_025_083, w_018_028);
  or2  I040_486(w_040_486, w_025_239, w_030_090);
  or2  I040_488(w_040_488, w_019_004, w_012_306);
  nand2 I040_493(w_040_493, w_007_166, w_031_490);
  or2  I040_497(w_040_497, w_034_030, w_018_015);
  nand2 I040_501(w_040_501, w_013_099, w_010_120);
  and2 I040_505(w_040_505, w_037_251, w_016_006);
  or2  I040_509(w_040_509, w_035_009, w_008_173);
  nand2 I040_514(w_040_514, w_024_120, w_013_029);
  nand2 I040_515(w_040_515, w_034_074, w_020_356);
  not1 I040_519(w_040_519, w_003_040);
  not1 I040_520(w_040_520, w_004_235);
  or2  I040_521(w_040_521, w_020_065, w_014_056);
  not1 I040_524(w_040_524, w_012_338);
  or2  I040_539(w_040_539, w_033_522, w_017_394);
  or2  I040_542(w_040_542, w_001_016, w_029_080);
  not1 I040_549(w_040_549, w_005_065);
  not1 I040_551(w_040_551, w_006_005);
  nand2 I040_553(w_040_553, w_005_242, w_002_596);
  and2 I040_554(w_040_554, w_021_193, w_038_397);
  and2 I040_555(w_040_555, w_039_524, w_005_113);
  or2  I040_558(w_040_558, w_005_033, w_007_172);
  nand2 I040_565(w_040_565, w_006_100, w_031_101);
  or2  I040_568(w_040_568, w_014_102, w_036_022);
  nand2 I040_571(w_040_571, w_003_006, w_000_716);
  or2  I040_582(w_040_582, w_033_335, w_003_015);
  nand2 I040_583(w_040_583, w_038_397, w_009_105);
  or2  I040_592(w_040_592, w_017_655, w_037_217);
  or2  I040_594(w_040_594, w_014_010, w_011_594);
  and2 I040_599(w_040_599, w_006_200, w_032_368);
  and2 I040_601(w_040_601, w_007_456, w_013_275);
  or2  I040_607(w_040_607, w_028_456, w_012_007);
  or2  I040_609(w_040_609, w_011_070, w_023_186);
  nand2 I040_611(w_040_611, w_008_147, w_027_181);
  nand2 I040_614(w_040_614, w_028_134, w_003_024);
  nand2 I040_616(w_040_616, w_007_091, w_025_261);
  not1 I040_617(w_040_617, w_032_509);
  nand2 I040_623(w_040_623, w_008_545, w_019_020);
  nand2 I040_630(w_040_630, w_036_064, w_030_201);
  not1 I040_632(w_040_632, w_015_426);
  or2  I040_639(w_040_639, w_021_204, w_029_048);
  or2  I040_644(w_040_644, w_025_108, w_026_188);
  not1 I040_646(w_040_646, w_035_076);
  and2 I040_660(w_040_660, w_026_055, w_008_312);
  and2 I040_663(w_040_663, w_027_114, w_018_023);
  nand2 I040_667(w_040_667, w_036_305, w_032_025);
  nand2 I040_670(w_040_670, w_002_017, w_034_016);
  and2 I040_682(w_040_682, w_011_435, w_007_296);
  not1 I040_689(w_040_689, w_039_306);
  and2 I040_691(w_040_691, w_026_430, w_007_028);
  not1 I040_692(w_040_692, w_029_083);
  not1 I040_693(w_040_693, w_015_069);
  or2  I040_698(w_040_698, w_004_225, w_039_466);
  and2 I040_699(w_040_699, w_029_044, w_013_132);
  not1 I040_704(w_040_704, w_037_158);
  nand2 I040_705(w_040_705, w_033_735, w_002_019);
  not1 I040_713(w_040_713, w_005_083);
  nand2 I040_718(w_040_720, w_040_719, w_019_001);
  not1 I040_719(w_040_721, w_040_720);
  not1 I040_720(w_040_722, w_040_721);
  and2 I040_721(w_040_723, w_014_243, w_040_722);
  and2 I040_722(w_040_724, w_030_226, w_040_723);
  not1 I040_723(w_040_725, w_040_724);
  not1 I040_724(w_040_726, w_040_725);
  nand2 I040_725(w_040_727, w_017_048, w_040_726);
  nand2 I040_726(w_040_728, w_006_137, w_040_727);
  nand2 I040_727(w_040_729, w_008_659, w_040_728);
  and2 I040_728(w_040_730, w_040_729, w_033_336);
  nand2 I040_729(w_040_719, w_040_730, w_006_160);
  not1 I041_007(w_041_007, w_028_354);
  nand2 I041_010(w_041_010, w_017_609, w_039_214);
  or2  I041_011(w_041_011, w_008_015, w_018_033);
  and2 I041_013(w_041_013, w_017_007, w_019_016);
  nand2 I041_016(w_041_016, w_024_300, w_023_106);
  not1 I041_023(w_041_023, w_019_017);
  nand2 I041_024(w_041_024, w_035_052, w_019_016);
  nand2 I041_026(w_041_026, w_004_446, w_015_060);
  nand2 I041_029(w_041_029, w_018_043, w_018_044);
  or2  I041_032(w_041_032, w_038_019, w_025_241);
  not1 I041_035(w_041_035, w_036_153);
  or2  I041_036(w_041_036, w_015_286, w_035_110);
  nand2 I041_037(w_041_037, w_008_211, w_030_106);
  nand2 I041_038(w_041_038, w_031_086, w_039_478);
  not1 I041_041(w_041_041, w_009_510);
  or2  I041_046(w_041_046, w_020_450, w_013_548);
  nand2 I041_048(w_041_048, w_027_094, w_005_015);
  or2  I041_051(w_041_051, w_004_123, w_012_000);
  nand2 I041_052(w_041_052, w_015_105, w_037_034);
  or2  I041_053(w_041_053, w_000_437, w_008_278);
  not1 I041_054(w_041_054, w_012_350);
  nand2 I041_055(w_041_055, w_019_012, w_027_039);
  and2 I041_057(w_041_057, w_020_205, w_026_333);
  or2  I041_060(w_041_060, w_037_050, w_024_057);
  not1 I041_062(w_041_062, w_012_346);
  or2  I041_070(w_041_070, w_005_114, w_014_097);
  or2  I041_073(w_041_073, w_001_024, w_038_333);
  not1 I041_077(w_041_077, w_025_124);
  or2  I041_079(w_041_079, w_015_660, w_018_011);
  nand2 I041_081(w_041_081, w_022_252, w_014_068);
  and2 I041_083(w_041_083, w_003_042, w_032_000);
  nand2 I041_086(w_041_086, w_025_105, w_005_047);
  not1 I041_088(w_041_088, w_000_676);
  or2  I041_090(w_041_090, w_000_403, w_000_250);
  nand2 I041_097(w_041_097, w_035_069, w_028_203);
  not1 I041_100(w_041_100, w_030_107);
  not1 I041_102(w_041_102, w_035_114);
  nand2 I041_104(w_041_104, w_033_251, w_002_634);
  and2 I041_106(w_041_106, w_021_091, w_028_090);
  nand2 I041_110(w_041_110, w_016_004, w_020_181);
  not1 I041_113(w_041_113, w_010_282);
  and2 I041_116(w_041_116, w_030_144, w_033_452);
  nand2 I041_117(w_041_117, w_009_098, w_007_222);
  and2 I041_128(w_041_128, w_014_153, w_026_393);
  nand2 I041_131(w_041_131, w_029_060, w_011_310);
  not1 I041_138(w_041_138, w_012_286);
  not1 I041_154(w_041_154, w_005_139);
  and2 I041_160(w_041_160, w_038_575, w_001_030);
  nand2 I041_166(w_041_166, w_019_011, w_037_228);
  and2 I041_172(w_041_172, w_038_052, w_038_064);
  and2 I041_178(w_041_178, w_003_003, w_001_030);
  nand2 I041_181(w_041_181, w_014_127, w_037_339);
  not1 I041_185(w_041_185, w_028_366);
  nand2 I041_189(w_041_189, w_014_245, w_031_231);
  and2 I041_194(w_041_194, w_020_297, w_032_077);
  not1 I041_197(w_041_197, w_026_093);
  nand2 I041_206(w_041_206, w_040_184, w_031_593);
  not1 I041_212(w_041_212, w_011_026);
  nand2 I041_220(w_041_220, w_015_271, w_035_044);
  or2  I041_226(w_041_226, w_006_232, w_013_199);
  or2  I041_228(w_041_228, w_032_599, w_032_433);
  nand2 I041_231(w_041_231, w_015_091, w_017_406);
  nand2 I041_234(w_041_234, w_012_299, w_015_205);
  not1 I041_241(w_041_241, w_029_086);
  nand2 I041_243(w_041_243, w_028_154, w_028_052);
  or2  I041_244(w_041_244, w_028_262, w_019_010);
  or2  I041_246(w_041_246, w_032_193, w_002_453);
  nand2 I041_248(w_041_248, w_000_531, w_014_193);
  or2  I041_257(w_041_257, w_017_356, w_012_229);
  or2  I041_263(w_041_263, w_036_019, w_017_492);
  or2  I041_275(w_041_275, w_019_000, w_010_759);
  or2  I041_276(w_041_276, w_033_558, w_040_632);
  not1 I041_279(w_041_279, w_034_026);
  and2 I041_282(w_041_282, w_031_126, w_000_743);
  nand2 I041_288(w_041_288, w_024_146, w_016_000);
  not1 I041_293(w_041_293, w_030_242);
  and2 I041_298(w_041_298, w_017_010, w_009_249);
  nand2 I041_300(w_041_300, w_005_113, w_023_153);
  and2 I041_304(w_041_304, w_007_478, w_024_125);
  not1 I041_305(w_041_305, w_002_135);
  or2  I041_306(w_041_306, w_021_127, w_027_149);
  nand2 I041_315(w_041_315, w_003_046, w_027_175);
  not1 I041_326(w_041_326, w_009_150);
  nand2 I041_334(w_041_334, w_023_212, w_026_122);
  not1 I041_336(w_041_336, w_008_149);
  and2 I041_337(w_041_337, w_012_090, w_033_382);
  not1 I041_338(w_041_338, w_024_312);
  and2 I041_339(w_041_339, w_017_066, w_013_259);
  not1 I041_340(w_041_340, w_036_151);
  not1 I041_342(w_041_342, w_005_135);
  not1 I041_345(w_041_345, w_012_203);
  and2 I041_346(w_041_346, w_038_383, w_024_119);
  not1 I041_349(w_041_349, w_016_005);
  or2  I041_354(w_041_354, w_040_322, w_028_170);
  not1 I041_355(w_041_355, w_040_133);
  not1 I041_359(w_041_359, w_000_543);
  not1 I041_378(w_041_378, w_024_388);
  or2  I041_380(w_041_380, w_001_013, w_010_108);
  not1 I041_389(w_041_389, w_015_502);
  not1 I041_392(w_041_392, w_010_058);
  or2  I041_397(w_041_397, w_016_001, w_030_414);
  or2  I041_399(w_041_399, w_029_091, w_008_487);
  not1 I041_403(w_041_403, w_004_427);
  or2  I041_408(w_041_408, w_022_126, w_027_009);
  and2 I041_409(w_041_409, w_031_223, w_017_010);
  not1 I041_412(w_041_412, w_021_222);
  and2 I041_414(w_041_414, w_029_078, w_016_000);
  and2 I041_429(w_041_429, w_019_018, w_023_100);
  nand2 I041_432(w_041_432, w_001_031, w_033_487);
  not1 I041_433(w_041_433, w_000_351);
  or2  I041_434(w_041_434, w_028_522, w_005_058);
  or2  I041_439(w_041_439, w_012_350, w_001_029);
  or2  I041_441(w_041_441, w_021_194, w_039_327);
  or2  I041_444(w_041_444, w_005_251, w_034_069);
  not1 I041_446(w_041_446, w_012_282);
  and2 I041_453(w_041_453, w_025_039, w_022_036);
  or2  I041_457(w_041_457, w_024_195, w_039_219);
  or2  I041_460(w_041_460, w_036_324, w_024_105);
  and2 I041_463(w_041_463, w_014_055, w_039_348);
  nand2 I041_476(w_041_476, w_010_765, w_008_710);
  or2  I041_482(w_041_482, w_021_240, w_018_037);
  or2  I041_485(w_041_485, w_001_010, w_040_609);
  nand2 I041_488(w_041_488, w_040_304, w_021_105);
  or2  I041_489(w_041_489, w_003_002, w_027_091);
  and2 I041_491(w_041_491, w_018_006, w_003_049);
  or2  I041_494(w_041_494, w_002_227, w_040_040);
  and2 I041_496(w_041_496, w_002_515, w_007_127);
  and2 I041_497(w_041_497, w_029_109, w_004_162);
  not1 I041_499(w_041_499, w_006_039);
  or2  I041_504(w_041_504, w_007_112, w_025_141);
  or2  I041_507(w_041_507, w_014_017, w_032_037);
  not1 I041_510(w_041_510, w_020_416);
  nand2 I041_511(w_041_511, w_029_056, w_019_004);
  or2  I041_512(w_041_512, w_010_520, w_014_261);
  not1 I041_513(w_041_513, w_011_385);
  or2  I041_515(w_041_515, w_031_265, w_014_047);
  or2  I041_524(w_041_524, w_024_036, w_022_185);
  not1 I041_525(w_041_525, w_027_041);
  or2  I041_528(w_041_528, w_038_211, w_040_243);
  or2  I041_529(w_041_529, w_012_019, w_005_114);
  and2 I041_531(w_041_531, w_014_259, w_039_561);
  or2  I041_532(w_041_532, w_000_289, w_005_123);
  or2  I041_535(w_041_535, w_031_069, w_024_346);
  or2  I041_537(w_041_537, w_027_070, w_008_602);
  and2 I041_541(w_041_541, w_040_462, w_032_451);
  or2  I041_548(w_041_548, w_032_060, w_013_015);
  nand2 I041_549(w_041_549, w_032_153, w_029_050);
  not1 I041_561(w_041_561, w_013_079);
  nand2 I041_576(w_041_576, w_023_123, w_005_005);
  not1 I041_579(w_041_579, w_009_370);
  not1 I041_581(w_041_581, w_025_283);
  and2 I041_583(w_041_583, w_019_012, w_036_284);
  not1 I041_587(w_041_587, w_029_022);
  nand2 I041_589(w_041_589, w_037_218, w_026_211);
  not1 I041_593(w_041_593, w_022_011);
  not1 I041_594(w_041_594, w_026_381);
  not1 I041_604(w_041_604, w_039_061);
  or2  I041_606(w_041_606, w_004_265, w_023_023);
  and2 I041_610(w_041_610, w_038_431, w_011_046);
  nand2 I041_614(w_041_614, w_036_430, w_027_097);
  and2 I041_618(w_041_618, w_026_149, w_022_360);
  or2  I041_623(w_041_623, w_000_735, w_003_029);
  or2  I041_625(w_041_625, w_034_027, w_036_432);
  or2  I041_627(w_041_627, w_016_001, w_034_060);
  or2  I041_628(w_041_628, w_024_421, w_027_002);
  or2  I041_630(w_041_630, w_006_068, w_005_112);
  and2 I041_632(w_041_632, w_013_117, w_020_078);
  and2 I041_647(w_041_647, w_019_008, w_024_355);
  nand2 I041_659(w_041_659, w_021_194, w_023_105);
  and2 I041_661(w_041_661, w_039_078, w_023_181);
  and2 I041_663(w_041_663, w_016_007, w_016_006);
  and2 I041_664(w_041_664, w_011_457, w_026_695);
  not1 I041_665(w_041_665, w_013_256);
  nand2 I041_668(w_041_668, w_004_499, w_031_154);
  or2  I041_670(w_041_670, w_035_030, w_003_044);
  or2  I041_673(w_041_673, w_036_164, w_030_355);
  and2 I041_676(w_041_676, w_002_091, w_019_000);
  or2  I041_683(w_041_683, w_010_303, w_008_685);
  not1 I041_685(w_041_685, w_031_153);
  or2  I041_692(w_041_692, w_030_205, w_020_084);
  or2  I041_698(w_041_698, w_036_359, w_025_018);
  nand2 I041_713(w_041_713, w_012_198, w_020_067);
  nand2 I041_714(w_041_714, w_030_309, w_007_092);
  not1 I041_721(w_041_721, w_024_307);
  and2 I042_000(w_042_000, w_029_068, w_015_071);
  not1 I042_001(w_042_001, w_035_047);
  not1 I042_002(w_042_002, w_034_026);
  or2  I042_005(w_042_005, w_011_359, w_012_038);
  nand2 I042_006(w_042_006, w_021_036, w_011_030);
  nand2 I042_008(w_042_008, w_008_035, w_003_067);
  nand2 I042_010(w_042_010, w_026_675, w_014_294);
  and2 I042_012(w_042_012, w_041_097, w_034_052);
  not1 I042_013(w_042_013, w_025_155);
  or2  I042_018(w_042_018, w_037_150, w_039_530);
  nand2 I042_023(w_042_023, w_021_042, w_025_141);
  or2  I042_024(w_042_024, w_002_022, w_039_037);
  and2 I042_025(w_042_025, w_007_001, w_003_066);
  and2 I042_026(w_042_026, w_003_047, w_006_132);
  not1 I042_034(w_042_034, w_035_099);
  not1 I042_035(w_042_035, w_000_770);
  and2 I042_036(w_042_036, w_035_078, w_015_677);
  not1 I042_038(w_042_038, w_013_229);
  not1 I042_039(w_042_039, w_012_115);
  not1 I042_041(w_042_041, w_011_315);
  or2  I042_043(w_042_043, w_006_192, w_003_055);
  not1 I042_044(w_042_044, w_038_047);
  nand2 I042_045(w_042_045, w_008_283, w_011_110);
  not1 I042_050(w_042_050, w_020_059);
  and2 I042_052(w_042_052, w_033_406, w_033_587);
  or2  I042_056(w_042_056, w_009_396, w_013_174);
  not1 I042_057(w_042_057, w_033_369);
  not1 I042_059(w_042_059, w_007_235);
  nand2 I042_061(w_042_061, w_011_120, w_003_021);
  and2 I042_062(w_042_062, w_002_094, w_026_488);
  and2 I042_066(w_042_066, w_008_295, w_032_497);
  and2 I042_071(w_042_071, w_003_078, w_037_320);
  nand2 I042_072(w_042_072, w_020_057, w_038_462);
  nand2 I042_076(w_042_076, w_023_112, w_039_620);
  or2  I042_077(w_042_077, w_037_210, w_026_039);
  or2  I042_081(w_042_081, w_025_066, w_002_276);
  nand2 I042_082(w_042_082, w_041_392, w_032_158);
  not1 I042_084(w_042_084, w_014_163);
  not1 I042_090(w_042_090, w_037_229);
  and2 I042_092(w_042_092, w_007_099, w_010_476);
  nand2 I042_094(w_042_094, w_038_079, w_015_344);
  nand2 I042_095(w_042_095, w_032_465, w_013_373);
  or2  I042_099(w_042_099, w_000_714, w_009_027);
  and2 I042_101(w_042_101, w_023_110, w_019_017);
  nand2 I042_102(w_042_102, w_032_060, w_041_345);
  or2  I042_103(w_042_103, w_033_451, w_031_370);
  nand2 I042_104(w_042_104, w_000_292, w_015_019);
  nand2 I042_109(w_042_109, w_003_032, w_035_069);
  or2  I042_110(w_042_110, w_000_054, w_016_001);
  not1 I042_111(w_042_111, w_031_465);
  and2 I042_112(w_042_112, w_037_010, w_035_052);
  and2 I042_113(w_042_113, w_004_143, w_002_421);
  nand2 I042_116(w_042_116, w_017_594, w_013_399);
  and2 I042_117(w_042_117, w_029_032, w_018_027);
  nand2 I042_121(w_042_121, w_023_120, w_004_349);
  and2 I042_123(w_042_123, w_020_076, w_016_008);
  and2 I042_124(w_042_124, w_033_396, w_022_026);
  not1 I042_125(w_042_125, w_011_594);
  and2 I042_126(w_042_126, w_015_669, w_039_404);
  or2  I042_127(w_042_127, w_011_054, w_022_080);
  not1 I042_130(w_042_130, w_009_365);
  not1 I042_132(w_042_132, w_008_709);
  nand2 I042_133(w_042_133, w_030_308, w_039_072);
  or2  I042_134(w_042_134, w_000_239, w_011_309);
  nand2 I042_135(w_042_135, w_008_449, w_039_052);
  nand2 I042_138(w_042_138, w_026_038, w_011_132);
  or2  I042_139(w_042_139, w_019_020, w_036_269);
  or2  I042_144(w_042_144, w_015_333, w_013_323);
  and2 I042_146(w_042_146, w_034_060, w_034_010);
  and2 I042_147(w_042_147, w_025_171, w_018_023);
  not1 I042_148(w_042_148, w_022_031);
  and2 I042_150(w_042_150, w_028_206, w_014_286);
  or2  I042_152(w_042_152, w_011_510, w_017_495);
  not1 I042_155(w_042_155, w_015_229);
  or2  I042_156(w_042_156, w_004_438, w_029_001);
  and2 I042_157(w_042_157, w_026_549, w_004_184);
  nand2 I042_158(w_042_158, w_004_275, w_008_232);
  nand2 I042_159(w_042_159, w_015_346, w_036_227);
  and2 I042_162(w_042_162, w_003_075, w_021_233);
  and2 I042_165(w_042_165, w_006_185, w_022_117);
  and2 I042_169(w_042_169, w_028_393, w_036_049);
  or2  I042_171(w_042_171, w_034_013, w_012_252);
  or2  I042_172(w_042_172, w_007_035, w_022_144);
  and2 I042_178(w_042_178, w_034_034, w_009_594);
  not1 I042_180(w_042_180, w_007_213);
  nand2 I042_181(w_042_181, w_018_018, w_004_288);
  nand2 I042_182(w_042_182, w_004_173, w_031_444);
  not1 I042_184(w_042_184, w_001_008);
  not1 I042_185(w_042_185, w_009_000);
  nand2 I042_186(w_042_186, w_027_143, w_019_005);
  and2 I042_191(w_042_191, w_004_284, w_023_011);
  not1 I042_192(w_042_192, w_002_094);
  and2 I042_194(w_042_194, w_041_683, w_017_027);
  nand2 I042_195(w_042_195, w_005_101, w_040_068);
  nand2 I042_197(w_042_197, w_029_035, w_001_007);
  and2 I042_198(w_042_198, w_024_096, w_010_384);
  nand2 I042_199(w_042_199, w_020_003, w_027_001);
  or2  I042_201(w_042_201, w_028_147, w_002_500);
  nand2 I042_203(w_042_203, w_013_035, w_006_197);
  or2  I042_206(w_042_206, w_033_095, w_031_602);
  and2 I042_209(w_042_209, w_026_648, w_023_074);
  not1 I042_215(w_042_215, w_034_018);
  not1 I042_217(w_042_217, w_014_044);
  not1 I042_219(w_042_219, w_026_305);
  not1 I042_220(w_042_220, w_004_354);
  nand2 I042_222(w_042_222, w_000_436, w_037_013);
  nand2 I042_226(w_042_226, w_028_425, w_035_000);
  nand2 I042_227(w_042_227, w_040_482, w_024_506);
  or2  I042_229(w_042_229, w_031_175, w_019_001);
  or2  I042_232(w_042_232, w_021_177, w_008_021);
  and2 I042_233(w_042_233, w_002_115, w_040_440);
  or2  I042_237(w_042_237, w_018_036, w_014_129);
  nand2 I042_252(w_042_252, w_012_203, w_005_022);
  and2 I042_255(w_042_255, w_027_014, w_013_471);
  nand2 I042_257(w_042_257, w_011_460, w_011_548);
  nand2 I042_258(w_042_258, w_039_581, w_003_053);
  and2 I042_260(w_042_260, w_007_139, w_021_244);
  and2 I042_261(w_042_261, w_007_015, w_022_195);
  or2  I042_264(w_042_264, w_035_039, w_035_025);
  or2  I042_265(w_042_265, w_036_461, w_038_598);
  not1 I042_267(w_042_267, w_010_737);
  nand2 I042_268(w_042_268, w_006_105, w_027_155);
  or2  I042_271(w_042_271, w_032_330, w_016_004);
  nand2 I042_272(w_042_272, w_008_726, w_013_552);
  and2 I042_275(w_042_275, w_013_534, w_010_766);
  or2  I042_276(w_042_276, w_025_019, w_011_025);
  not1 I042_278(w_042_278, w_018_017);
  and2 I042_279(w_042_279, w_030_040, w_038_588);
  not1 I042_281(w_042_281, w_004_126);
  not1 I042_282(w_042_282, w_000_643);
  and2 I042_286(w_042_286, w_022_012, w_020_342);
  not1 I042_288(w_042_288, w_033_059);
  or2  I042_290(w_042_290, w_033_119, w_038_079);
  nand2 I042_292(w_042_292, w_017_020, w_008_089);
  or2  I042_293(w_042_293, w_028_512, w_019_009);
  or2  I042_295(w_042_295, w_036_129, w_014_049);
  not1 I042_297(w_042_297, w_019_008);
  and2 I042_298(w_042_298, w_019_004, w_033_510);
  and2 I042_304(w_042_304, w_003_068, w_030_185);
  not1 I042_305(w_042_305, w_020_058);
  not1 I042_307(w_042_307, w_003_032);
  nand2 I042_309(w_042_309, w_012_006, w_004_022);
  or2  I042_310(w_042_310, w_028_324, w_005_195);
  or2  I042_311(w_042_311, w_006_246, w_033_608);
  nand2 I042_312(w_042_312, w_009_482, w_000_051);
  not1 I042_316(w_042_316, w_009_402);
  nand2 I042_317(w_042_317, w_037_279, w_018_026);
  and2 I042_318(w_042_318, w_022_160, w_009_238);
  nand2 I042_319(w_042_319, w_017_272, w_016_005);
  or2  I042_320(w_042_320, w_022_282, w_003_053);
  and2 I042_321(w_042_321, w_036_094, w_027_056);
  nand2 I042_323(w_042_323, w_011_152, w_036_311);
  nand2 I042_325(w_042_325, w_010_678, w_016_003);
  nand2 I042_327(w_042_327, w_023_114, w_014_050);
  and2 I042_328(w_042_328, w_018_020, w_039_221);
  nand2 I042_331(w_042_331, w_007_137, w_029_008);
  not1 I042_332(w_042_332, w_003_076);
  nand2 I042_334(w_042_334, w_033_216, w_012_183);
  or2  I042_339(w_042_339, w_014_224, w_034_035);
  nand2 I042_340(w_042_340, w_028_037, w_026_499);
  not1 I042_343(w_042_343, w_021_212);
  not1 I042_346(w_042_346, w_006_160);
  nand2 I042_356(w_042_356, w_016_003, w_028_001);
  nand2 I042_358(w_042_358, w_011_072, w_022_287);
  or2  I042_359(w_042_359, w_031_520, w_038_315);
  or2  I042_362(w_042_362, w_002_441, w_032_508);
  not1 I042_367(w_042_367, w_036_182);
  and2 I042_368(w_042_368, w_010_230, w_041_618);
  nand2 I042_369(w_042_369, w_030_252, w_005_252);
  nand2 I042_377(w_042_377, w_035_024, w_011_140);
  not1 I042_384(w_042_384, w_028_479);
  nand2 I042_385(w_042_385, w_041_336, w_030_194);
  and2 I042_389(w_042_389, w_027_170, w_013_060);
  nand2 I042_401(w_042_401, w_033_580, w_003_031);
  not1 I042_402(w_042_402, w_008_182);
  nand2 I042_404(w_042_404, w_037_149, w_037_020);
  and2 I042_406(w_042_406, w_002_695, w_010_618);
  nand2 I042_409(w_042_409, w_028_567, w_014_047);
  nand2 I042_413(w_042_413, w_017_123, w_017_336);
  and2 I042_414(w_042_414, w_026_028, w_041_632);
  and2 I042_415(w_042_415, w_020_217, w_015_112);
  nand2 I042_422(w_042_422, w_041_029, w_022_264);
  or2  I042_423(w_042_423, w_008_561, w_001_032);
  or2  I042_427(w_042_427, w_015_172, w_037_131);
  and2 I042_428(w_042_428, w_000_010, w_041_293);
  nand2 I042_432(w_042_432, w_039_544, w_037_071);
  or2  I042_433(w_042_433, w_020_058, w_006_080);
  nand2 I042_437(w_042_437, w_026_572, w_026_361);
  not1 I042_443(w_042_443, w_001_020);
  or2  I042_451(w_042_451, w_029_016, w_035_094);
  or2  I042_453(w_042_453, w_018_044, w_028_408);
  and2 I042_455(w_042_455, w_025_132, w_021_264);
  or2  I042_456(w_042_456, w_036_357, w_013_054);
  or2  I043_000(w_043_000, w_006_034, w_030_073);
  not1 I043_001(w_043_001, w_039_606);
  and2 I043_002(w_043_002, w_032_089, w_015_277);
  nand2 I043_003(w_043_003, w_038_054, w_025_174);
  not1 I043_004(w_043_004, w_014_243);
  nand2 I043_005(w_043_005, w_032_261, w_019_005);
  and2 I043_006(w_043_006, w_042_307, w_026_107);
  or2  I043_007(w_043_007, w_032_046, w_015_290);
  not1 I043_008(w_043_008, w_003_011);
  not1 I043_009(w_043_009, w_027_134);
  not1 I043_010(w_043_010, w_025_075);
  not1 I043_011(w_043_011, w_023_029);
  or2  I043_012(w_043_012, w_003_028, w_029_062);
  not1 I043_013(w_043_013, w_035_124);
  not1 I043_014(w_043_014, w_019_005);
  not1 I043_015(w_043_015, w_002_596);
  and2 I043_016(w_043_016, w_034_064, w_030_222);
  not1 I043_017(w_043_017, w_033_297);
  and2 I043_018(w_043_018, w_018_008, w_027_093);
  nand2 I043_019(w_043_019, w_012_282, w_002_601);
  nand2 I043_020(w_043_020, w_038_415, w_032_377);
  not1 I043_021(w_043_021, w_029_097);
  or2  I043_022(w_043_022, w_025_042, w_023_028);
  not1 I043_023(w_043_023, w_014_024);
  and2 I043_024(w_043_024, w_009_338, w_042_010);
  not1 I043_025(w_043_025, w_017_207);
  and2 I043_026(w_043_026, w_002_023, w_003_073);
  or2  I043_027(w_043_027, w_035_066, w_019_005);
  not1 I043_028(w_043_028, w_023_065);
  not1 I043_029(w_043_029, w_042_199);
  nand2 I043_030(w_043_030, w_006_208, w_009_469);
  nand2 I043_031(w_043_031, w_009_035, w_028_310);
  and2 I043_032(w_043_032, w_032_041, w_011_084);
  or2  I043_033(w_043_033, w_005_112, w_033_194);
  and2 I043_034(w_043_034, w_025_069, w_001_036);
  nand2 I043_035(w_043_035, w_024_492, w_031_420);
  and2 I043_036(w_043_036, w_021_003, w_034_016);
  or2  I043_037(w_043_037, w_010_368, w_002_646);
  nand2 I043_038(w_043_038, w_039_718, w_030_113);
  or2  I043_039(w_043_039, w_024_064, w_006_071);
  nand2 I043_040(w_043_040, w_031_415, w_026_532);
  and2 I043_041(w_043_041, w_033_515, w_038_150);
  nand2 I043_042(w_043_042, w_016_002, w_028_042);
  nand2 I043_043(w_043_043, w_028_187, w_002_406);
  or2  I043_044(w_043_044, w_029_056, w_015_116);
  or2  I043_045(w_043_045, w_013_104, w_033_201);
  nand2 I043_046(w_043_046, w_003_057, w_028_301);
  or2  I043_047(w_043_047, w_027_121, w_013_348);
  nand2 I044_000(w_044_000, w_036_126, w_026_523);
  and2 I044_002(w_044_002, w_013_564, w_007_294);
  or2  I044_013(w_044_013, w_016_006, w_038_504);
  not1 I044_014(w_044_014, w_002_503);
  not1 I044_019(w_044_019, w_015_120);
  or2  I044_021(w_044_021, w_028_140, w_030_411);
  nand2 I044_022(w_044_022, w_018_036, w_036_318);
  not1 I044_026(w_044_026, w_039_580);
  or2  I044_027(w_044_027, w_021_004, w_010_042);
  not1 I044_029(w_044_029, w_039_063);
  or2  I044_030(w_044_030, w_024_035, w_039_158);
  not1 I044_033(w_044_033, w_033_238);
  not1 I044_036(w_044_036, w_023_005);
  nand2 I044_040(w_044_040, w_031_367, w_004_053);
  nand2 I044_041(w_044_041, w_035_008, w_024_319);
  nand2 I044_046(w_044_046, w_039_612, w_038_455);
  and2 I044_048(w_044_048, w_015_087, w_031_509);
  nand2 I044_050(w_044_050, w_005_301, w_036_283);
  not1 I044_054(w_044_054, w_007_025);
  and2 I044_055(w_044_055, w_017_063, w_007_077);
  and2 I044_058(w_044_058, w_005_067, w_037_189);
  not1 I044_062(w_044_062, w_028_120);
  not1 I044_070(w_044_070, w_023_084);
  nand2 I044_072(w_044_072, w_016_007, w_034_064);
  and2 I044_080(w_044_080, w_009_310, w_001_023);
  not1 I044_082(w_044_082, w_042_102);
  or2  I044_093(w_044_093, w_029_047, w_006_014);
  or2  I044_098(w_044_098, w_033_719, w_037_074);
  or2  I044_100(w_044_100, w_006_220, w_019_007);
  nand2 I044_109(w_044_109, w_005_028, w_031_171);
  and2 I044_110(w_044_110, w_040_366, w_017_006);
  or2  I044_115(w_044_115, w_013_076, w_032_478);
  nand2 I044_119(w_044_119, w_041_116, w_007_188);
  nand2 I044_122(w_044_122, w_003_058, w_023_108);
  or2  I044_127(w_044_127, w_021_111, w_005_042);
  and2 I044_128(w_044_128, w_015_333, w_027_146);
  and2 I044_137(w_044_137, w_026_189, w_023_088);
  nand2 I044_139(w_044_139, w_022_048, w_017_421);
  not1 I044_154(w_044_154, w_036_310);
  and2 I044_158(w_044_158, w_013_166, w_043_009);
  not1 I044_159(w_044_159, w_023_115);
  or2  I044_160(w_044_160, w_022_010, w_035_003);
  not1 I044_165(w_044_165, w_041_713);
  and2 I044_169(w_044_169, w_019_001, w_023_003);
  or2  I044_175(w_044_175, w_004_344, w_003_063);
  and2 I044_180(w_044_180, w_013_103, w_000_337);
  and2 I044_181(w_044_181, w_010_051, w_017_114);
  nand2 I044_191(w_044_191, w_029_087, w_002_317);
  not1 I044_195(w_044_195, w_016_003);
  and2 I044_197(w_044_197, w_030_177, w_023_117);
  not1 I044_199(w_044_199, w_018_005);
  not1 I044_201(w_044_201, w_006_074);
  or2  I044_206(w_044_206, w_032_011, w_011_405);
  not1 I044_209(w_044_209, w_041_100);
  and2 I044_219(w_044_219, w_022_165, w_000_044);
  and2 I044_223(w_044_223, w_001_009, w_011_089);
  or2  I044_225(w_044_225, w_008_117, w_010_406);
  and2 I044_229(w_044_229, w_024_210, w_008_473);
  nand2 I044_243(w_044_243, w_037_063, w_029_096);
  or2  I044_248(w_044_248, w_039_599, w_019_015);
  not1 I044_261(w_044_261, w_028_160);
  and2 I044_267(w_044_267, w_009_393, w_004_294);
  and2 I044_268(w_044_268, w_017_288, w_036_278);
  nand2 I044_273(w_044_273, w_000_526, w_025_182);
  not1 I044_276(w_044_276, w_001_013);
  or2  I044_284(w_044_284, w_005_090, w_035_060);
  nand2 I044_286(w_044_286, w_003_079, w_037_303);
  not1 I044_289(w_044_289, w_043_036);
  nand2 I044_290(w_044_290, w_031_160, w_036_273);
  and2 I044_292(w_044_292, w_042_084, w_003_025);
  and2 I044_293(w_044_293, w_040_328, w_027_112);
  or2  I044_295(w_044_295, w_023_048, w_043_035);
  and2 I044_296(w_044_296, w_034_018, w_029_031);
  nand2 I044_301(w_044_301, w_009_078, w_000_364);
  nand2 I044_303(w_044_303, w_030_199, w_000_461);
  nand2 I044_306(w_044_306, w_043_001, w_028_038);
  or2  I044_312(w_044_312, w_010_716, w_016_001);
  or2  I044_322(w_044_322, w_025_009, w_034_036);
  not1 I044_331(w_044_331, w_010_579);
  or2  I044_332(w_044_332, w_020_498, w_009_033);
  nand2 I044_335(w_044_335, w_016_004, w_011_173);
  not1 I044_338(w_044_338, w_035_066);
  not1 I044_341(w_044_341, w_043_041);
  and2 I044_344(w_044_344, w_031_148, w_010_359);
  and2 I044_347(w_044_347, w_032_225, w_042_023);
  nand2 I044_348(w_044_348, w_017_249, w_025_036);
  not1 I044_366(w_044_366, w_018_016);
  not1 I044_367(w_044_367, w_014_132);
  or2  I044_371(w_044_371, w_024_563, w_003_015);
  not1 I044_373(w_044_373, w_003_061);
  not1 I044_375(w_044_375, w_006_071);
  nand2 I044_377(w_044_377, w_021_155, w_002_592);
  or2  I044_384(w_044_384, w_004_125, w_012_013);
  not1 I044_390(w_044_390, w_036_078);
  not1 I044_395(w_044_395, w_035_003);
  not1 I044_398(w_044_398, w_014_134);
  not1 I044_402(w_044_402, w_032_430);
  not1 I044_403(w_044_403, w_016_004);
  and2 I044_405(w_044_405, w_003_065, w_017_569);
  nand2 I044_407(w_044_407, w_009_302, w_016_003);
  or2  I044_414(w_044_414, w_035_005, w_003_084);
  and2 I044_418(w_044_418, w_037_083, w_000_772);
  and2 I044_419(w_044_419, w_038_152, w_012_108);
  and2 I044_424(w_044_424, w_013_257, w_016_006);
  nand2 I044_435(w_044_435, w_008_693, w_010_443);
  not1 I044_447(w_044_447, w_025_167);
  or2  I044_449(w_044_449, w_032_553, w_024_180);
  or2  I044_450(w_044_450, w_019_008, w_006_106);
  or2  I044_452(w_044_452, w_007_021, w_034_032);
  not1 I044_454(w_044_454, w_039_208);
  or2  I044_457(w_044_457, w_043_003, w_039_072);
  or2  I044_458(w_044_458, w_005_282, w_038_160);
  not1 I044_459(w_044_459, w_004_496);
  nand2 I044_460(w_044_460, w_023_104, w_014_094);
  and2 I044_461(w_044_461, w_010_599, w_024_359);
  nand2 I044_465(w_044_465, w_031_175, w_012_002);
  not1 I044_473(w_044_473, w_043_009);
  or2  I044_475(w_044_475, w_008_211, w_025_100);
  not1 I044_487(w_044_487, w_004_305);
  not1 I044_496(w_044_496, w_007_362);
  nand2 I044_497(w_044_497, w_017_036, w_022_031);
  and2 I044_499(w_044_499, w_027_037, w_034_048);
  or2  I044_500(w_044_500, w_004_213, w_022_097);
  not1 I044_502(w_044_502, w_035_059);
  nand2 I044_507(w_044_507, w_039_371, w_021_085);
  nand2 I044_510(w_044_510, w_017_190, w_032_512);
  not1 I044_514(w_044_514, w_017_343);
  or2  I044_518(w_044_518, w_002_093, w_019_012);
  not1 I044_521(w_044_521, w_032_186);
  and2 I044_532(w_044_532, w_009_338, w_012_150);
  not1 I044_534(w_044_534, w_015_110);
  nand2 I044_535(w_044_535, w_026_110, w_012_061);
  not1 I044_540(w_044_540, w_007_282);
  not1 I044_544(w_044_544, w_033_512);
  and2 I044_559(w_044_559, w_007_281, w_031_422);
  or2  I044_562(w_044_562, w_026_152, w_007_449);
  nand2 I044_563(w_044_563, w_030_399, w_018_043);
  or2  I044_564(w_044_564, w_001_004, w_023_144);
  or2  I044_569(w_044_569, w_018_043, w_012_228);
  not1 I044_571(w_044_571, w_012_076);
  and2 I044_573(w_044_573, w_002_537, w_001_004);
  and2 I044_574(w_044_574, w_033_407, w_026_049);
  or2  I044_577(w_044_577, w_016_002, w_027_040);
  or2  I044_583(w_044_583, w_020_252, w_024_015);
  or2  I044_587(w_044_587, w_018_037, w_020_063);
  nand2 I044_588(w_044_588, w_021_039, w_030_219);
  not1 I044_589(w_044_589, w_006_025);
  and2 I044_598(w_044_598, w_002_596, w_037_045);
  not1 I044_599(w_044_599, w_006_241);
  and2 I044_603(w_044_603, w_039_578, w_009_315);
  or2  I044_608(w_044_608, w_034_056, w_011_378);
  or2  I044_610(w_044_610, w_023_181, w_007_265);
  and2 I044_611(w_044_611, w_001_031, w_034_050);
  and2 I044_616(w_044_616, w_040_070, w_030_152);
  or2  I044_628(w_044_628, w_001_036, w_015_653);
  or2  I044_632(w_044_632, w_023_042, w_017_370);
  nand2 I044_643(w_044_643, w_040_294, w_003_048);
  and2 I044_646(w_044_646, w_007_040, w_008_726);
  not1 I044_650(w_044_650, w_031_154);
  nand2 I044_652(w_044_652, w_037_154, w_032_163);
  not1 I044_653(w_044_653, w_040_691);
  or2  I044_657(w_044_657, w_022_041, w_037_338);
  not1 I044_658(w_044_658, w_003_001);
  not1 I044_662(w_044_662, w_015_093);
  and2 I044_663(w_044_663, w_034_000, w_036_091);
  or2  I044_666(w_044_666, w_021_202, w_008_692);
  or2  I044_670(w_044_670, w_036_012, w_032_568);
  and2 I044_673(w_044_673, w_017_211, w_041_334);
  not1 I044_675(w_044_675, w_037_008);
  and2 I044_681(w_044_681, w_007_258, w_018_025);
  not1 I044_684(w_044_684, w_031_520);
  or2  I044_686(w_044_686, w_018_015, w_021_236);
  nand2 I044_687(w_044_687, w_020_175, w_001_002);
  and2 I044_689(w_044_689, w_000_174, w_038_012);
  or2  I044_690(w_044_690, w_011_011, w_010_697);
  and2 I044_691(w_044_691, w_017_099, w_038_234);
  nand2 I044_694(w_044_694, w_043_045, w_007_104);
  and2 I044_705(w_044_705, w_010_178, w_032_219);
  not1 I044_710(w_044_710, w_039_258);
  nand2 I044_712(w_044_712, w_023_196, w_040_542);
  not1 I044_713(w_044_713, w_005_131);
  nand2 I044_719(w_044_719, w_009_523, w_022_349);
  or2  I044_721(w_044_721, w_012_211, w_007_029);
  or2  I044_722(w_044_722, w_039_003, w_004_158);
  and2 I044_723(w_044_723, w_016_007, w_020_171);
  or2  I044_740(w_044_740, w_029_026, w_016_007);
  not1 I044_743(w_044_743, w_043_003);
  not1 I044_746(w_044_746, w_042_139);
  or2  I045_000(w_045_000, w_025_234, w_041_185);
  nand2 I045_001(w_045_001, w_000_366, w_037_064);
  not1 I045_002(w_045_002, w_013_578);
  or2  I045_003(w_045_003, w_010_209, w_031_116);
  nand2 I045_005(w_045_005, w_021_231, w_021_230);
  not1 I045_006(w_045_006, w_020_255);
  nand2 I045_007(w_045_007, w_007_041, w_010_004);
  or2  I045_009(w_045_009, w_029_061, w_025_166);
  or2  I045_012(w_045_012, w_027_169, w_041_528);
  and2 I045_013(w_045_013, w_010_775, w_018_027);
  and2 I045_014(w_045_014, w_035_001, w_024_191);
  not1 I045_016(w_045_016, w_000_516);
  nand2 I045_017(w_045_017, w_019_017, w_028_503);
  or2  I045_020(w_045_020, w_033_493, w_014_043);
  and2 I045_023(w_045_023, w_001_012, w_042_197);
  nand2 I045_024(w_045_024, w_025_083, w_035_036);
  and2 I045_026(w_045_026, w_016_000, w_001_025);
  and2 I045_029(w_045_029, w_027_058, w_038_077);
  nand2 I045_034(w_045_034, w_017_028, w_009_539);
  not1 I045_038(w_045_038, w_041_086);
  nand2 I045_039(w_045_039, w_036_074, w_029_114);
  or2  I045_041(w_045_041, w_015_354, w_041_231);
  and2 I045_043(w_045_043, w_040_486, w_008_125);
  not1 I045_044(w_045_044, w_030_022);
  not1 I045_047(w_045_047, w_028_070);
  nand2 I045_048(w_045_048, w_005_245, w_015_543);
  and2 I045_049(w_045_049, w_000_017, w_001_032);
  or2  I045_050(w_045_050, w_003_059, w_040_373);
  nand2 I045_052(w_045_052, w_032_092, w_018_011);
  not1 I045_055(w_045_055, w_008_650);
  and2 I045_057(w_045_057, w_039_668, w_027_008);
  not1 I045_060(w_045_060, w_040_235);
  not1 I045_063(w_045_063, w_022_125);
  not1 I045_067(w_045_067, w_013_330);
  and2 I045_068(w_045_068, w_013_090, w_030_078);
  nand2 I045_069(w_045_069, w_020_476, w_040_343);
  nand2 I045_071(w_045_071, w_041_663, w_019_014);
  and2 I045_074(w_045_074, w_009_476, w_012_221);
  nand2 I045_075(w_045_075, w_004_202, w_030_275);
  nand2 I045_083(w_045_083, w_007_094, w_039_459);
  and2 I045_084(w_045_084, w_005_043, w_001_015);
  and2 I045_088(w_045_088, w_017_187, w_007_219);
  not1 I045_091(w_045_091, w_015_591);
  and2 I045_092(w_045_092, w_030_224, w_022_030);
  nand2 I045_100(w_045_100, w_011_351, w_026_502);
  not1 I045_102(w_045_102, w_042_455);
  not1 I045_105(w_045_105, w_022_168);
  nand2 I045_106(w_045_106, w_006_166, w_028_201);
  or2  I045_108(w_045_108, w_037_088, w_014_158);
  not1 I045_109(w_045_109, w_019_019);
  or2  I045_117(w_045_117, w_043_014, w_026_012);
  or2  I045_118(w_045_118, w_028_173, w_026_007);
  nand2 I045_124(w_045_124, w_030_226, w_044_564);
  or2  I045_126(w_045_126, w_019_005, w_018_003);
  and2 I045_129(w_045_129, w_022_263, w_000_078);
  or2  I045_130(w_045_130, w_039_145, w_028_005);
  nand2 I045_131(w_045_131, w_028_569, w_025_219);
  or2  I045_138(w_045_138, w_018_043, w_041_593);
  nand2 I045_139(w_045_139, w_032_143, w_016_004);
  and2 I045_144(w_045_144, w_040_163, w_017_430);
  nand2 I045_148(w_045_148, w_026_395, w_038_185);
  not1 I045_149(w_045_149, w_002_239);
  not1 I045_151(w_045_151, w_010_722);
  not1 I045_157(w_045_157, w_002_253);
  nand2 I045_158(w_045_158, w_005_070, w_036_178);
  or2  I045_160(w_045_160, w_041_625, w_018_036);
  nand2 I045_161(w_045_161, w_029_012, w_039_161);
  nand2 I045_166(w_045_166, w_023_076, w_000_618);
  nand2 I045_167(w_045_167, w_032_209, w_015_417);
  not1 I045_168(w_045_168, w_024_182);
  and2 I045_169(w_045_169, w_030_307, w_013_046);
  or2  I045_170(w_045_170, w_042_229, w_022_297);
  not1 I045_172(w_045_172, w_004_160);
  or2  I045_174(w_045_174, w_027_199, w_020_189);
  not1 I045_176(w_045_176, w_036_459);
  not1 I045_177(w_045_177, w_000_768);
  and2 I045_180(w_045_180, w_021_023, w_038_402);
  and2 I045_181(w_045_181, w_037_312, w_010_451);
  nand2 I045_182(w_045_182, w_020_162, w_018_009);
  and2 I045_186(w_045_186, w_000_689, w_024_496);
  not1 I045_189(w_045_189, w_038_066);
  nand2 I045_191(w_045_191, w_019_016, w_009_161);
  and2 I045_196(w_045_196, w_029_110, w_036_348);
  or2  I045_197(w_045_197, w_030_047, w_013_526);
  or2  I045_198(w_045_198, w_008_011, w_004_004);
  or2  I045_199(w_045_199, w_012_125, w_044_160);
  not1 I045_204(w_045_204, w_017_132);
  nand2 I045_205(w_045_205, w_026_109, w_009_117);
  nand2 I045_206(w_045_206, w_021_149, w_037_093);
  not1 I045_210(w_045_210, w_019_000);
  nand2 I045_212(w_045_212, w_006_018, w_006_055);
  or2  I045_215(w_045_215, w_036_330, w_044_502);
  or2  I045_219(w_045_219, w_014_002, w_012_214);
  or2  I045_220(w_045_220, w_008_067, w_020_244);
  not1 I045_224(w_045_224, w_027_049);
  or2  I045_225(w_045_225, w_008_414, w_044_559);
  not1 I045_226(w_045_226, w_018_026);
  nand2 I045_227(w_045_227, w_034_062, w_024_517);
  nand2 I045_228(w_045_228, w_024_209, w_040_371);
  not1 I045_230(w_045_230, w_019_005);
  nand2 I045_231(w_045_231, w_018_041, w_030_184);
  and2 I045_235(w_045_235, w_004_133, w_020_347);
  or2  I045_239(w_045_239, w_021_026, w_024_253);
  and2 I045_242(w_045_242, w_011_443, w_039_108);
  and2 I045_245(w_045_245, w_015_051, w_030_017);
  and2 I045_255(w_045_255, w_015_421, w_006_134);
  not1 I045_258(w_045_258, w_040_080);
  not1 I045_259(w_045_259, w_032_280);
  nand2 I045_260(w_045_260, w_007_033, w_002_221);
  or2  I045_264(w_045_264, w_018_015, w_019_020);
  nand2 I045_265(w_045_265, w_014_142, w_035_020);
  or2  I045_266(w_045_266, w_015_082, w_039_185);
  nand2 I045_267(w_045_267, w_042_267, w_000_117);
  not1 I045_268(w_045_268, w_026_295);
  and2 I045_269(w_045_269, w_003_051, w_036_165);
  and2 I045_270(w_045_270, w_000_314, w_036_060);
  not1 I045_271(w_045_271, w_010_416);
  not1 I045_272(w_045_272, w_031_055);
  nand2 I045_274(w_045_274, w_021_102, w_033_256);
  and2 I045_276(w_045_276, w_041_339, w_044_562);
  not1 I045_277(w_045_277, w_028_491);
  not1 I045_280(w_045_280, w_032_039);
  and2 I045_282(w_045_282, w_000_514, w_004_218);
  not1 I045_283(w_045_283, w_018_016);
  and2 I045_284(w_045_284, w_014_201, w_000_208);
  and2 I045_286(w_045_286, w_019_008, w_002_069);
  or2  I045_287(w_045_287, w_034_034, w_026_038);
  not1 I045_289(w_045_289, w_041_194);
  and2 I045_290(w_045_290, w_015_435, w_018_034);
  or2  I045_291(w_045_291, w_025_157, w_033_718);
  not1 I045_292(w_045_292, w_025_290);
  nand2 I045_293(w_045_293, w_000_474, w_006_158);
  nand2 I045_294(w_045_294, w_002_673, w_025_012);
  or2  I045_296(w_045_296, w_022_294, w_010_059);
  nand2 I045_300(w_045_300, w_021_001, w_033_094);
  and2 I045_304(w_045_304, w_031_581, w_022_134);
  nand2 I045_305(w_045_305, w_027_047, w_042_050);
  not1 I045_307(w_045_307, w_027_007);
  nand2 I045_308(w_045_308, w_003_028, w_012_131);
  not1 I045_310(w_045_310, w_012_243);
  nand2 I045_311(w_045_311, w_033_100, w_007_306);
  not1 I045_314(w_045_314, w_027_099);
  and2 I045_315(w_045_315, w_039_302, w_015_017);
  and2 I045_317(w_045_317, w_002_368, w_033_084);
  nand2 I045_319(w_045_319, w_012_335, w_036_271);
  or2  I045_321(w_045_321, w_016_006, w_001_013);
  or2  I045_323(w_045_323, w_039_522, w_030_392);
  not1 I045_326(w_045_326, w_002_055);
  or2  I045_327(w_045_327, w_038_368, w_020_288);
  or2  I045_330(w_045_330, w_015_346, w_010_369);
  and2 I045_331(w_045_331, w_007_459, w_003_057);
  or2  I045_332(w_045_332, w_028_283, w_038_152);
  not1 I045_333(w_045_333, w_000_447);
  nand2 I045_334(w_045_334, w_028_149, w_037_210);
  nand2 I045_335(w_045_335, w_024_101, w_004_017);
  not1 I045_336(w_045_336, w_021_015);
  and2 I045_337(w_045_337, w_043_041, w_002_342);
  or2  I045_338(w_045_338, w_016_002, w_012_140);
  nand2 I045_344(w_045_344, w_009_573, w_000_474);
  nand2 I045_345(w_045_345, w_016_008, w_002_343);
  and2 I045_348(w_045_348, w_028_248, w_044_646);
  or2  I045_353(w_045_353, w_011_043, w_003_052);
  nand2 I045_358(w_045_358, w_008_170, w_044_158);
  and2 I045_359(w_045_359, w_005_077, w_015_051);
  not1 I045_361(w_045_361, w_043_040);
  and2 I045_362(w_045_362, w_041_178, w_017_073);
  not1 I045_366(w_045_366, w_026_617);
  not1 I045_367(w_045_367, w_006_107);
  and2 I045_368(w_045_368, w_035_059, w_006_007);
  and2 I045_369(w_045_369, w_009_144, w_011_007);
  not1 I045_375(w_045_375, w_039_519);
  and2 I045_378(w_045_378, w_002_170, w_031_059);
  nand2 I045_379(w_045_379, w_044_267, w_028_252);
  or2  I045_381(w_045_381, w_016_007, w_014_269);
  nand2 I045_386(w_045_386, w_029_077, w_024_188);
  and2 I045_388(w_045_388, w_012_127, w_044_268);
  and2 I045_389(w_045_389, w_014_015, w_001_032);
  and2 I045_390(w_045_390, w_029_078, w_031_520);
  or2  I045_400(w_045_400, w_012_327, w_028_270);
  not1 I045_401(w_045_401, w_034_039);
  and2 I045_405(w_045_405, w_030_268, w_007_367);
  not1 I045_407(w_045_407, w_040_713);
  nand2 I045_409(w_045_411, w_015_580, w_045_410);
  not1 I045_410(w_045_412, w_045_411);
  nand2 I045_411(w_045_413, w_045_412, w_012_084);
  and2 I045_412(w_045_414, w_045_413, w_045_429);
  nand2 I045_413(w_045_410, w_006_094, w_045_414);
  nand2 I045_414(w_045_419, w_007_332, w_045_418);
  or2  I045_415(w_045_420, w_045_419, w_025_251);
  and2 I045_416(w_045_421, w_045_420, w_040_704);
  or2  I045_417(w_045_422, w_043_009, w_045_421);
  or2  I045_418(w_045_423, w_045_422, w_037_345);
  not1 I045_419(w_045_424, w_045_423);
  and2 I045_420(w_045_425, w_009_501, w_045_424);
  or2  I045_421(w_045_426, w_045_425, w_008_344);
  and2 I045_422(w_045_427, w_027_148, w_045_426);
  not1 I045_423(w_045_418, w_045_414);
  and2 I045_424(w_045_429, w_015_259, w_045_427);
  nand2 I046_002(w_046_002, w_017_429, w_043_033);
  nand2 I046_009(w_046_009, w_016_005, w_000_610);
  and2 I046_010(w_046_010, w_041_206, w_008_548);
  nand2 I046_013(w_046_013, w_025_104, w_045_118);
  nand2 I046_015(w_046_015, w_034_020, w_000_371);
  or2  I046_023(w_046_023, w_024_010, w_000_035);
  or2  I046_024(w_046_024, w_003_017, w_037_030);
  and2 I046_025(w_046_025, w_029_103, w_026_358);
  or2  I046_028(w_046_028, w_034_015, w_010_227);
  not1 I046_029(w_046_029, w_021_232);
  nand2 I046_031(w_046_031, w_004_463, w_000_206);
  nand2 I046_033(w_046_033, w_016_002, w_009_126);
  and2 I046_037(w_046_037, w_043_001, w_043_043);
  not1 I046_039(w_046_039, w_040_698);
  nand2 I046_041(w_046_041, w_019_002, w_042_181);
  nand2 I046_042(w_046_042, w_045_100, w_034_065);
  not1 I046_047(w_046_047, w_015_020);
  or2  I046_050(w_046_050, w_020_472, w_022_298);
  or2  I046_052(w_046_052, w_021_098, w_035_110);
  and2 I046_057(w_046_057, w_029_006, w_002_214);
  or2  I046_058(w_046_058, w_002_608, w_036_265);
  and2 I046_059(w_046_059, w_019_001, w_006_206);
  or2  I046_061(w_046_061, w_042_132, w_042_195);
  nand2 I046_062(w_046_062, w_035_037, w_036_066);
  or2  I046_068(w_046_068, w_038_308, w_000_245);
  and2 I046_073(w_046_073, w_010_241, w_042_010);
  not1 I046_074(w_046_074, w_025_099);
  nand2 I046_082(w_046_082, w_036_044, w_028_475);
  nand2 I046_085(w_046_085, w_033_011, w_017_430);
  or2  I046_092(w_046_092, w_021_062, w_018_005);
  nand2 I046_096(w_046_096, w_007_121, w_018_024);
  not1 I046_097(w_046_097, w_004_444);
  and2 I046_099(w_046_099, w_022_401, w_042_320);
  not1 I046_100(w_046_100, w_029_015);
  or2  I046_101(w_046_101, w_007_016, w_041_046);
  and2 I046_104(w_046_104, w_009_094, w_039_103);
  not1 I046_106(w_046_106, w_004_058);
  not1 I046_110(w_046_110, w_011_150);
  and2 I046_118(w_046_118, w_044_373, w_018_011);
  not1 I046_120(w_046_120, w_004_115);
  or2  I046_121(w_046_121, w_030_258, w_028_368);
  not1 I046_127(w_046_127, w_009_135);
  and2 I046_129(w_046_129, w_011_486, w_016_003);
  not1 I046_132(w_046_132, w_045_068);
  and2 I046_137(w_046_137, w_011_119, w_009_025);
  and2 I046_143(w_046_143, w_014_008, w_040_096);
  and2 I046_164(w_046_164, w_044_165, w_020_096);
  and2 I046_168(w_046_168, w_026_136, w_042_178);
  nand2 I046_171(w_046_171, w_028_526, w_044_461);
  or2  I046_172(w_046_172, w_024_119, w_034_044);
  and2 I046_174(w_046_174, w_004_048, w_009_145);
  not1 I046_176(w_046_176, w_019_010);
  or2  I046_184(w_046_184, w_031_259, w_027_090);
  and2 I046_189(w_046_189, w_033_310, w_035_006);
  and2 I046_194(w_046_194, w_023_002, w_045_348);
  not1 I046_196(w_046_196, w_011_088);
  or2  I046_197(w_046_197, w_002_500, w_023_078);
  and2 I046_201(w_046_201, w_045_174, w_012_047);
  not1 I046_209(w_046_209, w_024_535);
  nand2 I046_210(w_046_210, w_038_396, w_040_166);
  or2  I046_211(w_046_211, w_036_006, w_020_166);
  not1 I046_222(w_046_222, w_005_159);
  or2  I046_229(w_046_229, w_022_036, w_035_096);
  or2  I046_230(w_046_230, w_015_476, w_015_413);
  or2  I046_232(w_046_232, w_012_037, w_002_229);
  not1 I046_234(w_046_234, w_038_597);
  not1 I046_236(w_046_236, w_037_313);
  nand2 I046_238(w_046_238, w_025_124, w_027_045);
  and2 I046_240(w_046_240, w_040_086, w_017_166);
  or2  I046_246(w_046_246, w_018_007, w_003_059);
  and2 I046_247(w_046_247, w_027_167, w_018_029);
  or2  I046_248(w_046_248, w_040_393, w_005_134);
  and2 I046_250(w_046_250, w_018_034, w_014_124);
  nand2 I046_255(w_046_255, w_001_021, w_005_091);
  and2 I046_261(w_046_261, w_017_314, w_006_109);
  and2 I046_263(w_046_263, w_018_035, w_028_550);
  and2 I046_264(w_046_264, w_036_240, w_042_346);
  nand2 I046_267(w_046_267, w_020_080, w_017_013);
  nand2 I046_270(w_046_270, w_008_475, w_001_030);
  nand2 I046_272(w_046_272, w_020_135, w_040_257);
  not1 I046_279(w_046_279, w_041_315);
  or2  I046_284(w_046_284, w_000_216, w_016_002);
  and2 I046_288(w_046_288, w_015_544, w_009_502);
  or2  I046_292(w_046_292, w_037_147, w_031_136);
  and2 I046_294(w_046_294, w_032_197, w_032_221);
  nand2 I046_297(w_046_297, w_024_057, w_024_166);
  and2 I046_298(w_046_298, w_024_482, w_015_046);
  not1 I046_299(w_046_299, w_040_221);
  and2 I046_300(w_046_300, w_007_396, w_016_008);
  not1 I046_302(w_046_302, w_015_131);
  or2  I046_303(w_046_303, w_041_354, w_035_051);
  not1 I046_304(w_046_304, w_013_400);
  nand2 I046_314(w_046_314, w_022_005, w_025_228);
  or2  I046_318(w_046_318, w_042_165, w_040_299);
  and2 I046_319(w_046_319, w_007_342, w_008_221);
  and2 I046_323(w_046_323, w_044_159, w_036_296);
  nand2 I046_330(w_046_330, w_033_207, w_002_042);
  or2  I046_334(w_046_334, w_036_251, w_029_055);
  not1 I046_336(w_046_336, w_011_302);
  not1 I046_338(w_046_338, w_030_203);
  or2  I046_339(w_046_339, w_021_165, w_021_066);
  or2  I046_341(w_046_341, w_032_052, w_021_175);
  nand2 I046_346(w_046_346, w_040_609, w_039_360);
  or2  I046_351(w_046_351, w_009_426, w_009_186);
  nand2 I046_356(w_046_356, w_034_020, w_028_152);
  or2  I046_360(w_046_360, w_018_010, w_011_090);
  nand2 I046_372(w_046_372, w_000_751, w_042_099);
  and2 I046_373(w_046_373, w_035_097, w_022_214);
  or2  I046_377(w_046_377, w_021_201, w_029_061);
  or2  I046_387(w_046_387, w_042_293, w_002_549);
  or2  I046_389(w_046_389, w_032_192, w_040_367);
  and2 I046_390(w_046_390, w_030_064, w_008_411);
  nand2 I046_394(w_046_394, w_040_316, w_020_086);
  not1 I046_397(w_046_397, w_017_517);
  and2 I046_401(w_046_401, w_040_519, w_019_019);
  not1 I046_414(w_046_414, w_008_030);
  and2 I046_422(w_046_422, w_016_006, w_035_085);
  and2 I046_425(w_046_425, w_039_604, w_044_347);
  or2  I046_427(w_046_427, w_005_021, w_036_120);
  not1 I046_429(w_046_429, w_005_052);
  nand2 I046_432(w_046_432, w_029_077, w_024_207);
  nand2 I046_435(w_046_435, w_003_074, w_023_210);
  and2 I046_436(w_046_436, w_044_093, w_016_001);
  nand2 I046_443(w_046_443, w_008_128, w_034_064);
  not1 I046_447(w_046_447, w_002_368);
  or2  I046_450(w_046_450, w_044_013, w_035_126);
  nand2 I046_452(w_046_452, w_010_459, w_017_629);
  nand2 I046_456(w_046_456, w_013_148, w_008_202);
  and2 I046_459(w_046_459, w_027_046, w_017_597);
  not1 I046_463(w_046_463, w_012_112);
  or2  I046_467(w_046_467, w_043_000, w_019_009);
  not1 I046_472(w_046_472, w_044_563);
  nand2 I046_477(w_046_477, w_018_025, w_026_551);
  and2 I046_478(w_046_478, w_042_414, w_007_033);
  not1 I046_480(w_046_480, w_019_009);
  nand2 I046_483(w_046_483, w_012_062, w_008_046);
  or2  I046_484(w_046_484, w_034_066, w_007_094);
  and2 I046_494(w_046_494, w_042_023, w_029_023);
  or2  I046_496(w_046_496, w_023_208, w_007_016);
  and2 I046_509(w_046_509, w_001_005, w_003_041);
  nand2 I046_515(w_046_515, w_015_546, w_034_069);
  not1 I046_516(w_046_516, w_035_074);
  or2  I046_517(w_046_517, w_015_633, w_025_038);
  not1 I046_525(w_046_525, w_015_521);
  nand2 I046_526(w_046_526, w_039_714, w_008_381);
  nand2 I046_532(w_046_532, w_020_181, w_030_355);
  or2  I046_545(w_046_545, w_041_628, w_014_256);
  nand2 I046_551(w_046_551, w_008_358, w_006_002);
  not1 I046_561(w_046_561, w_034_060);
  nand2 I046_562(w_046_562, w_001_017, w_022_175);
  or2  I046_564(w_046_564, w_035_104, w_005_053);
  and2 I046_571(w_046_571, w_030_179, w_007_109);
  nand2 I046_575(w_046_575, w_018_030, w_027_054);
  nand2 I046_576(w_046_576, w_012_225, w_041_336);
  not1 I046_580(w_046_580, w_030_132);
  and2 I046_583(w_046_583, w_033_363, w_043_005);
  not1 I046_593(w_046_593, w_036_035);
  and2 I046_598(w_046_598, w_018_042, w_045_071);
  not1 I046_599(w_046_599, w_008_557);
  not1 I046_604(w_046_604, w_000_606);
  and2 I046_606(w_046_606, w_023_113, w_042_018);
  not1 I046_608(w_046_608, w_028_287);
  or2  I046_609(w_046_609, w_013_436, w_040_324);
  not1 I046_611(w_046_611, w_012_125);
  nand2 I046_612(w_046_612, w_024_229, w_022_376);
  and2 I046_616(w_046_616, w_041_282, w_029_110);
  or2  I046_619(w_046_619, w_038_149, w_032_574);
  or2  I046_620(w_046_620, w_033_236, w_025_148);
  nand2 I046_625(w_046_625, w_027_178, w_043_041);
  and2 I046_627(w_046_627, w_003_079, w_015_198);
  and2 I046_630(w_046_630, w_008_524, w_044_681);
  not1 I046_631(w_046_631, w_019_003);
  not1 I046_632(w_046_632, w_000_153);
  nand2 I046_637(w_046_637, w_026_669, w_007_354);
  or2  I046_646(w_046_646, w_035_039, w_034_012);
  nand2 I046_647(w_046_647, w_023_066, w_028_013);
  and2 I046_655(w_046_655, w_039_069, w_010_009);
  not1 I046_659(w_046_659, w_042_125);
  nand2 I046_660(w_046_660, w_024_176, w_016_003);
  not1 I046_662(w_046_662, w_039_267);
  or2  I046_677(w_046_677, w_040_440, w_006_039);
  not1 I046_686(w_046_686, w_009_036);
  and2 I046_698(w_046_698, w_007_130, w_044_332);
  and2 I046_699(w_046_699, w_033_590, w_013_164);
  or2  I046_702(w_046_702, w_027_118, w_040_129);
  and2 I046_704(w_046_704, w_010_002, w_033_698);
  nand2 I046_712(w_046_712, w_013_069, w_022_006);
  nand2 I047_001(w_047_001, w_022_316, w_018_033);
  not1 I047_002(w_047_002, w_005_226);
  or2  I047_005(w_047_005, w_025_253, w_009_342);
  or2  I047_006(w_047_006, w_038_005, w_034_039);
  or2  I047_007(w_047_007, w_034_000, w_042_116);
  nand2 I047_008(w_047_008, w_043_000, w_027_194);
  and2 I047_013(w_047_013, w_024_126, w_038_456);
  nand2 I047_014(w_047_014, w_004_388, w_035_000);
  nand2 I047_018(w_047_018, w_008_268, w_046_459);
  nand2 I047_021(w_047_021, w_023_071, w_015_481);
  nand2 I047_023(w_047_023, w_020_462, w_034_058);
  and2 I047_024(w_047_024, w_011_492, w_006_020);
  or2  I047_031(w_047_031, w_027_078, w_024_275);
  nand2 I047_032(w_047_032, w_030_364, w_030_053);
  nand2 I047_033(w_047_033, w_026_570, w_027_007);
  or2  I047_038(w_047_038, w_017_659, w_006_077);
  or2  I047_040(w_047_040, w_005_312, w_008_688);
  and2 I047_042(w_047_042, w_046_050, w_026_550);
  and2 I047_045(w_047_045, w_004_098, w_013_161);
  or2  I047_047(w_047_047, w_003_060, w_026_494);
  not1 I047_049(w_047_049, w_007_254);
  nand2 I047_050(w_047_050, w_004_329, w_001_032);
  and2 I047_051(w_047_051, w_023_054, w_013_087);
  nand2 I047_054(w_047_054, w_011_626, w_045_005);
  nand2 I047_065(w_047_065, w_001_005, w_012_102);
  and2 I047_070(w_047_070, w_032_189, w_004_335);
  or2  I047_072(w_047_072, w_019_001, w_026_154);
  or2  I047_073(w_047_073, w_009_370, w_042_295);
  nand2 I047_077(w_047_077, w_042_034, w_000_682);
  and2 I047_080(w_047_080, w_029_015, w_002_503);
  not1 I047_087(w_047_087, w_019_010);
  nand2 I047_088(w_047_088, w_036_009, w_005_314);
  and2 I047_090(w_047_090, w_028_392, w_026_126);
  nand2 I047_099(w_047_099, w_044_390, w_020_391);
  not1 I047_105(w_047_105, w_045_180);
  or2  I047_106(w_047_106, w_042_123, w_013_183);
  or2  I047_107(w_047_107, w_007_444, w_001_015);
  not1 I047_113(w_047_113, w_015_168);
  nand2 I047_115(w_047_115, w_013_511, w_041_212);
  or2  I047_116(w_047_116, w_005_043, w_046_432);
  and2 I047_118(w_047_118, w_036_004, w_020_209);
  or2  I047_119(w_047_119, w_035_039, w_023_122);
  or2  I047_121(w_047_121, w_004_374, w_031_463);
  nand2 I047_124(w_047_124, w_028_006, w_028_441);
  not1 I047_125(w_047_125, w_001_021);
  nand2 I047_126(w_047_126, w_015_369, w_015_386);
  nand2 I047_129(w_047_129, w_010_692, w_038_559);
  or2  I047_132(w_047_132, w_013_102, w_045_049);
  and2 I047_134(w_047_134, w_016_000, w_011_583);
  and2 I047_136(w_047_136, w_007_020, w_026_660);
  and2 I047_137(w_047_137, w_031_256, w_009_159);
  not1 I047_139(w_047_139, w_026_178);
  not1 I047_140(w_047_140, w_038_047);
  not1 I047_141(w_047_141, w_033_065);
  and2 I047_142(w_047_142, w_016_007, w_030_235);
  and2 I047_147(w_047_147, w_016_008, w_026_660);
  or2  I047_148(w_047_148, w_042_290, w_029_103);
  and2 I047_152(w_047_152, w_043_041, w_019_010);
  nand2 I047_154(w_047_154, w_044_033, w_007_389);
  nand2 I047_155(w_047_155, w_036_163, w_027_008);
  or2  I047_158(w_047_158, w_028_433, w_025_088);
  and2 I047_174(w_047_174, w_001_021, w_040_689);
  or2  I047_177(w_047_177, w_011_222, w_035_006);
  nand2 I047_185(w_047_185, w_008_720, w_021_141);
  not1 I047_188(w_047_188, w_020_173);
  and2 I047_191(w_047_191, w_035_021, w_000_116);
  not1 I047_192(w_047_192, w_002_495);
  not1 I047_197(w_047_197, w_030_265);
  and2 I047_199(w_047_199, w_036_298, w_014_141);
  and2 I047_201(w_047_201, w_028_022, w_041_537);
  nand2 I047_205(w_047_205, w_036_146, w_005_168);
  not1 I047_206(w_047_206, w_020_012);
  and2 I047_207(w_047_207, w_007_316, w_002_511);
  not1 I047_208(w_047_208, w_043_008);
  and2 I047_209(w_047_209, w_017_102, w_005_318);
  not1 I047_210(w_047_210, w_042_401);
  and2 I047_211(w_047_211, w_046_302, w_000_061);
  and2 I047_214(w_047_214, w_028_044, w_000_391);
  nand2 I047_215(w_047_215, w_023_191, w_036_099);
  or2  I047_219(w_047_219, w_042_413, w_041_444);
  and2 I047_220(w_047_220, w_041_172, w_029_087);
  or2  I047_221(w_047_221, w_009_478, w_013_156);
  not1 I047_224(w_047_224, w_023_024);
  not1 I047_225(w_047_225, w_007_074);
  or2  I047_229(w_047_229, w_004_486, w_017_601);
  not1 I047_230(w_047_230, w_045_315);
  not1 I047_232(w_047_232, w_042_209);
  or2  I047_237(w_047_237, w_021_177, w_029_063);
  not1 I047_238(w_047_238, w_007_044);
  nand2 I047_239(w_047_239, w_029_023, w_041_181);
  nand2 I047_245(w_047_245, w_042_237, w_042_292);
  nand2 I047_246(w_047_246, w_022_309, w_025_296);
  nand2 I047_248(w_047_248, w_026_448, w_037_303);
  not1 I047_249(w_047_249, w_032_072);
  not1 I047_251(w_047_251, w_017_631);
  nand2 I047_254(w_047_254, w_040_246, w_003_029);
  and2 I047_255(w_047_255, w_032_022, w_023_081);
  not1 I047_256(w_047_256, w_020_291);
  and2 I047_263(w_047_263, w_029_114, w_042_362);
  nand2 I047_265(w_047_265, w_044_571, w_014_021);
  not1 I047_267(w_047_267, w_033_329);
  nand2 I047_268(w_047_268, w_000_197, w_026_712);
  not1 I047_270(w_047_270, w_042_304);
  and2 I047_273(w_047_273, w_035_065, w_005_138);
  not1 I047_275(w_047_275, w_036_336);
  not1 I047_276(w_047_276, w_036_313);
  and2 I047_277(w_047_277, w_033_486, w_045_068);
  not1 I047_279(w_047_279, w_037_010);
  or2  I047_280(w_047_280, w_021_142, w_020_494);
  nand2 I047_283(w_047_283, w_010_739, w_011_151);
  and2 I047_287(w_047_287, w_001_015, w_031_390);
  not1 I047_288(w_047_288, w_021_106);
  or2  I047_290(w_047_290, w_005_210, w_038_385);
  nand2 I047_291(w_047_291, w_027_156, w_016_001);
  not1 I047_294(w_047_294, w_017_023);
  and2 I047_295(w_047_295, w_015_040, w_045_231);
  nand2 I047_298(w_047_298, w_006_030, w_014_026);
  or2  I047_299(w_047_299, w_022_367, w_015_269);
  or2  I047_305(w_047_305, w_008_710, w_009_011);
  nand2 I047_306(w_047_306, w_046_304, w_034_003);
  nand2 I047_307(w_047_307, w_025_127, w_046_284);
  or2  I047_309(w_047_309, w_035_022, w_023_189);
  or2  I047_311(w_047_311, w_041_685, w_018_016);
  and2 I047_317(w_047_317, w_043_010, w_039_055);
  nand2 I047_318(w_047_318, w_033_740, w_034_030);
  nand2 I047_320(w_047_320, w_008_024, w_026_431);
  nand2 I047_323(w_047_323, w_004_380, w_013_209);
  or2  I047_325(w_047_325, w_017_108, w_042_456);
  and2 I047_327(w_047_327, w_029_099, w_044_746);
  or2  I047_329(w_047_329, w_009_070, w_037_122);
  or2  I047_330(w_047_330, w_020_050, w_034_037);
  and2 I047_340(w_047_340, w_038_508, w_017_186);
  nand2 I047_341(w_047_341, w_042_428, w_020_090);
  and2 I047_342(w_047_342, w_007_196, w_044_514);
  not1 I047_350(w_047_350, w_005_162);
  not1 I047_359(w_047_359, w_003_008);
  not1 I047_360(w_047_360, w_010_109);
  and2 I047_362(w_047_362, w_036_256, w_018_022);
  nand2 I047_367(w_047_367, w_015_087, w_015_319);
  and2 I047_370(w_047_370, w_007_241, w_044_414);
  or2  I047_379(w_047_379, w_035_069, w_016_008);
  not1 I047_383(w_047_383, w_018_005);
  nand2 I047_390(w_047_390, w_029_010, w_019_004);
  and2 I047_394(w_047_394, w_023_065, w_044_616);
  or2  I047_396(w_047_396, w_020_203, w_042_072);
  and2 I047_399(w_047_399, w_041_661, w_018_009);
  not1 I047_404(w_047_404, w_010_581);
  not1 I047_407(w_047_407, w_014_187);
  nand2 I047_413(w_047_413, w_009_374, w_020_404);
  nand2 I047_419(w_047_419, w_015_127, w_032_092);
  not1 I047_420(w_047_420, w_017_017);
  nand2 I047_422(w_047_422, w_028_186, w_026_238);
  or2  I047_428(w_047_428, w_017_460, w_026_424);
  not1 I047_436(w_047_436, w_005_001);
  or2  I047_443(w_047_443, w_046_330, w_023_139);
  not1 I047_454(w_047_454, w_029_042);
  or2  I047_458(w_047_458, w_042_288, w_018_034);
  and2 I047_465(w_047_465, w_035_074, w_004_130);
  or2  I047_469(w_047_469, w_021_124, w_004_310);
  nand2 I048_000(w_048_000, w_023_102, w_004_135);
  not1 I048_001(w_048_001, w_010_566);
  not1 I048_002(w_048_002, w_039_061);
  and2 I048_003(w_048_003, w_039_267, w_025_096);
  not1 I048_004(w_048_004, w_043_039);
  or2  I048_005(w_048_005, w_044_673, w_015_120);
  nand2 I048_006(w_048_006, w_042_182, w_022_195);
  or2  I048_007(w_048_007, w_022_164, w_044_273);
  and2 I048_008(w_048_008, w_035_031, w_019_004);
  or2  I048_009(w_048_009, w_010_359, w_017_274);
  nand2 I048_010(w_048_010, w_042_265, w_029_066);
  or2  I048_011(w_048_011, w_027_088, w_010_746);
  not1 I048_012(w_048_012, w_017_086);
  not1 I048_013(w_048_013, w_008_562);
  nand2 I048_014(w_048_014, w_030_278, w_028_196);
  not1 I048_015(w_048_015, w_015_335);
  or2  I048_016(w_048_016, w_009_016, w_028_021);
  not1 I048_017(w_048_017, w_046_435);
  and2 I048_018(w_048_018, w_032_449, w_002_297);
  and2 I048_019(w_048_019, w_005_019, w_022_117);
  and2 I049_002(w_049_002, w_001_029, w_010_458);
  nand2 I049_003(w_049_003, w_012_300, w_046_609);
  and2 I049_004(w_049_004, w_038_610, w_028_374);
  not1 I049_005(w_049_005, w_013_161);
  or2  I049_006(w_049_006, w_031_574, w_010_121);
  nand2 I049_009(w_049_009, w_008_583, w_032_105);
  and2 I049_011(w_049_011, w_002_032, w_030_240);
  nand2 I049_012(w_049_012, w_042_297, w_035_097);
  and2 I049_016(w_049_016, w_012_313, w_039_588);
  nand2 I049_017(w_049_017, w_039_348, w_009_328);
  and2 I049_018(w_049_018, w_045_138, w_024_365);
  or2  I049_019(w_049_019, w_015_526, w_021_188);
  not1 I049_020(w_049_020, w_024_280);
  and2 I049_021(w_049_021, w_046_058, w_031_470);
  not1 I049_022(w_049_022, w_030_200);
  not1 I049_023(w_049_023, w_047_042);
  nand2 I049_024(w_049_024, w_018_025, w_036_298);
  and2 I049_025(w_049_025, w_038_604, w_026_383);
  nand2 I049_026(w_049_026, w_015_102, w_038_516);
  not1 I049_029(w_049_029, w_041_513);
  not1 I049_033(w_049_033, w_018_032);
  or2  I049_035(w_049_035, w_021_171, w_035_013);
  nand2 I049_036(w_049_036, w_023_043, w_005_144);
  not1 I049_041(w_049_041, w_034_017);
  or2  I049_045(w_049_045, w_005_015, w_007_058);
  or2  I049_047(w_049_047, w_039_586, w_001_028);
  or2  I049_049(w_049_049, w_040_045, w_016_001);
  not1 I049_060(w_049_060, w_001_011);
  or2  I049_065(w_049_065, w_001_004, w_032_533);
  not1 I049_066(w_049_066, w_032_134);
  or2  I049_070(w_049_070, w_016_000, w_008_702);
  nand2 I049_074(w_049_074, w_028_011, w_043_024);
  or2  I049_076(w_049_076, w_004_062, w_008_668);
  not1 I049_079(w_049_079, w_002_443);
  or2  I049_081(w_049_081, w_029_005, w_006_077);
  not1 I049_083(w_049_083, w_032_191);
  or2  I049_093(w_049_093, w_012_143, w_021_225);
  not1 I049_095(w_049_095, w_038_059);
  and2 I049_101(w_049_101, w_022_370, w_026_225);
  nand2 I049_104(w_049_104, w_031_083, w_037_242);
  not1 I049_107(w_049_107, w_007_204);
  not1 I049_110(w_049_110, w_009_247);
  or2  I049_111(w_049_111, w_024_180, w_047_239);
  not1 I049_112(w_049_112, w_020_246);
  nand2 I049_116(w_049_116, w_039_634, w_010_674);
  nand2 I049_119(w_049_119, w_004_225, w_020_230);
  or2  I049_120(w_049_120, w_034_011, w_044_292);
  and2 I049_121(w_049_121, w_012_031, w_021_169);
  nand2 I049_124(w_049_124, w_022_268, w_031_033);
  and2 I049_130(w_049_130, w_013_478, w_021_045);
  nand2 I049_131(w_049_131, w_003_011, w_013_197);
  or2  I049_134(w_049_134, w_022_211, w_016_005);
  and2 I049_135(w_049_135, w_018_016, w_044_670);
  not1 I049_140(w_049_140, w_027_180);
  or2  I049_144(w_049_144, w_027_170, w_015_192);
  not1 I049_153(w_049_153, w_010_314);
  nand2 I049_154(w_049_154, w_030_070, w_018_035);
  and2 I049_161(w_049_161, w_015_664, w_047_224);
  nand2 I049_162(w_049_162, w_019_009, w_012_024);
  or2  I049_164(w_049_164, w_038_418, w_033_492);
  nand2 I049_165(w_049_165, w_008_121, w_007_294);
  and2 I049_166(w_049_166, w_031_095, w_042_201);
  nand2 I049_168(w_049_168, w_026_471, w_038_163);
  not1 I049_171(w_049_171, w_011_546);
  or2  I049_172(w_049_172, w_019_016, w_043_008);
  nand2 I049_174(w_049_174, w_032_559, w_005_130);
  nand2 I049_175(w_049_175, w_048_003, w_038_457);
  not1 I049_177(w_049_177, w_000_559);
  or2  I049_178(w_049_178, w_011_014, w_047_070);
  or2  I049_179(w_049_179, w_047_469, w_025_126);
  nand2 I049_182(w_049_182, w_032_013, w_006_059);
  or2  I049_184(w_049_184, w_027_049, w_039_300);
  nand2 I049_187(w_049_187, w_030_241, w_033_085);
  and2 I049_189(w_049_189, w_000_067, w_023_003);
  or2  I049_190(w_049_190, w_003_053, w_033_143);
  nand2 I049_192(w_049_192, w_025_002, w_003_044);
  nand2 I049_200(w_049_200, w_009_359, w_018_005);
  not1 I049_202(w_049_202, w_038_550);
  nand2 I049_204(w_049_204, w_000_443, w_024_518);
  or2  I049_207(w_049_207, w_044_687, w_000_582);
  and2 I049_209(w_049_209, w_009_086, w_035_069);
  and2 I049_210(w_049_210, w_001_005, w_048_016);
  and2 I049_217(w_049_217, w_030_215, w_028_070);
  not1 I049_220(w_049_220, w_043_009);
  not1 I049_222(w_049_222, w_044_507);
  not1 I049_223(w_049_223, w_029_059);
  or2  I049_231(w_049_231, w_033_537, w_000_702);
  or2  I049_232(w_049_232, w_035_067, w_047_107);
  and2 I049_233(w_049_233, w_038_465, w_024_121);
  and2 I049_236(w_049_236, w_008_409, w_043_007);
  not1 I049_237(w_049_237, w_019_013);
  and2 I049_238(w_049_238, w_020_561, w_033_442);
  and2 I049_239(w_049_239, w_036_101, w_011_162);
  not1 I049_240(w_049_240, w_040_283);
  not1 I049_246(w_049_246, w_037_117);
  nand2 I049_249(w_049_249, w_033_328, w_036_046);
  nand2 I049_252(w_049_252, w_015_499, w_031_066);
  and2 I049_253(w_049_253, w_031_218, w_003_000);
  and2 I049_254(w_049_254, w_037_062, w_046_515);
  not1 I049_256(w_049_256, w_039_471);
  and2 I049_259(w_049_259, w_038_458, w_020_042);
  and2 I049_260(w_049_260, w_013_556, w_031_410);
  and2 I049_263(w_049_263, w_016_004, w_040_139);
  or2  I049_267(w_049_267, w_000_012, w_029_091);
  not1 I049_268(w_049_268, w_037_123);
  and2 I049_269(w_049_269, w_007_262, w_008_722);
  or2  I049_271(w_049_271, w_019_011, w_010_586);
  nand2 I049_272(w_049_272, w_042_220, w_025_228);
  or2  I049_277(w_049_277, w_013_217, w_036_114);
  nand2 I049_278(w_049_278, w_047_298, w_004_129);
  not1 I049_279(w_049_279, w_031_147);
  not1 I049_280(w_049_280, w_002_672);
  not1 I049_281(w_049_281, w_007_316);
  and2 I049_282(w_049_282, w_006_147, w_008_285);
  nand2 I049_285(w_049_285, w_044_652, w_021_234);
  or2  I049_288(w_049_288, w_029_092, w_038_508);
  or2  I049_290(w_049_290, w_011_052, w_009_027);
  or2  I049_292(w_049_292, w_015_139, w_002_213);
  not1 I049_294(w_049_294, w_023_093);
  and2 I049_299(w_049_299, w_013_134, w_032_281);
  nand2 I049_303(w_049_303, w_030_214, w_039_429);
  nand2 I049_304(w_049_304, w_009_442, w_010_398);
  and2 I049_305(w_049_305, w_021_263, w_013_043);
  not1 I049_309(w_049_309, w_001_032);
  not1 I049_312(w_049_312, w_033_321);
  or2  I049_313(w_049_313, w_029_001, w_033_756);
  nand2 I049_320(w_049_320, w_024_183, w_035_029);
  nand2 I049_322(w_049_322, w_006_083, w_006_124);
  or2  I049_324(w_049_324, w_019_010, w_003_029);
  or2  I049_334(w_049_334, w_036_050, w_025_133);
  and2 I049_335(w_049_335, w_018_026, w_035_025);
  not1 I049_337(w_049_337, w_012_330);
  nand2 I049_338(w_049_338, w_048_003, w_010_370);
  or2  I049_341(w_049_341, w_033_539, w_023_166);
  or2  I049_342(w_049_342, w_015_339, w_020_602);
  not1 I049_347(w_049_347, w_041_587);
  and2 I049_348(w_049_348, w_026_326, w_002_417);
  or2  I049_358(w_049_358, w_030_318, w_043_040);
  nand2 I049_362(w_049_362, w_029_078, w_020_331);
  or2  I049_363(w_049_363, w_021_022, w_000_520);
  nand2 I049_372(w_049_372, w_039_213, w_028_465);
  and2 I049_373(w_049_373, w_010_412, w_004_126);
  not1 I049_386(w_049_386, w_003_020);
  nand2 I049_389(w_049_389, w_011_080, w_038_188);
  nand2 I049_397(w_049_397, w_033_340, w_040_663);
  and2 I049_411(w_049_411, w_005_084, w_021_193);
  not1 I050_004(w_050_004, w_046_025);
  not1 I050_007(w_050_007, w_034_034);
  and2 I050_008(w_050_008, w_000_451, w_025_006);
  nand2 I050_009(w_050_009, w_036_112, w_031_604);
  or2  I050_010(w_050_010, w_043_003, w_004_043);
  or2  I050_011(w_050_011, w_002_045, w_029_108);
  not1 I050_012(w_050_012, w_039_559);
  and2 I050_016(w_050_016, w_018_039, w_013_463);
  not1 I050_017(w_050_017, w_019_001);
  and2 I050_021(w_050_021, w_000_459, w_008_521);
  and2 I050_024(w_050_024, w_021_023, w_003_034);
  or2  I050_027(w_050_027, w_005_029, w_047_106);
  or2  I050_030(w_050_030, w_040_049, w_035_122);
  and2 I050_031(w_050_031, w_039_506, w_014_043);
  and2 I050_032(w_050_032, w_045_016, w_003_053);
  or2  I050_034(w_050_034, w_002_313, w_024_029);
  and2 I050_035(w_050_035, w_027_062, w_048_017);
  or2  I050_036(w_050_036, w_041_659, w_033_329);
  or2  I050_037(w_050_037, w_033_318, w_030_172);
  or2  I050_041(w_050_041, w_035_084, w_043_040);
  or2  I050_042(w_050_042, w_026_427, w_000_059);
  nand2 I050_045(w_050_045, w_009_042, w_026_718);
  and2 I050_046(w_050_046, w_013_001, w_040_015);
  or2  I050_047(w_050_047, w_034_020, w_034_039);
  and2 I050_048(w_050_048, w_029_047, w_047_005);
  nand2 I050_050(w_050_050, w_020_530, w_007_273);
  or2  I050_054(w_050_054, w_011_109, w_012_289);
  not1 I050_056(w_050_056, w_045_124);
  nand2 I050_058(w_050_058, w_022_320, w_036_075);
  and2 I050_062(w_050_062, w_006_068, w_000_715);
  and2 I050_064(w_050_064, w_003_084, w_036_289);
  not1 I050_069(w_050_069, w_019_007);
  or2  I050_071(w_050_071, w_038_115, w_023_154);
  nand2 I050_072(w_050_072, w_010_291, w_032_183);
  not1 I050_079(w_050_079, w_024_183);
  or2  I050_080(w_050_080, w_017_325, w_042_044);
  or2  I050_082(w_050_082, w_006_217, w_047_132);
  and2 I050_085(w_050_085, w_045_311, w_018_004);
  or2  I050_091(w_050_091, w_046_435, w_044_301);
  nand2 I050_093(w_050_093, w_031_118, w_024_542);
  or2  I050_099(w_050_099, w_045_108, w_043_001);
  and2 I050_101(w_050_101, w_008_457, w_017_184);
  nand2 I050_103(w_050_103, w_010_532, w_011_177);
  and2 I050_105(w_050_105, w_000_292, w_035_055);
  and2 I050_106(w_050_106, w_028_216, w_003_057);
  or2  I050_110(w_050_110, w_023_160, w_022_098);
  not1 I050_112(w_050_112, w_033_762);
  not1 I050_117(w_050_117, w_047_290);
  not1 I050_119(w_050_119, w_004_415);
  and2 I050_120(w_050_120, w_037_185, w_025_104);
  nand2 I050_121(w_050_121, w_021_154, w_014_000);
  and2 I050_123(w_050_123, w_015_019, w_031_214);
  and2 I050_127(w_050_127, w_011_233, w_044_684);
  and2 I050_130(w_050_130, w_017_070, w_047_458);
  and2 I050_131(w_050_131, w_018_012, w_041_035);
  not1 I050_133(w_050_133, w_047_360);
  or2  I050_135(w_050_135, w_033_149, w_010_039);
  not1 I050_136(w_050_136, w_014_179);
  and2 I050_138(w_050_138, w_044_497, w_008_136);
  nand2 I050_141(w_050_141, w_011_219, w_020_457);
  nand2 I050_148(w_050_148, w_020_002, w_029_109);
  and2 I050_149(w_050_149, w_004_213, w_024_202);
  or2  I050_152(w_050_152, w_038_575, w_018_015);
  or2  I050_161(w_050_161, w_022_124, w_008_223);
  and2 I050_164(w_050_164, w_036_328, w_009_397);
  or2  I050_175(w_050_175, w_014_167, w_006_021);
  and2 I050_177(w_050_177, w_007_210, w_039_317);
  nand2 I050_186(w_050_186, w_011_263, w_040_312);
  and2 I050_199(w_050_199, w_013_270, w_032_279);
  nand2 I050_205(w_050_205, w_005_019, w_011_137);
  not1 I050_207(w_050_207, w_010_230);
  and2 I050_211(w_050_211, w_014_264, w_046_564);
  and2 I050_222(w_050_222, w_030_240, w_017_102);
  or2  I050_226(w_050_226, w_039_422, w_042_072);
  and2 I050_234(w_050_234, w_023_006, w_045_235);
  and2 I050_236(w_050_236, w_008_572, w_040_295);
  nand2 I050_237(w_050_237, w_014_248, w_013_235);
  or2  I050_238(w_050_238, w_013_168, w_019_008);
  not1 I050_242(w_050_242, w_027_109);
  not1 I050_247(w_050_247, w_013_091);
  not1 I050_257(w_050_257, w_041_670);
  nand2 I050_259(w_050_259, w_016_005, w_016_007);
  not1 I050_263(w_050_263, w_032_425);
  and2 I050_264(w_050_264, w_023_077, w_014_053);
  not1 I050_266(w_050_266, w_024_007);
  or2  I050_267(w_050_267, w_039_428, w_025_008);
  nand2 I050_271(w_050_271, w_032_185, w_033_587);
  or2  I050_274(w_050_274, w_018_002, w_006_027);
  and2 I050_280(w_050_280, w_044_137, w_034_017);
  nand2 I050_292(w_050_292, w_011_398, w_009_463);
  or2  I050_295(w_050_295, w_029_020, w_020_013);
  nand2 I050_305(w_050_305, w_017_453, w_022_052);
  or2  I050_306(w_050_306, w_017_365, w_011_344);
  nand2 I050_309(w_050_309, w_011_462, w_035_015);
  and2 I050_312(w_050_312, w_042_101, w_023_012);
  not1 I050_317(w_050_317, w_011_094);
  and2 I050_322(w_050_322, w_003_077, w_000_065);
  not1 I050_323(w_050_323, w_046_010);
  and2 I050_333(w_050_333, w_016_000, w_025_126);
  or2  I050_334(w_050_334, w_030_049, w_019_013);
  or2  I050_344(w_050_344, w_034_026, w_026_657);
  not1 I050_348(w_050_348, w_011_206);
  or2  I050_359(w_050_359, w_015_126, w_032_195);
  nand2 I050_363(w_050_363, w_016_007, w_039_175);
  and2 I050_365(w_050_365, w_004_378, w_014_089);
  or2  I050_367(w_050_367, w_006_021, w_034_004);
  nand2 I050_373(w_050_373, w_007_455, w_049_269);
  nand2 I050_376(w_050_376, w_007_001, w_007_324);
  or2  I050_377(w_050_377, w_044_276, w_012_308);
  and2 I050_384(w_050_384, w_011_265, w_044_719);
  or2  I050_385(w_050_385, w_005_010, w_020_038);
  and2 I050_386(w_050_386, w_030_097, w_019_010);
  and2 I050_388(w_050_388, w_006_056, w_000_345);
  and2 I050_392(w_050_392, w_011_026, w_024_301);
  and2 I050_398(w_050_398, w_014_190, w_041_589);
  nand2 I050_399(w_050_399, w_048_006, w_020_429);
  nand2 I050_401(w_050_401, w_024_276, w_046_346);
  or2  I050_404(w_050_404, w_027_098, w_025_094);
  not1 I050_405(w_050_405, w_019_011);
  or2  I050_406(w_050_406, w_017_429, w_012_198);
  not1 I050_407(w_050_407, w_046_580);
  or2  I050_408(w_050_408, w_026_720, w_044_002);
  not1 I050_412(w_050_412, w_047_137);
  and2 I050_415(w_050_415, w_036_082, w_005_255);
  not1 I050_416(w_050_416, w_027_189);
  and2 I050_417(w_050_417, w_045_041, w_005_239);
  not1 I050_427(w_050_427, w_007_367);
  or2  I050_435(w_050_435, w_027_120, w_040_670);
  nand2 I050_437(w_050_437, w_020_087, w_001_011);
  nand2 I050_440(w_050_440, w_049_004, w_049_076);
  not1 I050_446(w_050_446, w_048_017);
  or2  I050_454(w_050_454, w_019_020, w_028_104);
  nand2 I050_460(w_050_460, w_015_082, w_038_385);
  or2  I050_461(w_050_461, w_018_006, w_033_121);
  and2 I050_470(w_050_470, w_029_046, w_037_146);
  or2  I050_475(w_050_475, w_011_288, w_037_011);
  nand2 I050_479(w_050_479, w_025_117, w_012_210);
  or2  I050_480(w_050_480, w_020_588, w_043_034);
  not1 I050_488(w_050_488, w_034_016);
  not1 I050_493(w_050_493, w_011_260);
  nand2 I050_500(w_050_500, w_043_006, w_030_106);
  and2 I050_510(w_050_510, w_001_031, w_018_029);
  or2  I050_514(w_050_514, w_022_117, w_032_173);
  not1 I050_520(w_050_520, w_004_478);
  or2  I050_526(w_050_526, w_007_025, w_024_193);
  and2 I050_532(w_050_532, w_044_030, w_033_253);
  and2 I050_533(w_050_533, w_009_169, w_001_034);
  not1 I050_534(w_050_534, w_023_178);
  and2 I050_537(w_050_537, w_041_673, w_027_037);
  not1 I050_543(w_050_543, w_003_074);
  nand2 I050_546(w_050_546, w_034_056, w_018_036);
  not1 I050_570(w_050_570, w_021_172);
  or2  I050_571(w_050_571, w_042_261, w_013_316);
  nand2 I050_573(w_050_573, w_024_092, w_004_453);
  or2  I050_578(w_050_578, w_004_008, w_008_409);
  and2 I050_584(w_050_584, w_048_019, w_043_018);
  nand2 I050_589(w_050_589, w_025_060, w_032_234);
  and2 I050_593(w_050_593, w_010_753, w_024_083);
  and2 I050_597(w_050_597, w_047_155, w_040_405);
  and2 I050_602(w_050_602, w_045_300, w_039_559);
  and2 I050_610(w_050_610, w_033_545, w_027_164);
  and2 I050_611(w_050_611, w_017_623, w_011_013);
  nand2 I050_612(w_050_612, w_035_120, w_001_008);
  or2  I050_621(w_050_621, w_042_317, w_026_071);
  and2 I050_626(w_050_626, w_022_388, w_035_091);
  not1 I050_627(w_050_627, w_020_517);
  nand2 I050_630(w_050_630, w_042_195, w_037_316);
  not1 I050_646(w_050_646, w_013_311);
  nand2 I051_003(w_051_003, w_033_545, w_041_433);
  nand2 I051_005(w_051_005, w_029_067, w_046_655);
  not1 I051_006(w_051_006, w_024_513);
  and2 I051_008(w_051_008, w_046_625, w_010_139);
  and2 I051_009(w_051_009, w_020_151, w_045_105);
  nand2 I051_011(w_051_011, w_050_510, w_020_003);
  and2 I051_013(w_051_013, w_030_134, w_045_108);
  nand2 I051_014(w_051_014, w_025_247, w_050_589);
  not1 I051_017(w_051_017, w_032_443);
  or2  I051_019(w_051_019, w_049_025, w_032_464);
  or2  I051_021(w_051_021, w_026_289, w_036_029);
  nand2 I051_023(w_051_023, w_032_109, w_020_098);
  or2  I051_024(w_051_024, w_026_357, w_011_104);
  nand2 I051_025(w_051_025, w_011_411, w_001_011);
  or2  I051_027(w_051_027, w_011_120, w_012_068);
  or2  I051_028(w_051_028, w_016_008, w_033_516);
  or2  I051_031(w_051_031, w_025_142, w_045_049);
  not1 I051_033(w_051_033, w_019_003);
  or2  I051_036(w_051_036, w_004_048, w_039_598);
  not1 I051_037(w_051_037, w_047_320);
  or2  I051_041(w_051_041, w_011_043, w_002_170);
  or2  I051_044(w_051_044, w_033_171, w_001_027);
  and2 I051_045(w_051_045, w_001_036, w_020_361);
  and2 I051_051(w_051_051, w_021_089, w_012_111);
  not1 I051_052(w_051_052, w_004_168);
  and2 I051_053(w_051_053, w_022_236, w_023_176);
  or2  I051_055(w_051_055, w_013_453, w_033_574);
  not1 I051_061(w_051_061, w_022_062);
  not1 I051_062(w_051_062, w_035_042);
  and2 I051_063(w_051_063, w_008_490, w_006_005);
  or2  I051_067(w_051_067, w_044_295, w_013_311);
  and2 I051_069(w_051_069, w_019_003, w_000_400);
  or2  I051_073(w_051_073, w_017_036, w_015_200);
  and2 I051_074(w_051_074, w_008_048, w_034_023);
  not1 I051_075(w_051_075, w_044_662);
  nand2 I051_078(w_051_078, w_021_262, w_017_434);
  and2 I051_080(w_051_080, w_012_089, w_001_028);
  or2  I051_081(w_051_081, w_010_298, w_034_035);
  nand2 I051_084(w_051_084, w_039_057, w_003_024);
  and2 I051_090(w_051_090, w_027_187, w_008_226);
  or2  I051_092(w_051_092, w_031_423, w_042_082);
  not1 I051_094(w_051_094, w_007_340);
  or2  I051_095(w_051_095, w_023_026, w_013_178);
  not1 I051_096(w_051_096, w_048_007);
  not1 I051_098(w_051_098, w_036_144);
  or2  I051_103(w_051_103, w_025_101, w_038_064);
  nand2 I051_105(w_051_105, w_012_233, w_042_039);
  not1 I051_106(w_051_106, w_020_322);
  nand2 I051_107(w_051_107, w_035_052, w_039_092);
  or2  I051_113(w_051_113, w_016_003, w_030_353);
  nand2 I051_115(w_051_115, w_032_129, w_033_251);
  not1 I051_117(w_051_117, w_018_002);
  and2 I051_120(w_051_120, w_044_569, w_013_274);
  nand2 I051_121(w_051_121, w_043_020, w_038_123);
  and2 I051_126(w_051_126, w_023_016, w_016_005);
  not1 I051_136(w_051_136, w_046_210);
  or2  I051_137(w_051_137, w_003_077, w_022_240);
  nand2 I051_138(w_051_138, w_022_288, w_044_632);
  not1 I051_140(w_051_140, w_021_215);
  or2  I051_141(w_051_141, w_031_150, w_011_583);
  not1 I051_147(w_051_147, w_040_238);
  nand2 I051_148(w_051_148, w_020_549, w_047_224);
  nand2 I051_150(w_051_150, w_028_374, w_013_163);
  or2  I051_157(w_051_157, w_019_002, w_008_062);
  or2  I051_159(w_051_159, w_041_349, w_007_386);
  or2  I051_162(w_051_162, w_013_323, w_043_005);
  and2 I051_165(w_051_165, w_035_105, w_004_360);
  nand2 I051_166(w_051_166, w_046_261, w_044_367);
  not1 I051_167(w_051_167, w_023_215);
  and2 I051_170(w_051_170, w_043_022, w_002_027);
  or2  I051_171(w_051_171, w_017_004, w_040_318);
  and2 I051_172(w_051_172, w_025_263, w_004_118);
  not1 I051_173(w_051_173, w_024_441);
  and2 I051_181(w_051_181, w_002_098, w_016_008);
  nand2 I051_183(w_051_183, w_018_035, w_016_002);
  not1 I051_185(w_051_185, w_034_004);
  not1 I051_186(w_051_186, w_049_282);
  or2  I051_188(w_051_188, w_036_103, w_017_229);
  not1 I051_189(w_051_189, w_001_000);
  or2  I051_195(w_051_195, w_026_056, w_050_611);
  not1 I051_196(w_051_196, w_033_012);
  nand2 I051_199(w_051_199, w_011_631, w_032_116);
  not1 I051_200(w_051_200, w_019_010);
  or2  I051_203(w_051_203, w_040_014, w_004_268);
  and2 I051_204(w_051_204, w_029_064, w_004_456);
  not1 I051_206(w_051_206, w_022_397);
  not1 I051_208(w_051_208, w_044_062);
  or2  I051_210(w_051_210, w_028_128, w_012_035);
  and2 I051_215(w_051_215, w_048_004, w_046_346);
  not1 I051_218(w_051_218, w_034_012);
  not1 I051_222(w_051_222, w_037_273);
  nand2 I051_225(w_051_225, w_004_012, w_047_002);
  nand2 I051_226(w_051_226, w_043_032, w_007_219);
  not1 I051_230(w_051_230, w_033_354);
  nand2 I051_231(w_051_231, w_003_045, w_047_309);
  or2  I051_232(w_051_232, w_017_663, w_043_006);
  and2 I051_233(w_051_233, w_024_243, w_044_610);
  or2  I051_235(w_051_235, w_050_042, w_043_002);
  or2  I051_237(w_051_237, w_004_391, w_050_292);
  not1 I051_242(w_051_242, w_009_568);
  or2  I051_243(w_051_243, w_007_124, w_033_059);
  or2  I051_244(w_051_244, w_006_198, w_007_216);
  nand2 I051_246(w_051_246, w_030_196, w_003_031);
  or2  I051_248(w_051_248, w_041_054, w_042_282);
  not1 I051_249(w_051_249, w_000_050);
  nand2 I051_250(w_051_250, w_032_208, w_003_051);
  not1 I051_256(w_051_256, w_028_483);
  and2 I051_260(w_051_260, w_045_007, w_025_009);
  not1 I051_262(w_051_262, w_008_693);
  not1 I051_263(w_051_263, w_045_083);
  and2 I051_265(w_051_265, w_024_029, w_027_040);
  not1 I051_268(w_051_268, w_031_239);
  or2  I051_275(w_051_275, w_013_185, w_012_252);
  or2  I051_279(w_051_279, w_046_031, w_001_003);
  nand2 I051_282(w_051_282, w_013_072, w_016_005);
  not1 I051_286(w_051_286, w_014_130);
  or2  I051_291(w_051_291, w_036_132, w_042_422);
  and2 I051_298(w_051_298, w_010_733, w_031_086);
  and2 I051_301(w_051_301, w_005_054, w_027_082);
  nand2 I051_303(w_051_303, w_029_101, w_034_043);
  or2  I051_307(w_051_307, w_002_302, w_022_220);
  not1 I051_308(w_051_308, w_045_002);
  and2 I051_309(w_051_309, w_014_136, w_041_342);
  not1 I051_312(w_051_312, w_047_359);
  or2  I051_313(w_051_313, w_006_029, w_016_002);
  not1 I051_317(w_051_317, w_020_183);
  nand2 I051_318(w_051_318, w_022_395, w_031_281);
  or2  I051_319(w_051_319, w_049_011, w_022_258);
  or2  I051_320(w_051_320, w_028_053, w_018_007);
  not1 I051_322(w_051_322, w_032_184);
  not1 I051_323(w_051_323, w_040_439);
  and2 I051_326(w_051_326, w_030_312, w_010_684);
  or2  I051_330(w_051_330, w_028_252, w_042_126);
  not1 I051_333(w_051_333, w_043_019);
  not1 I051_337(w_051_337, w_048_004);
  and2 I051_340(w_051_340, w_000_430, w_017_078);
  and2 I051_342(w_051_342, w_008_012, w_006_234);
  and2 I051_343(w_051_343, w_005_141, w_000_776);
  and2 I051_346(w_051_346, w_037_026, w_018_003);
  nand2 I051_348(w_051_348, w_030_316, w_046_387);
  not1 I051_349(w_051_349, w_026_621);
  and2 I051_351(w_051_351, w_005_092, w_013_301);
  and2 I051_353(w_051_353, w_042_099, w_000_777);
  or2  I051_354(w_051_354, w_035_101, w_034_012);
  not1 I051_358(w_051_358, w_050_010);
  or2  I051_366(w_051_366, w_009_088, w_003_010);
  nand2 I051_367(w_051_367, w_020_009, w_041_263);
  nand2 I051_369(w_051_369, w_004_066, w_032_011);
  nand2 I051_370(w_051_370, w_008_193, w_039_073);
  nand2 I051_372(w_051_372, w_013_545, w_016_000);
  not1 I051_378(w_051_378, w_009_239);
  not1 I051_380(w_051_380, w_013_215);
  not1 I051_381(w_051_381, w_048_016);
  not1 I051_395(w_051_395, w_037_028);
  or2  I051_398(w_051_398, w_041_326, w_014_096);
  not1 I051_406(w_051_406, w_024_056);
  and2 I052_000(w_052_000, w_011_551, w_006_242);
  not1 I052_001(w_052_001, w_028_163);
  not1 I052_002(w_052_002, w_024_103);
  not1 I052_003(w_052_003, w_046_074);
  and2 I052_004(w_052_004, w_040_386, w_029_068);
  not1 I052_005(w_052_005, w_017_127);
  nand2 I052_006(w_052_006, w_022_034, w_015_389);
  or2  I052_007(w_052_007, w_048_016, w_013_220);
  nand2 I052_008(w_052_008, w_044_418, w_008_555);
  nand2 I052_009(w_052_009, w_006_181, w_019_008);
  not1 I052_011(w_052_011, w_049_024);
  and2 I052_012(w_052_012, w_014_077, w_003_073);
  or2  I052_013(w_052_013, w_019_006, w_002_303);
  not1 I052_014(w_052_014, w_043_027);
  not1 I052_015(w_052_015, w_036_032);
  and2 I052_017(w_052_017, w_036_090, w_018_034);
  not1 I052_018(w_052_018, w_010_419);
  and2 I052_019(w_052_019, w_016_006, w_021_213);
  nand2 I052_020(w_052_020, w_011_148, w_008_244);
  nand2 I052_021(w_052_021, w_043_026, w_026_605);
  not1 I052_022(w_052_022, w_002_579);
  not1 I052_023(w_052_023, w_048_017);
  or2  I052_024(w_052_024, w_041_138, w_017_038);
  and2 I052_025(w_052_025, w_032_404, w_003_026);
  and2 I052_026(w_052_026, w_047_265, w_013_000);
  and2 I052_027(w_052_027, w_001_030, w_005_277);
  and2 I052_028(w_052_028, w_024_192, w_011_533);
  not1 I052_029(w_052_029, w_041_665);
  and2 I052_030(w_052_030, w_037_074, w_029_088);
  and2 I052_031(w_052_031, w_022_351, w_029_048);
  nand2 I052_032(w_052_032, w_008_490, w_028_527);
  nand2 I052_033(w_052_033, w_041_664, w_016_006);
  or2  I052_034(w_052_034, w_021_029, w_025_272);
  and2 I052_035(w_052_035, w_012_315, w_050_377);
  nand2 I052_036(w_052_036, w_046_662, w_006_058);
  and2 I052_037(w_052_037, w_018_014, w_020_383);
  nand2 I052_038(w_052_038, w_031_539, w_026_033);
  nand2 I052_039(w_052_039, w_021_126, w_023_143);
  nand2 I052_040(w_052_040, w_012_214, w_003_019);
  nand2 I052_041(w_052_041, w_027_015, w_022_229);
  nand2 I052_042(w_052_042, w_017_291, w_042_451);
  not1 I052_043(w_052_043, w_034_034);
  nand2 I052_044(w_052_044, w_030_226, w_051_298);
  or2  I052_045(w_052_045, w_025_257, w_004_302);
  not1 I052_046(w_052_046, w_003_046);
  nand2 I053_000(w_053_000, w_007_473, w_028_191);
  or2  I053_001(w_053_001, w_018_004, w_007_080);
  or2  I053_004(w_053_004, w_040_047, w_030_134);
  and2 I053_005(w_053_005, w_038_054, w_017_115);
  and2 I053_006(w_053_006, w_050_305, w_003_046);
  not1 I053_007(w_053_007, w_011_631);
  and2 I053_009(w_053_009, w_041_036, w_024_108);
  nand2 I053_010(w_053_010, w_011_133, w_024_013);
  nand2 I053_013(w_053_013, w_015_001, w_029_004);
  and2 I053_014(w_053_014, w_006_002, w_000_415);
  nand2 I053_015(w_053_015, w_052_024, w_024_541);
  nand2 I053_017(w_053_017, w_044_181, w_016_003);
  or2  I053_018(w_053_018, w_045_317, w_006_166);
  nand2 I053_020(w_053_020, w_010_606, w_045_158);
  and2 I053_021(w_053_021, w_045_126, w_037_051);
  nand2 I053_023(w_053_023, w_024_212, w_000_214);
  or2  I053_024(w_053_024, w_048_005, w_021_091);
  nand2 I053_025(w_053_025, w_007_359, w_013_517);
  or2  I053_026(w_053_026, w_036_272, w_046_620);
  nand2 I053_028(w_053_028, w_023_058, w_017_381);
  nand2 I053_029(w_053_029, w_004_221, w_051_113);
  not1 I053_031(w_053_031, w_051_073);
  and2 I053_033(w_053_033, w_017_260, w_051_173);
  and2 I053_034(w_053_034, w_032_471, w_004_163);
  or2  I053_035(w_053_035, w_001_023, w_013_263);
  not1 I053_037(w_053_037, w_027_183);
  and2 I053_038(w_053_038, w_025_048, w_022_382);
  or2  I053_040(w_053_040, w_036_186, w_046_002);
  and2 I053_041(w_053_041, w_030_090, w_016_008);
  not1 I053_042(w_053_042, w_029_004);
  nand2 I053_044(w_053_044, w_029_071, w_024_565);
  and2 I053_046(w_053_046, w_005_068, w_028_449);
  and2 I053_047(w_053_047, w_021_176, w_047_245);
  and2 I053_048(w_053_048, w_010_717, w_046_660);
  not1 I053_049(w_053_049, w_033_771);
  nand2 I053_050(w_053_050, w_035_027, w_033_209);
  or2  I053_051(w_053_051, w_036_312, w_014_286);
  not1 I053_053(w_053_053, w_051_121);
  not1 I053_054(w_053_054, w_052_030);
  not1 I053_055(w_053_055, w_029_055);
  nand2 I053_056(w_053_056, w_017_532, w_038_140);
  or2  I053_058(w_053_058, w_032_437, w_003_009);
  not1 I053_060(w_053_060, w_006_125);
  not1 I053_061(w_053_061, w_009_382);
  and2 I053_062(w_053_062, w_045_368, w_041_623);
  or2  I053_065(w_053_065, w_011_424, w_000_360);
  not1 I053_066(w_053_066, w_039_648);
  not1 I053_067(w_053_067, w_050_271);
  and2 I053_069(w_053_069, w_021_266, w_019_012);
  nand2 I053_070(w_053_070, w_020_125, w_031_107);
  nand2 I053_071(w_053_071, w_002_167, w_002_681);
  and2 I053_072(w_053_072, w_013_074, w_037_319);
  and2 I053_073(w_053_073, w_002_519, w_048_007);
  nand2 I053_074(w_053_074, w_051_067, w_016_003);
  or2  I053_075(w_053_075, w_010_412, w_048_014);
  or2  I053_076(w_053_076, w_012_029, w_010_431);
  and2 I053_077(w_053_077, w_018_012, w_033_509);
  nand2 I053_078(w_053_078, w_017_468, w_004_116);
  nand2 I053_079(w_053_079, w_029_023, w_013_544);
  not1 I053_080(w_053_080, w_044_371);
  or2  I053_081(w_053_081, w_007_475, w_032_028);
  and2 I053_082(w_053_082, w_006_176, w_043_038);
  and2 I053_083(w_053_083, w_032_357, w_052_031);
  and2 I053_085(w_053_085, w_034_018, w_003_077);
  not1 I053_086(w_053_086, w_048_009);
  and2 I053_087(w_053_087, w_040_692, w_029_062);
  nand2 I053_088(w_053_088, w_008_598, w_038_020);
  nand2 I053_089(w_053_089, w_008_746, w_000_513);
  nand2 I053_090(w_053_090, w_031_356, w_032_109);
  and2 I053_091(w_053_091, w_009_127, w_046_039);
  nand2 I053_092(w_053_092, w_028_264, w_000_160);
  or2  I053_093(w_053_093, w_049_179, w_042_404);
  and2 I053_094(w_053_094, w_034_041, w_050_404);
  or2  I053_095(w_053_095, w_037_301, w_048_017);
  not1 I053_096(w_053_096, w_004_045);
  not1 I053_097(w_053_097, w_016_001);
  not1 I053_098(w_053_098, w_004_111);
  not1 I053_099(w_053_099, w_006_194);
  not1 I053_101(w_053_101, w_028_008);
  not1 I053_102(w_053_102, w_044_191);
  nand2 I053_103(w_053_103, w_042_138, w_052_040);
  and2 I053_105(w_053_105, w_027_176, w_025_120);
  and2 I053_106(w_053_106, w_031_134, w_015_589);
  and2 I053_108(w_053_108, w_007_143, w_051_186);
  nand2 I053_109(w_053_109, w_025_079, w_044_338);
  not1 I053_110(w_053_110, w_023_158);
  or2  I053_111(w_053_111, w_007_070, w_035_019);
  nand2 I053_112(w_053_112, w_039_203, w_043_001);
  not1 I053_113(w_053_113, w_006_129);
  not1 I053_114(w_053_114, w_018_001);
  and2 I053_115(w_053_115, w_022_348, w_003_031);
  not1 I053_116(w_053_116, w_034_034);
  not1 I053_119(w_053_119, w_050_488);
  or2  I053_120(w_053_120, w_001_007, w_020_055);
  or2  I053_126(w_053_126, w_030_312, w_011_102);
  not1 I053_129(w_053_129, w_003_005);
  nand2 I053_131(w_053_131, w_028_094, w_021_271);
  or2  I053_132(w_053_132, w_023_146, w_049_144);
  nand2 I053_134(w_053_134, w_041_606, w_033_692);
  not1 I053_135(w_053_135, w_011_481);
  not1 I053_136(w_053_136, w_050_048);
  nand2 I053_137(w_053_137, w_041_698, w_042_271);
  not1 I053_139(w_053_139, w_006_151);
  and2 I053_140(w_053_140, w_042_146, w_001_016);
  nand2 I053_143(w_053_143, w_040_120, w_022_149);
  nand2 I053_144(w_053_144, w_043_016, w_018_024);
  nand2 I053_149(w_053_149, w_024_146, w_024_418);
  or2  I053_151(w_053_151, w_036_058, w_051_078);
  or2  I053_152(w_053_152, w_013_118, w_036_335);
  and2 I053_153(w_053_153, w_040_521, w_001_014);
  and2 I053_154(w_053_154, w_040_063, w_020_008);
  nand2 I053_155(w_053_155, w_037_257, w_035_047);
  nand2 I053_156(w_053_156, w_006_149, w_000_696);
  not1 I053_158(w_053_158, w_043_042);
  or2  I053_161(w_053_161, w_003_021, w_005_292);
  nand2 I054_001(w_054_001, w_034_009, w_002_044);
  not1 I054_003(w_054_003, w_043_006);
  and2 I054_004(w_054_004, w_035_094, w_028_056);
  nand2 I054_009(w_054_009, w_016_000, w_046_627);
  not1 I054_013(w_054_013, w_024_118);
  not1 I054_020(w_054_020, w_022_348);
  or2  I054_021(w_054_021, w_049_272, w_049_231);
  and2 I054_024(w_054_024, w_028_177, w_040_180);
  and2 I054_026(w_054_026, w_043_007, w_012_036);
  or2  I054_029(w_054_029, w_043_019, w_032_033);
  nand2 I054_033(w_054_033, w_046_598, w_027_039);
  or2  I054_035(w_054_035, w_026_136, w_048_019);
  or2  I054_041(w_054_041, w_015_565, w_028_299);
  and2 I054_043(w_054_043, w_027_060, w_036_194);
  nand2 I054_049(w_054_049, w_030_174, w_019_006);
  not1 I054_051(w_054_051, w_007_454);
  nand2 I054_055(w_054_055, w_029_067, w_014_102);
  and2 I054_058(w_054_058, w_003_059, w_005_124);
  or2  I054_061(w_054_061, w_001_020, w_041_026);
  and2 I054_066(w_054_066, w_036_079, w_044_663);
  or2  I054_068(w_054_068, w_050_017, w_012_198);
  and2 I054_071(w_054_071, w_006_157, w_012_083);
  and2 I054_073(w_054_073, w_008_426, w_022_251);
  or2  I054_074(w_054_074, w_022_261, w_045_310);
  nand2 I054_077(w_054_077, w_035_031, w_020_199);
  not1 I054_078(w_054_078, w_048_010);
  not1 I054_081(w_054_081, w_024_141);
  nand2 I054_082(w_054_082, w_043_029, w_041_628);
  nand2 I054_084(w_054_084, w_011_308, w_004_428);
  and2 I054_085(w_054_085, w_029_115, w_050_526);
  and2 I054_088(w_054_088, w_031_446, w_016_004);
  nand2 I054_089(w_054_089, w_003_058, w_005_039);
  and2 I054_095(w_054_095, w_053_074, w_018_011);
  and2 I054_096(w_054_096, w_023_064, w_028_150);
  not1 I054_098(w_054_098, w_022_234);
  and2 I054_102(w_054_102, w_009_552, w_049_009);
  or2  I054_104(w_054_104, w_016_002, w_034_008);
  nand2 I054_106(w_054_106, w_051_346, w_012_247);
  nand2 I054_109(w_054_109, w_014_234, w_013_235);
  or2  I054_114(w_054_114, w_048_007, w_032_411);
  or2  I054_116(w_054_116, w_044_475, w_012_009);
  not1 I054_122(w_054_122, w_015_220);
  or2  I054_126(w_054_126, w_022_020, w_007_374);
  or2  I054_131(w_054_131, w_011_351, w_034_066);
  nand2 I054_133(w_054_133, w_014_219, w_028_097);
  and2 I054_137(w_054_137, w_006_225, w_031_112);
  or2  I054_138(w_054_138, w_003_050, w_016_006);
  or2  I054_141(w_054_141, w_040_433, w_036_314);
  not1 I054_144(w_054_144, w_039_043);
  and2 I054_145(w_054_145, w_017_267, w_014_094);
  or2  I054_146(w_054_146, w_021_023, w_024_064);
  nand2 I054_148(w_054_148, w_019_002, w_003_037);
  nand2 I054_149(w_054_149, w_040_288, w_030_298);
  nand2 I054_150(w_054_150, w_050_627, w_019_003);
  not1 I054_151(w_054_151, w_020_065);
  not1 I054_155(w_054_155, w_025_296);
  and2 I054_157(w_054_157, w_021_195, w_006_204);
  and2 I054_161(w_054_161, w_037_246, w_003_003);
  nand2 I054_162(w_054_162, w_044_100, w_031_302);
  or2  I054_164(w_054_164, w_015_026, w_005_220);
  or2  I054_166(w_054_166, w_014_103, w_019_000);
  not1 I054_167(w_054_167, w_027_102);
  and2 I054_169(w_054_169, w_017_056, w_046_197);
  and2 I054_170(w_054_170, w_017_436, w_009_435);
  nand2 I054_173(w_054_173, w_023_162, w_032_540);
  and2 I054_176(w_054_176, w_036_295, w_048_013);
  or2  I054_178(w_054_178, w_035_006, w_016_000);
  nand2 I054_184(w_054_184, w_024_175, w_002_606);
  not1 I054_186(w_054_186, w_051_092);
  nand2 I054_190(w_054_190, w_029_063, w_022_382);
  not1 I054_194(w_054_194, w_031_472);
  not1 I054_199(w_054_199, w_043_022);
  and2 I054_203(w_054_203, w_043_030, w_017_415);
  and2 I054_214(w_054_214, w_031_153, w_013_463);
  or2  I054_228(w_054_228, w_005_244, w_040_119);
  nand2 I054_230(w_054_230, w_018_015, w_020_474);
  and2 I054_231(w_054_231, w_053_060, w_018_009);
  not1 I054_234(w_054_234, w_042_453);
  and2 I054_239(w_054_239, w_001_028, w_039_706);
  nand2 I054_240(w_054_240, w_004_468, w_007_008);
  or2  I054_252(w_054_252, w_013_521, w_035_012);
  and2 I054_256(w_054_256, w_051_055, w_027_030);
  nand2 I054_258(w_054_258, w_050_323, w_003_052);
  and2 I054_262(w_054_262, w_051_081, w_040_004);
  and2 I054_274(w_054_274, w_045_130, w_027_034);
  not1 I054_276(w_054_276, w_024_231);
  nand2 I054_279(w_054_279, w_041_441, w_045_407);
  nand2 I054_283(w_054_283, w_047_422, w_045_034);
  or2  I054_284(w_054_284, w_024_263, w_015_019);
  and2 I054_305(w_054_305, w_029_046, w_021_274);
  or2  I054_310(w_054_310, w_002_642, w_023_184);
  nand2 I054_314(w_054_314, w_041_226, w_021_100);
  and2 I054_319(w_054_319, w_010_127, w_027_189);
  nand2 I054_323(w_054_323, w_014_272, w_035_024);
  not1 I054_332(w_054_332, w_041_593);
  and2 I054_344(w_054_344, w_029_024, w_029_002);
  nand2 I054_346(w_054_346, w_048_004, w_028_022);
  nand2 I054_347(w_054_347, w_030_262, w_026_613);
  nand2 I054_365(w_054_365, w_042_025, w_010_086);
  or2  I054_394(w_054_394, w_033_002, w_036_156);
  and2 I054_410(w_054_410, w_039_099, w_047_428);
  or2  I054_412(w_054_412, w_036_304, w_048_018);
  or2  I054_415(w_054_415, w_013_414, w_017_485);
  nand2 I054_417(w_054_417, w_007_240, w_035_117);
  and2 I054_425(w_054_425, w_022_077, w_028_041);
  and2 I054_431(w_054_431, w_048_012, w_026_698);
  or2  I054_439(w_054_439, w_029_048, w_040_032);
  not1 I054_440(w_054_440, w_002_043);
  nand2 I054_456(w_054_456, w_048_003, w_033_068);
  and2 I054_463(w_054_463, w_036_336, w_039_534);
  nand2 I054_466(w_054_466, w_006_002, w_034_055);
  and2 I054_467(w_054_467, w_020_154, w_035_122);
  nand2 I054_472(w_054_472, w_005_282, w_019_017);
  nand2 I054_486(w_054_486, w_000_653, w_033_715);
  or2  I054_490(w_054_490, w_018_013, w_005_134);
  nand2 I054_494(w_054_494, w_033_703, w_020_361);
  or2  I054_502(w_054_502, w_020_260, w_033_427);
  nand2 I054_508(w_054_508, w_020_301, w_015_191);
  nand2 I054_510(w_054_510, w_047_306, w_022_389);
  nand2 I054_515(w_054_515, w_048_018, w_004_102);
  and2 I054_521(w_054_521, w_017_589, w_039_309);
  not1 I054_533(w_054_533, w_024_205);
  nand2 I054_534(w_054_534, w_044_070, w_015_144);
  nand2 I054_542(w_054_542, w_004_160, w_020_077);
  not1 I054_545(w_054_545, w_018_018);
  or2  I054_549(w_054_549, w_048_015, w_018_024);
  not1 I054_557(w_054_557, w_041_032);
  not1 I054_569(w_054_569, w_008_016);
  or2  I054_581(w_054_581, w_030_345, w_038_435);
  not1 I054_588(w_054_588, w_038_082);
  or2  I054_590(w_054_590, w_051_115, w_050_571);
  and2 I055_000(w_055_000, w_006_011, w_046_612);
  not1 I055_006(w_055_006, w_024_008);
  not1 I055_007(w_055_007, w_017_599);
  and2 I055_014(w_055_014, w_015_120, w_001_012);
  or2  I055_015(w_055_015, w_052_024, w_044_583);
  nand2 I055_018(w_055_018, w_023_009, w_047_295);
  not1 I055_022(w_055_022, w_022_084);
  not1 I055_023(w_055_023, w_052_024);
  or2  I055_027(w_055_027, w_003_034, w_004_031);
  nand2 I055_029(w_055_029, w_009_065, w_002_574);
  and2 I055_030(w_055_030, w_048_009, w_001_034);
  and2 I055_033(w_055_033, w_004_214, w_023_215);
  and2 I055_034(w_055_034, w_014_011, w_010_387);
  not1 I055_035(w_055_035, w_007_106);
  or2  I055_036(w_055_036, w_017_523, w_048_013);
  or2  I055_038(w_055_038, w_010_277, w_023_107);
  nand2 I055_039(w_055_039, w_000_465, w_013_447);
  nand2 I055_040(w_055_040, w_023_214, w_052_028);
  not1 I055_041(w_055_041, w_049_320);
  and2 I055_042(w_055_042, w_002_067, w_022_386);
  not1 I055_043(w_055_043, w_015_281);
  nand2 I055_045(w_055_045, w_004_337, w_008_676);
  and2 I055_046(w_055_046, w_045_260, w_033_207);
  and2 I055_047(w_055_047, w_012_088, w_033_001);
  or2  I055_049(w_055_049, w_047_001, w_008_658);
  or2  I055_051(w_055_051, w_007_260, w_049_223);
  not1 I055_052(w_055_052, w_053_113);
  or2  I055_053(w_055_053, w_047_329, w_026_234);
  and2 I055_057(w_055_057, w_023_003, w_029_035);
  not1 I055_058(w_055_058, w_023_158);
  and2 I055_059(w_055_059, w_022_079, w_017_419);
  and2 I055_061(w_055_061, w_026_127, w_002_701);
  nand2 I055_064(w_055_064, w_013_179, w_037_164);
  not1 I055_066(w_055_066, w_045_314);
  not1 I055_068(w_055_068, w_012_077);
  nand2 I055_072(w_055_072, w_040_091, w_031_309);
  not1 I055_074(w_055_074, w_003_048);
  and2 I055_076(w_055_076, w_028_313, w_017_178);
  nand2 I055_077(w_055_077, w_028_173, w_040_428);
  and2 I055_078(w_055_078, w_012_058, w_000_757);
  not1 I055_080(w_055_080, w_039_652);
  nand2 I055_082(w_055_082, w_045_013, w_019_019);
  not1 I055_084(w_055_084, w_009_070);
  nand2 I055_085(w_055_085, w_021_205, w_030_308);
  or2  I055_088(w_055_088, w_020_080, w_005_107);
  not1 I055_089(w_055_089, w_025_082);
  not1 I055_090(w_055_090, w_048_019);
  not1 I055_091(w_055_091, w_045_369);
  not1 I055_094(w_055_094, w_048_001);
  and2 I055_095(w_055_095, w_021_029, w_013_272);
  or2  I055_096(w_055_096, w_009_042, w_053_161);
  or2  I055_097(w_055_097, w_028_050, w_033_278);
  or2  I055_103(w_055_103, w_035_009, w_039_007);
  nand2 I055_104(w_055_104, w_041_060, w_022_280);
  nand2 I055_106(w_055_106, w_035_072, w_005_121);
  or2  I055_108(w_055_108, w_015_469, w_000_131);
  nand2 I055_110(w_055_110, w_022_152, w_007_084);
  and2 I055_114(w_055_114, w_021_168, w_039_538);
  or2  I055_116(w_055_116, w_016_000, w_011_021);
  and2 I055_122(w_055_122, w_030_050, w_001_019);
  not1 I055_123(w_055_123, w_017_525);
  not1 I055_124(w_055_124, w_043_012);
  nand2 I055_127(w_055_127, w_030_157, w_036_201);
  not1 I055_129(w_055_129, w_002_438);
  and2 I055_131(w_055_131, w_014_111, w_039_361);
  and2 I055_132(w_055_132, w_043_030, w_007_283);
  or2  I055_133(w_055_133, w_034_051, w_025_002);
  or2  I055_137(w_055_137, w_011_167, w_012_297);
  not1 I055_138(w_055_138, w_051_243);
  not1 I055_139(w_055_139, w_039_016);
  or2  I055_140(w_055_140, w_032_191, w_029_012);
  and2 I055_142(w_055_142, w_000_636, w_031_453);
  and2 I055_145(w_055_145, w_046_632, w_035_020);
  or2  I055_154(w_055_154, w_010_265, w_017_089);
  or2  I055_155(w_055_155, w_043_009, w_046_704);
  nand2 I055_156(w_055_156, w_051_024, w_043_016);
  or2  I055_161(w_055_161, w_035_010, w_028_109);
  or2  I055_164(w_055_164, w_021_072, w_005_095);
  and2 I055_165(w_055_165, w_043_021, w_050_079);
  or2  I055_168(w_055_168, w_049_202, w_031_287);
  or2  I055_174(w_055_174, w_027_024, w_033_016);
  and2 I055_180(w_055_180, w_041_007, w_012_219);
  or2  I055_181(w_055_181, w_014_043, w_043_033);
  and2 I055_183(w_055_183, w_023_108, w_020_278);
  or2  I055_185(w_055_185, w_024_377, w_053_140);
  nand2 I055_187(w_055_187, w_053_066, w_015_091);
  or2  I055_191(w_055_191, w_000_295, w_010_335);
  or2  I055_192(w_055_192, w_045_131, w_041_512);
  or2  I055_197(w_055_197, w_021_158, w_025_169);
  nand2 I055_200(w_055_200, w_005_014, w_019_000);
  or2  I055_202(w_055_202, w_023_104, w_018_024);
  nand2 I055_204(w_055_204, w_015_276, w_040_346);
  nand2 I055_207(w_055_207, w_054_151, w_007_437);
  not1 I055_213(w_055_213, w_048_002);
  or2  I055_215(w_055_215, w_019_004, w_036_165);
  not1 I055_219(w_055_219, w_023_007);
  nand2 I055_220(w_055_220, w_037_033, w_010_164);
  and2 I055_225(w_055_225, w_012_003, w_047_132);
  or2  I055_226(w_055_226, w_003_037, w_028_160);
  or2  I055_227(w_055_227, w_052_003, w_035_030);
  not1 I055_234(w_055_234, w_027_182);
  not1 I055_236(w_055_236, w_029_086);
  not1 I055_239(w_055_239, w_022_381);
  not1 I055_240(w_055_240, w_035_060);
  or2  I055_241(w_055_241, w_052_006, w_049_140);
  not1 I055_242(w_055_242, w_041_026);
  or2  I055_243(w_055_243, w_000_130, w_054_314);
  or2  I055_254(w_055_254, w_004_019, w_051_320);
  not1 I055_255(w_055_255, w_026_396);
  not1 I055_257(w_055_257, w_029_026);
  or2  I055_258(w_055_258, w_029_081, w_020_007);
  not1 I055_259(w_055_259, w_016_007);
  nand2 I055_262(w_055_262, w_000_143, w_016_002);
  nand2 I055_265(w_055_265, w_047_211, w_003_060);
  nand2 I055_266(w_055_266, w_018_027, w_012_016);
  nand2 I055_267(w_055_267, w_025_307, w_042_077);
  or2  I055_276(w_055_276, w_031_136, w_035_050);
  or2  I055_279(w_055_279, w_030_375, w_001_025);
  nand2 I055_282(w_055_282, w_017_314, w_043_027);
  and2 I055_285(w_055_285, w_043_009, w_014_042);
  or2  I055_286(w_055_286, w_021_225, w_012_006);
  not1 I055_287(w_055_287, w_047_065);
  not1 I055_290(w_055_290, w_036_190);
  or2  I055_294(w_055_294, w_007_198, w_052_017);
  or2  I055_297(w_055_297, w_002_012, w_047_125);
  or2  I055_298(w_055_298, w_024_275, w_038_135);
  nand2 I055_302(w_055_302, w_026_267, w_028_091);
  not1 I055_307(w_055_307, w_013_293);
  and2 I055_309(w_055_309, w_046_303, w_037_044);
  and2 I055_312(w_055_312, w_028_277, w_014_168);
  nand2 I055_313(w_055_313, w_042_135, w_050_398);
  not1 I055_316(w_055_316, w_033_076);
  or2  I055_324(w_055_324, w_043_035, w_025_124);
  not1 I055_330(w_055_330, w_053_077);
  or2  I055_337(w_055_337, w_046_015, w_021_170);
  not1 I055_339(w_055_339, w_016_000);
  not1 I055_344(w_055_344, w_039_415);
  or2  I055_345(w_055_345, w_010_042, w_054_515);
  and2 I056_007(w_056_007, w_023_016, w_012_002);
  nand2 I056_008(w_056_008, w_035_081, w_011_112);
  nand2 I056_009(w_056_009, w_008_172, w_032_124);
  nand2 I056_012(w_056_012, w_033_323, w_025_012);
  nand2 I056_016(w_056_016, w_044_284, w_039_143);
  and2 I056_017(w_056_017, w_040_014, w_030_350);
  nand2 I056_020(w_056_020, w_025_209, w_023_200);
  not1 I056_022(w_056_022, w_016_006);
  or2  I056_030(w_056_030, w_028_115, w_040_484);
  or2  I056_033(w_056_033, w_012_258, w_009_625);
  nand2 I056_035(w_056_035, w_027_090, w_038_043);
  and2 I056_037(w_056_037, w_042_150, w_017_001);
  or2  I056_038(w_056_038, w_012_127, w_027_032);
  nand2 I056_039(w_056_039, w_044_033, w_002_445);
  and2 I056_044(w_056_044, w_032_240, w_026_015);
  and2 I056_046(w_056_046, w_049_334, w_006_005);
  and2 I056_048(w_056_048, w_036_146, w_020_463);
  and2 I056_049(w_056_049, w_031_204, w_010_559);
  and2 I056_051(w_056_051, w_036_033, w_001_013);
  or2  I056_057(w_056_057, w_009_190, w_040_565);
  and2 I056_058(w_056_058, w_032_449, w_045_020);
  or2  I056_069(w_056_069, w_042_275, w_010_228);
  not1 I056_070(w_056_070, w_017_052);
  or2  I056_071(w_056_071, w_034_068, w_000_220);
  or2  I056_081(w_056_081, w_049_154, w_048_018);
  not1 I056_082(w_056_082, w_027_159);
  nand2 I056_084(w_056_084, w_020_177, w_034_071);
  not1 I056_088(w_056_088, w_000_066);
  nand2 I056_089(w_056_089, w_014_288, w_050_399);
  and2 I056_090(w_056_090, w_051_044, w_053_031);
  and2 I056_094(w_056_094, w_033_263, w_007_224);
  not1 I056_106(w_056_106, w_006_077);
  nand2 I056_108(w_056_108, w_052_004, w_034_075);
  and2 I056_119(w_056_119, w_041_529, w_026_114);
  and2 I056_120(w_056_120, w_030_089, w_029_116);
  not1 I056_123(w_056_123, w_055_312);
  or2  I056_129(w_056_129, w_023_013, w_029_097);
  nand2 I056_141(w_056_141, w_015_370, w_022_333);
  not1 I056_145(w_056_145, w_023_031);
  or2  I056_154(w_056_154, w_051_204, w_002_488);
  nand2 I056_172(w_056_172, w_012_118, w_029_051);
  not1 I056_176(w_056_176, w_043_028);
  nand2 I056_184(w_056_184, w_017_655, w_038_495);
  not1 I056_200(w_056_200, w_018_028);
  nand2 I056_214(w_056_214, w_029_020, w_055_265);
  and2 I056_224(w_056_224, w_014_088, w_049_285);
  or2  I056_229(w_056_229, w_038_601, w_033_184);
  nand2 I056_231(w_056_231, w_032_078, w_017_064);
  not1 I056_232(w_056_232, w_002_486);
  or2  I056_235(w_056_235, w_026_413, w_018_002);
  or2  I056_238(w_056_238, w_006_002, w_035_022);
  and2 I056_241(w_056_241, w_020_075, w_029_096);
  and2 I056_242(w_056_242, w_055_053, w_046_247);
  not1 I056_244(w_056_244, w_032_493);
  or2  I056_249(w_056_249, w_007_315, w_009_226);
  nand2 I056_250(w_056_250, w_010_542, w_042_201);
  or2  I056_252(w_056_252, w_048_013, w_014_140);
  nand2 I056_254(w_056_254, w_032_515, w_030_105);
  nand2 I056_255(w_056_255, w_039_553, w_050_312);
  and2 I056_267(w_056_267, w_053_074, w_009_151);
  or2  I056_280(w_056_280, w_019_004, w_043_016);
  nand2 I056_289(w_056_289, w_005_239, w_019_001);
  nand2 I056_303(w_056_303, w_052_039, w_048_010);
  and2 I056_314(w_056_314, w_053_075, w_005_040);
  not1 I056_317(w_056_317, w_031_072);
  or2  I056_323(w_056_323, w_030_053, w_055_077);
  or2  I056_332(w_056_332, w_013_322, w_012_246);
  and2 I056_348(w_056_348, w_031_160, w_049_168);
  and2 I056_357(w_056_357, w_026_027, w_053_081);
  or2  I056_365(w_056_365, w_012_069, w_028_102);
  nand2 I056_369(w_056_369, w_005_083, w_031_129);
  or2  I056_371(w_056_371, w_004_315, w_055_145);
  and2 I056_383(w_056_383, w_011_531, w_015_490);
  not1 I056_390(w_056_390, w_016_000);
  and2 I056_400(w_056_400, w_023_093, w_051_256);
  nand2 I056_412(w_056_412, w_001_009, w_047_299);
  and2 I056_427(w_056_427, w_013_059, w_030_015);
  and2 I056_434(w_056_434, w_017_073, w_035_043);
  or2  I056_438(w_056_438, w_045_361, w_040_480);
  or2  I056_457(w_056_457, w_017_386, w_020_408);
  or2  I056_462(w_056_462, w_029_071, w_054_415);
  and2 I056_463(w_056_463, w_047_307, w_049_095);
  and2 I056_465(w_056_465, w_047_205, w_024_059);
  nand2 I056_466(w_056_466, w_033_468, w_044_544);
  nand2 I056_476(w_056_476, w_024_215, w_036_117);
  nand2 I056_487(w_056_487, w_049_002, w_017_365);
  or2  I056_490(w_056_490, w_051_249, w_007_255);
  nand2 I056_491(w_056_491, w_031_546, w_012_087);
  not1 I056_493(w_056_493, w_027_060);
  and2 I056_499(w_056_499, w_008_222, w_050_435);
  or2  I056_500(w_056_500, w_010_768, w_048_016);
  or2  I056_501(w_056_501, w_041_038, w_007_126);
  and2 I056_505(w_056_505, w_035_035, w_035_093);
  not1 I056_507(w_056_507, w_040_196);
  nand2 I056_509(w_056_509, w_027_031, w_051_206);
  or2  I056_520(w_056_520, w_055_046, w_003_068);
  not1 I056_523(w_056_523, w_024_361);
  or2  I056_525(w_056_525, w_054_415, w_015_045);
  not1 I056_528(w_056_528, w_031_050);
  and2 I056_532(w_056_532, w_007_310, w_026_598);
  not1 I056_540(w_056_540, w_038_290);
  not1 I056_545(w_056_545, w_003_024);
  or2  I056_551(w_056_551, w_004_059, w_000_685);
  not1 I056_554(w_056_554, w_037_346);
  or2  I056_557(w_056_557, w_036_033, w_024_202);
  nand2 I056_567(w_056_567, w_046_608, w_024_433);
  and2 I056_579(w_056_579, w_001_011, w_055_290);
  and2 I056_586(w_056_586, w_021_097, w_012_207);
  nand2 I056_596(w_056_596, w_050_004, w_005_042);
  and2 I056_597(w_056_597, w_022_249, w_010_388);
  not1 I056_609(w_056_609, w_047_192);
  nand2 I056_610(w_056_610, w_052_037, w_015_347);
  not1 I056_615(w_056_615, w_043_026);
  or2  I056_620(w_056_620, w_027_056, w_000_053);
  and2 I056_622(w_056_622, w_003_063, w_021_182);
  not1 I056_623(w_056_623, w_014_088);
  nand2 I056_627(w_056_627, w_032_240, w_043_045);
  not1 I056_629(w_056_629, w_047_206);
  not1 I056_633(w_056_633, w_003_054);
  or2  I056_642(w_056_642, w_008_524, w_003_025);
  or2  I056_645(w_056_645, w_024_025, w_022_163);
  nand2 I056_655(w_056_655, w_028_131, w_025_297);
  not1 I056_661(w_056_661, w_017_318);
  not1 I056_663(w_056_663, w_002_390);
  and2 I056_665(w_056_665, w_039_515, w_012_050);
  nand2 I056_675(w_056_675, w_041_610, w_005_021);
  or2  I056_686(w_056_686, w_025_282, w_055_064);
  and2 I056_692(w_056_692, w_012_273, w_049_134);
  nand2 I056_702(w_056_702, w_030_339, w_020_408);
  or2  I056_703(w_056_703, w_040_210, w_050_259);
  not1 I056_709(w_056_709, w_007_127);
  and2 I056_710(w_056_710, w_051_027, w_029_080);
  not1 I056_713(w_056_713, w_026_132);
  and2 I056_721(w_056_721, w_020_023, w_044_041);
  and2 I056_723(w_056_723, w_043_028, w_044_577);
  not1 I056_724(w_056_724, w_004_170);
  and2 I056_736(w_056_736, w_016_003, w_029_039);
  or2  I057_000(w_057_000, w_029_080, w_038_044);
  or2  I057_001(w_057_001, w_053_096, w_033_517);
  or2  I057_002(w_057_002, w_021_108, w_017_461);
  nand2 I057_004(w_057_004, w_037_305, w_006_190);
  not1 I057_006(w_057_006, w_005_073);
  not1 I057_007(w_057_007, w_043_035);
  nand2 I057_008(w_057_008, w_039_024, w_042_191);
  and2 I057_010(w_057_010, w_013_411, w_017_640);
  and2 I057_013(w_057_013, w_050_593, w_027_065);
  and2 I057_018(w_057_018, w_026_098, w_031_382);
  or2  I057_019(w_057_019, w_012_055, w_029_061);
  and2 I057_022(w_057_022, w_050_136, w_013_178);
  not1 I057_023(w_057_023, w_038_606);
  and2 I057_025(w_057_025, w_046_211, w_030_367);
  or2  I057_028(w_057_028, w_049_294, w_042_275);
  nand2 I057_029(w_057_029, w_035_069, w_015_673);
  not1 I057_032(w_057_032, w_055_259);
  and2 I057_036(w_057_036, w_017_248, w_042_000);
  and2 I057_047(w_057_047, w_009_232, w_037_253);
  or2  I057_049(w_057_049, w_035_098, w_053_144);
  nand2 I057_052(w_057_052, w_020_177, w_023_135);
  not1 I057_053(w_057_053, w_056_721);
  not1 I057_055(w_057_055, w_028_147);
  not1 I057_056(w_057_056, w_041_083);
  and2 I057_057(w_057_057, w_004_214, w_012_298);
  or2  I057_058(w_057_058, w_048_011, w_034_042);
  nand2 I057_060(w_057_060, w_022_227, w_055_154);
  and2 I057_061(w_057_061, w_020_136, w_002_285);
  nand2 I057_062(w_057_062, w_031_571, w_050_012);
  not1 I057_063(w_057_063, w_042_062);
  not1 I057_066(w_057_066, w_002_370);
  nand2 I057_068(w_057_068, w_005_254, w_010_412);
  and2 I057_070(w_057_070, w_050_309, w_052_006);
  and2 I057_073(w_057_073, w_034_012, w_012_101);
  not1 I057_076(w_057_076, w_022_313);
  not1 I057_078(w_057_078, w_049_131);
  nand2 I057_081(w_057_081, w_012_167, w_017_024);
  nand2 I057_082(w_057_082, w_028_110, w_020_247);
  and2 I057_083(w_057_083, w_001_001, w_050_612);
  nand2 I057_084(w_057_084, w_033_541, w_052_017);
  and2 I057_085(w_057_085, w_007_096, w_006_066);
  and2 I057_086(w_057_086, w_039_348, w_013_320);
  and2 I057_087(w_057_087, w_030_413, w_024_426);
  and2 I057_088(w_057_088, w_000_462, w_052_042);
  or2  I057_092(w_057_092, w_056_123, w_053_070);
  nand2 I057_094(w_057_094, w_023_100, w_043_014);
  and2 I057_095(w_057_095, w_022_117, w_044_029);
  not1 I057_097(w_057_097, w_018_013);
  nand2 I057_099(w_057_099, w_025_060, w_008_239);
  nand2 I057_100(w_057_100, w_031_531, w_008_252);
  not1 I057_101(w_057_101, w_052_042);
  not1 I057_102(w_057_102, w_033_159);
  not1 I057_105(w_057_105, w_052_044);
  not1 I057_107(w_057_107, w_018_041);
  or2  I057_112(w_057_112, w_011_239, w_045_043);
  nand2 I057_114(w_057_114, w_038_317, w_023_047);
  or2  I057_117(w_057_117, w_003_029, w_050_373);
  and2 I057_121(w_057_121, w_045_170, w_001_007);
  not1 I057_123(w_057_123, w_042_041);
  and2 I057_124(w_057_124, w_035_126, w_017_257);
  not1 I057_126(w_057_126, w_031_442);
  and2 I057_131(w_057_131, w_050_101, w_039_063);
  and2 I057_135(w_057_135, w_052_011, w_040_583);
  not1 I057_137(w_057_137, w_028_058);
  nand2 I057_140(w_057_140, w_050_058, w_047_454);
  nand2 I057_141(w_057_141, w_042_026, w_023_079);
  not1 I057_143(w_057_143, w_024_181);
  nand2 I057_144(w_057_144, w_007_316, w_030_417);
  or2  I057_145(w_057_145, w_022_048, w_001_029);
  or2  I057_146(w_057_146, w_030_143, w_047_219);
  not1 I057_147(w_057_147, w_040_147);
  not1 I057_150(w_057_150, w_016_002);
  not1 I057_155(w_057_155, w_008_469);
  not1 I057_156(w_057_156, w_010_003);
  nand2 I057_160(w_057_160, w_052_015, w_033_710);
  or2  I057_171(w_057_171, w_012_205, w_040_039);
  and2 I057_174(w_057_174, w_050_407, w_031_553);
  or2  I057_175(w_057_175, w_027_018, w_038_489);
  nand2 I057_182(w_057_182, w_015_579, w_012_019);
  nand2 I057_185(w_057_185, w_039_658, w_010_640);
  not1 I057_187(w_057_187, w_022_142);
  and2 I057_194(w_057_194, w_009_239, w_011_458);
  and2 I057_200(w_057_200, w_012_327, w_040_070);
  and2 I057_203(w_057_203, w_049_124, w_013_391);
  not1 I057_210(w_057_210, w_025_241);
  or2  I057_213(w_057_213, w_024_292, w_008_713);
  and2 I057_215(w_057_215, w_006_016, w_016_002);
  nand2 I057_220(w_057_220, w_051_094, w_026_614);
  nand2 I057_228(w_057_228, w_013_165, w_044_180);
  nand2 I057_229(w_057_229, w_033_722, w_038_469);
  and2 I057_230(w_057_230, w_010_417, w_032_499);
  nand2 I057_235(w_057_235, w_018_019, w_034_073);
  and2 I057_236(w_057_236, w_034_006, w_035_066);
  or2  I057_237(w_057_237, w_002_572, w_009_094);
  and2 I057_239(w_057_239, w_044_058, w_044_402);
  or2  I057_241(w_057_241, w_015_527, w_049_335);
  nand2 I057_243(w_057_243, w_019_004, w_016_005);
  nand2 I057_246(w_057_246, w_035_056, w_018_027);
  or2  I057_250(w_057_250, w_049_172, w_047_360);
  nand2 I057_254(w_057_254, w_034_002, w_024_507);
  or2  I057_257(w_057_257, w_045_069, w_029_101);
  nand2 I057_258(w_057_258, w_028_107, w_021_099);
  and2 I057_262(w_057_262, w_014_280, w_044_424);
  or2  I057_268(w_057_268, w_001_021, w_033_638);
  or2  I057_271(w_057_271, w_001_004, w_011_618);
  or2  I057_273(w_057_273, w_029_113, w_044_611);
  not1 I057_274(w_057_274, w_042_013);
  not1 I057_279(w_057_279, w_005_108);
  nand2 I057_281(w_057_281, w_044_014, w_017_512);
  and2 I057_285(w_057_285, w_003_012, w_000_285);
  not1 I057_289(w_057_289, w_054_569);
  and2 I057_291(w_057_291, w_035_066, w_039_406);
  nand2 I057_293(w_057_293, w_056_232, w_004_000);
  not1 I057_296(w_057_296, w_035_102);
  and2 I057_307(w_057_307, w_050_056, w_048_004);
  not1 I057_313(w_057_313, w_019_015);
  not1 I058_005(w_058_005, w_025_028);
  nand2 I058_017(w_058_017, w_020_186, w_010_341);
  or2  I058_022(w_058_022, w_026_283, w_050_461);
  and2 I058_025(w_058_025, w_045_333, w_011_556);
  or2  I058_029(w_058_029, w_042_323, w_042_045);
  and2 I058_030(w_058_030, w_042_255, w_025_187);
  and2 I058_032(w_058_032, w_016_001, w_027_053);
  and2 I058_033(w_058_033, w_014_027, w_018_004);
  not1 I058_037(w_058_037, w_008_100);
  or2  I058_050(w_058_050, w_027_162, w_055_307);
  nand2 I058_056(w_058_056, w_053_140, w_000_030);
  not1 I058_060(w_058_060, w_057_200);
  and2 I058_061(w_058_061, w_018_011, w_033_569);
  not1 I058_065(w_058_065, w_009_134);
  nand2 I058_070(w_058_070, w_049_166, w_015_056);
  or2  I058_073(w_058_073, w_021_078, w_051_052);
  nand2 I058_074(w_058_074, w_004_218, w_049_119);
  or2  I058_075(w_058_075, w_049_029, w_051_062);
  or2  I058_081(w_058_081, w_001_032, w_006_205);
  nand2 I058_082(w_058_082, w_048_011, w_005_136);
  nand2 I058_085(w_058_085, w_008_539, w_056_487);
  nand2 I058_086(w_058_086, w_002_086, w_017_112);
  and2 I058_088(w_058_088, w_027_173, w_019_007);
  nand2 I058_090(w_058_090, w_012_264, w_053_060);
  or2  I058_092(w_058_092, w_055_286, w_020_412);
  nand2 I058_095(w_058_095, w_023_147, w_040_311);
  or2  I058_104(w_058_104, w_004_125, w_000_768);
  and2 I058_105(w_058_105, w_042_144, w_038_151);
  not1 I058_111(w_058_111, w_023_102);
  not1 I058_112(w_058_112, w_057_150);
  and2 I058_119(w_058_119, w_028_456, w_029_109);
  nand2 I058_123(w_058_123, w_003_079, w_036_283);
  not1 I058_132(w_058_132, w_023_033);
  not1 I058_134(w_058_134, w_010_263);
  nand2 I058_135(w_058_135, w_050_119, w_030_312);
  nand2 I058_136(w_058_136, w_001_022, w_029_001);
  not1 I058_140(w_058_140, w_014_129);
  or2  I058_148(w_058_148, w_044_331, w_019_002);
  or2  I058_156(w_058_156, w_048_001, w_029_111);
  not1 I058_159(w_058_159, w_022_272);
  or2  I058_161(w_058_161, w_026_145, w_022_357);
  and2 I058_162(w_058_162, w_052_014, w_041_079);
  or2  I058_164(w_058_164, w_015_151, w_036_177);
  nand2 I058_171(w_058_171, w_024_049, w_047_185);
  nand2 I058_174(w_058_174, w_046_172, w_040_219);
  not1 I058_179(w_058_179, w_009_094);
  nand2 I058_182(w_058_182, w_018_037, w_008_704);
  not1 I058_193(w_058_193, w_012_050);
  or2  I058_195(w_058_195, w_056_106, w_023_105);
  not1 I058_206(w_058_206, w_022_102);
  or2  I058_208(w_058_208, w_028_392, w_033_208);
  and2 I058_210(w_058_210, w_021_255, w_055_068);
  and2 I058_216(w_058_216, w_047_033, w_013_059);
  not1 I058_224(w_058_224, w_017_309);
  and2 I058_229(w_058_229, w_054_463, w_035_083);
  nand2 I058_235(w_058_235, w_012_130, w_044_449);
  nand2 I058_238(w_058_238, w_026_591, w_019_004);
  and2 I058_251(w_058_251, w_019_012, w_016_008);
  and2 I058_253(w_058_253, w_037_267, w_053_154);
  or2  I058_254(w_058_254, w_055_165, w_005_112);
  and2 I058_255(w_058_255, w_016_008, w_036_128);
  not1 I058_256(w_058_256, w_001_017);
  not1 I058_258(w_058_258, w_044_322);
  not1 I058_271(w_058_271, w_037_266);
  or2  I058_274(w_058_274, w_027_155, w_042_368);
  or2  I058_280(w_058_280, w_045_359, w_020_347);
  not1 I058_282(w_058_282, w_039_681);
  and2 I058_287(w_058_287, w_031_125, w_052_029);
  and2 I058_292(w_058_292, w_047_394, w_050_238);
  nand2 I058_295(w_058_295, w_026_643, w_027_075);
  not1 I058_304(w_058_304, w_024_399);
  nand2 I058_306(w_058_306, w_036_026, w_041_024);
  not1 I058_310(w_058_310, w_024_276);
  and2 I058_316(w_058_316, w_013_392, w_013_146);
  or2  I058_321(w_058_321, w_020_122, w_024_392);
  or2  I058_327(w_058_327, w_041_013, w_004_459);
  and2 I058_330(w_058_330, w_048_019, w_027_053);
  not1 I058_332(w_058_332, w_003_031);
  and2 I058_335(w_058_335, w_022_030, w_046_248);
  not1 I058_341(w_058_341, w_001_028);
  and2 I058_344(w_058_344, w_006_015, w_008_055);
  or2  I058_352(w_058_352, w_007_431, w_012_153);
  and2 I058_359(w_058_359, w_025_118, w_039_713);
  and2 I058_366(w_058_366, w_024_211, w_001_009);
  or2  I058_368(w_058_368, w_009_498, w_055_064);
  nand2 I058_376(w_058_376, w_010_415, w_006_222);
  not1 I058_379(w_058_379, w_054_284);
  and2 I058_383(w_058_383, w_039_440, w_049_305);
  or2  I058_402(w_058_402, w_023_041, w_043_005);
  and2 I058_404(w_058_404, w_028_178, w_000_704);
  not1 I058_416(w_058_416, w_020_092);
  not1 I058_420(w_058_420, w_014_137);
  or2  I058_423(w_058_423, w_046_132, w_032_444);
  or2  I058_425(w_058_425, w_033_646, w_042_220);
  nand2 I058_427(w_058_427, w_000_227, w_045_003);
  or2  I058_428(w_058_428, w_038_200, w_037_285);
  and2 I058_442(w_058_442, w_052_036, w_035_013);
  nand2 I058_447(w_058_447, w_055_131, w_055_183);
  or2  I058_453(w_058_453, w_025_102, w_018_009);
  nand2 I058_454(w_058_454, w_015_038, w_054_078);
  and2 I058_457(w_058_457, w_036_201, w_041_090);
  or2  I058_459(w_058_459, w_038_134, w_010_515);
  and2 I058_467(w_058_467, w_042_095, w_009_134);
  or2  I058_469(w_058_469, w_045_047, w_021_267);
  or2  I058_472(w_058_472, w_050_543, w_038_173);
  or2  I058_477(w_058_477, w_057_174, w_010_000);
  not1 I058_478(w_058_478, w_028_137);
  and2 I058_479(w_058_479, w_014_074, w_008_701);
  not1 I058_484(w_058_484, w_046_042);
  or2  I058_485(w_058_485, w_011_520, w_026_163);
  nand2 I058_493(w_058_493, w_038_317, w_052_021);
  or2  I058_498(w_058_498, w_032_442, w_039_046);
  not1 I058_503(w_058_503, w_042_428);
  and2 I058_504(w_058_504, w_023_198, w_015_163);
  nand2 I058_505(w_058_505, w_039_606, w_005_292);
  not1 I058_513(w_058_513, w_008_337);
  nand2 I058_515(w_058_515, w_053_135, w_037_245);
  nand2 I058_522(w_058_522, w_007_371, w_046_292);
  nand2 I058_527(w_058_527, w_052_008, w_010_369);
  and2 I058_534(w_058_534, w_001_025, w_018_018);
  nand2 I058_536(w_058_536, w_007_139, w_001_005);
  nand2 I058_538(w_058_538, w_054_283, w_029_023);
  or2  I058_540(w_058_540, w_048_015, w_011_004);
  or2  I058_541(w_058_541, w_041_429, w_022_185);
  not1 I058_550(w_058_550, w_016_004);
  not1 I058_555(w_058_555, w_033_291);
  nand2 I058_559(w_058_559, w_053_062, w_020_033);
  not1 I058_562(w_058_562, w_057_156);
  and2 I058_568(w_058_568, w_014_021, w_045_323);
  or2  I058_570(w_058_570, w_056_008, w_042_116);
  not1 I058_581(w_058_581, w_035_100);
  nand2 I058_589(w_058_589, w_025_044, w_009_216);
  or2  I058_590(w_058_590, w_017_133, w_043_015);
  not1 I058_593(w_058_593, w_011_075);
  or2  I058_594(w_058_594, w_054_581, w_027_020);
  and2 I058_596(w_058_596, w_010_060, w_055_287);
  not1 I058_597(w_058_597, w_032_526);
  and2 I058_602(w_058_602, w_005_042, w_028_489);
  and2 I058_607(w_058_607, w_037_095, w_031_213);
  and2 I058_635(w_058_635, w_017_071, w_038_447);
  nand2 I058_638(w_058_638, w_026_539, w_040_099);
  nand2 I058_645(w_058_645, w_026_105, w_032_187);
  not1 I058_647(w_058_647, w_015_287);
  not1 I058_655(w_058_655, w_039_719);
  not1 I058_656(w_058_656, w_010_417);
  nand2 I058_658(w_058_658, w_042_158, w_038_315);
  nand2 I058_660(w_058_660, w_048_012, w_020_138);
  not1 I058_664(w_058_664, w_046_129);
  not1 I058_673(w_058_673, w_008_553);
  not1 I058_681(w_058_681, w_036_033);
  not1 I058_683(w_058_683, w_015_246);
  nand2 I058_696(w_058_696, w_034_009, w_045_050);
  nand2 I058_699(w_058_699, w_053_120, w_007_032);
  nand2 I059_001(w_059_001, w_057_237, w_034_016);
  not1 I059_002(w_059_002, w_020_610);
  or2  I059_003(w_059_003, w_017_068, w_029_009);
  nand2 I059_005(w_059_005, w_007_357, w_008_441);
  nand2 I059_012(w_059_012, w_026_681, w_018_015);
  or2  I059_017(w_059_017, w_045_074, w_007_160);
  nand2 I059_026(w_059_026, w_020_004, w_028_077);
  or2  I059_029(w_059_029, w_015_045, w_007_172);
  or2  I059_032(w_059_032, w_007_167, w_029_080);
  and2 I059_043(w_059_043, w_026_257, w_002_018);
  not1 I059_045(w_059_045, w_003_001);
  or2  I059_049(w_059_049, w_021_139, w_019_002);
  and2 I059_052(w_059_052, w_017_657, w_013_043);
  or2  I059_055(w_059_055, w_046_571, w_029_074);
  and2 I059_056(w_059_056, w_046_606, w_040_644);
  or2  I059_057(w_059_057, w_040_582, w_034_057);
  or2  I059_060(w_059_060, w_032_243, w_008_515);
  or2  I059_061(w_059_061, w_009_030, w_010_442);
  not1 I059_066(w_059_066, w_027_160);
  not1 I059_084(w_059_084, w_053_050);
  nand2 I059_089(w_059_089, w_058_295, w_010_134);
  and2 I059_090(w_059_090, w_010_712, w_022_135);
  or2  I059_094(w_059_094, w_049_341, w_054_472);
  or2  I059_101(w_059_101, w_020_484, w_006_032);
  or2  I059_103(w_059_103, w_018_023, w_006_025);
  and2 I059_111(w_059_111, w_032_389, w_053_013);
  not1 I059_114(w_059_114, w_001_034);
  and2 I059_125(w_059_125, w_055_204, w_049_023);
  not1 I059_131(w_059_131, w_045_106);
  nand2 I059_135(w_059_135, w_053_020, w_056_224);
  not1 I059_140(w_059_140, w_034_007);
  or2  I059_146(w_059_146, w_019_015, w_018_019);
  not1 I059_147(w_059_147, w_056_709);
  and2 I059_150(w_059_150, w_034_035, w_010_365);
  not1 I059_157(w_059_157, w_048_003);
  nand2 I059_159(w_059_159, w_000_418, w_037_087);
  and2 I059_162(w_059_162, w_023_051, w_057_143);
  not1 I059_165(w_059_165, w_008_013);
  and2 I059_166(w_059_166, w_049_101, w_021_204);
  not1 I059_167(w_059_167, w_049_294);
  not1 I059_168(w_059_168, w_012_162);
  not1 I059_170(w_059_170, w_025_101);
  not1 I059_173(w_059_173, w_035_043);
  nand2 I059_174(w_059_174, w_028_175, w_048_002);
  not1 I059_178(w_059_178, w_001_031);
  or2  I059_181(w_059_181, w_007_007, w_051_051);
  and2 I059_183(w_059_183, w_000_379, w_058_032);
  or2  I059_184(w_059_184, w_002_545, w_047_073);
  and2 I059_186(w_059_186, w_012_171, w_031_097);
  or2  I059_196(w_059_196, w_013_020, w_042_006);
  or2  I059_200(w_059_200, w_045_327, w_051_308);
  not1 I059_201(w_059_201, w_021_217);
  not1 I059_202(w_059_202, w_020_119);
  and2 I059_209(w_059_209, w_056_724, w_044_195);
  nand2 I059_213(w_059_213, w_044_608, w_044_040);
  and2 I059_218(w_059_218, w_012_277, w_003_059);
  nand2 I059_220(w_059_220, w_002_434, w_033_114);
  and2 I059_233(w_059_233, w_035_063, w_007_138);
  nand2 I059_236(w_059_236, w_042_307, w_056_141);
  and2 I059_239(w_059_239, w_017_360, w_027_179);
  or2  I059_242(w_059_242, w_020_607, w_011_147);
  or2  I059_248(w_059_248, w_005_115, w_019_003);
  or2  I059_249(w_059_249, w_030_080, w_028_132);
  not1 I059_255(w_059_255, w_005_092);
  nand2 I059_258(w_059_258, w_012_262, w_040_442);
  not1 I059_260(w_059_260, w_009_122);
  and2 I059_278(w_059_278, w_011_121, w_014_136);
  or2  I059_286(w_059_286, w_031_440, w_030_284);
  not1 I059_288(w_059_288, w_039_148);
  nand2 I059_301(w_059_301, w_022_151, w_010_222);
  not1 I059_309(w_059_309, w_015_001);
  or2  I059_313(w_059_313, w_036_376, w_026_002);
  nand2 I059_315(w_059_315, w_021_013, w_011_407);
  and2 I059_321(w_059_321, w_025_072, w_008_763);
  or2  I059_328(w_059_328, w_055_180, w_017_664);
  and2 I059_337(w_059_337, w_017_206, w_022_050);
  and2 I059_340(w_059_340, w_000_496, w_036_120);
  not1 I059_348(w_059_348, w_055_133);
  or2  I059_354(w_059_354, w_009_388, w_055_042);
  or2  I059_355(w_059_355, w_016_002, w_010_319);
  not1 I059_364(w_059_364, w_041_432);
  nand2 I059_392(w_059_392, w_019_009, w_036_154);
  and2 I059_396(w_059_396, w_046_562, w_000_083);
  not1 I059_405(w_059_405, w_039_676);
  and2 I059_413(w_059_413, w_012_188, w_019_010);
  and2 I059_423(w_059_423, w_053_029, w_045_210);
  not1 I059_425(w_059_425, w_048_011);
  and2 I059_430(w_059_430, w_019_011, w_051_323);
  nand2 I059_431(w_059_431, w_044_395, w_047_340);
  not1 I059_432(w_059_432, w_036_243);
  and2 I059_439(w_059_439, w_040_325, w_051_232);
  not1 I059_444(w_059_444, w_058_515);
  nand2 I059_455(w_059_455, w_051_181, w_019_012);
  nand2 I059_459(w_059_459, w_058_541, w_005_103);
  or2  I059_462(w_059_462, w_008_115, w_050_234);
  not1 I059_479(w_059_479, w_002_225);
  or2  I059_482(w_059_482, w_012_315, w_017_141);
  or2  I059_489(w_059_489, w_048_015, w_047_105);
  nand2 I059_500(w_059_500, w_021_094, w_008_264);
  nand2 I059_501(w_059_501, w_020_193, w_015_257);
  or2  I059_507(w_059_507, w_028_122, w_024_143);
  and2 I059_508(w_059_508, w_048_008, w_013_186);
  or2  I059_512(w_059_512, w_032_067, w_032_275);
  nand2 I059_517(w_059_517, w_022_243, w_028_228);
  or2  I059_521(w_059_521, w_041_548, w_004_492);
  nand2 I059_522(w_059_522, w_027_014, w_017_122);
  and2 I059_533(w_059_533, w_045_291, w_052_031);
  nand2 I059_538(w_059_538, w_019_014, w_024_166);
  nand2 I059_550(w_059_550, w_037_124, w_003_084);
  nand2 I059_552(w_059_552, w_052_033, w_054_466);
  and2 I059_553(w_059_553, w_010_236, w_030_086);
  nand2 I059_554(w_059_554, w_025_177, w_018_021);
  and2 I059_555(w_059_555, w_000_713, w_012_183);
  not1 I059_559(w_059_559, w_053_001);
  nand2 I059_567(w_059_567, w_014_151, w_030_119);
  nand2 I059_578(w_059_578, w_028_335, w_009_532);
  or2  I059_587(w_059_587, w_052_039, w_046_686);
  not1 I059_588(w_059_588, w_057_032);
  not1 I059_589(w_059_589, w_052_033);
  or2  I059_596(w_059_596, w_023_108, w_015_371);
  or2  I059_600(w_059_600, w_013_436, w_046_647);
  or2  I059_612(w_059_612, w_038_087, w_044_206);
  nand2 I059_616(w_059_616, w_032_462, w_002_642);
  nand2 I059_633(w_059_633, w_028_231, w_035_070);
  not1 I059_636(w_059_636, w_043_025);
  and2 I059_637(w_059_637, w_009_160, w_045_265);
  nand2 I059_639(w_059_639, w_039_367, w_040_558);
  and2 I059_647(w_059_647, w_018_042, w_027_014);
  and2 I059_660(w_059_660, w_016_000, w_049_120);
  and2 I059_667(w_059_667, w_049_021, w_013_137);
  nand2 I059_683(w_059_683, w_035_062, w_023_027);
  and2 I059_695(w_059_695, w_009_520, w_041_397);
  or2  I059_698(w_059_698, w_001_012, w_044_673);
  and2 I059_702(w_059_702, w_005_190, w_029_042);
  not1 I059_708(w_059_708, w_052_032);
  and2 I059_722(w_059_722, w_023_100, w_051_337);
  not1 I059_724(w_059_724, w_022_281);
  not1 I059_727(w_059_727, w_036_087);
  or2  I059_730(w_059_730, w_032_490, w_057_274);
  not1 I059_734(w_059_734, w_053_153);
  not1 I060_003(w_060_003, w_052_007);
  or2  I060_009(w_060_009, w_020_076, w_027_153);
  and2 I060_012(w_060_012, w_041_604, w_051_003);
  or2  I060_016(w_060_016, w_053_103, w_048_008);
  nand2 I060_017(w_060_017, w_051_095, w_038_068);
  or2  I060_019(w_060_019, w_009_568, w_054_095);
  nand2 I060_020(w_060_020, w_014_197, w_006_019);
  nand2 I060_024(w_060_024, w_053_004, w_052_002);
  and2 I060_025(w_060_025, w_034_024, w_045_226);
  and2 I060_026(w_060_026, w_039_010, w_003_028);
  or2  I060_027(w_060_027, w_001_013, w_037_071);
  not1 I060_030(w_060_030, w_046_246);
  and2 I060_033(w_060_033, w_054_169, w_016_005);
  not1 I060_036(w_060_036, w_034_013);
  or2  I060_037(w_060_037, w_036_118, w_013_479);
  not1 I060_038(w_060_038, w_051_021);
  or2  I060_039(w_060_039, w_015_315, w_019_005);
  or2  I060_045(w_060_045, w_008_009, w_036_297);
  not1 I060_049(w_060_049, w_023_066);
  nand2 I060_050(w_060_050, w_020_255, w_052_015);
  not1 I060_053(w_060_053, w_042_152);
  or2  I060_058(w_060_058, w_056_528, w_025_000);
  nand2 I060_071(w_060_071, w_008_709, w_052_045);
  or2  I060_073(w_060_073, w_050_306, w_031_213);
  or2  I060_075(w_060_075, w_017_228, w_031_561);
  and2 I060_080(w_060_080, w_023_063, w_016_000);
  and2 I060_081(w_060_081, w_055_007, w_058_344);
  nand2 I060_085(w_060_085, w_009_562, w_021_146);
  not1 I060_086(w_060_086, w_053_015);
  or2  I060_088(w_060_088, w_041_052, w_024_223);
  nand2 I060_097(w_060_097, w_035_115, w_052_036);
  nand2 I060_098(w_060_098, w_027_158, w_041_288);
  nand2 I060_109(w_060_109, w_045_148, w_057_146);
  nand2 I060_112(w_060_112, w_054_043, w_011_280);
  or2  I060_114(w_060_114, w_023_007, w_047_283);
  not1 I060_116(w_060_116, w_044_181);
  or2  I060_118(w_060_118, w_057_293, w_001_035);
  and2 I060_119(w_060_119, w_047_350, w_052_033);
  or2  I060_122(w_060_122, w_033_748, w_051_322);
  or2  I060_123(w_060_123, w_038_024, w_015_434);
  and2 I060_125(w_060_125, w_025_187, w_030_409);
  and2 I060_126(w_060_126, w_048_001, w_018_029);
  nand2 I060_131(w_060_131, w_011_270, w_059_301);
  or2  I060_141(w_060_141, w_045_130, w_003_000);
  or2  I060_148(w_060_148, w_043_010, w_050_493);
  and2 I060_155(w_060_155, w_057_281, w_021_112);
  not1 I060_160(w_060_160, w_035_122);
  nand2 I060_161(w_060_161, w_039_051, w_010_589);
  or2  I060_164(w_060_164, w_041_581, w_039_014);
  and2 I060_167(w_060_167, w_024_055, w_019_010);
  nand2 I060_168(w_060_168, w_021_150, w_005_134);
  not1 I060_169(w_060_169, w_020_394);
  not1 I060_171(w_060_171, w_034_026);
  nand2 I060_176(w_060_176, w_019_019, w_051_013);
  or2  I060_189(w_060_189, w_016_005, w_025_050);
  or2  I060_190(w_060_190, w_035_073, w_023_007);
  not1 I060_194(w_060_194, w_053_083);
  not1 I060_198(w_060_198, w_049_278);
  and2 I060_204(w_060_204, w_055_240, w_005_100);
  nand2 I060_208(w_060_208, w_006_217, w_032_124);
  not1 I060_209(w_060_209, w_002_361);
  or2  I060_212(w_060_212, w_041_497, w_050_386);
  or2  I060_216(w_060_216, w_042_203, w_057_230);
  not1 I060_222(w_060_222, w_002_391);
  or2  I060_224(w_060_224, w_028_142, w_013_286);
  or2  I060_225(w_060_225, w_052_022, w_039_413);
  not1 I060_246(w_060_246, w_008_094);
  or2  I060_254(w_060_254, w_001_025, w_051_343);
  and2 I060_257(w_060_257, w_014_127, w_046_297);
  nand2 I060_259(w_060_259, w_005_206, w_044_225);
  nand2 I060_261(w_060_261, w_026_506, w_012_040);
  not1 I060_262(w_060_262, w_010_233);
  or2  I060_265(w_060_265, w_008_437, w_009_314);
  or2  I060_266(w_060_266, w_006_072, w_053_007);
  nand2 I060_268(w_060_268, w_050_348, w_007_119);
  or2  I060_272(w_060_272, w_030_162, w_022_276);
  nand2 I060_277(w_060_277, w_017_025, w_048_010);
  or2  I060_278(w_060_278, w_047_254, w_018_015);
  not1 I060_284(w_060_284, w_043_026);
  not1 I060_285(w_060_285, w_045_407);
  not1 I060_288(w_060_288, w_012_337);
  not1 I060_289(w_060_289, w_051_052);
  nand2 I060_290(w_060_290, w_021_200, w_006_035);
  nand2 I060_291(w_060_291, w_033_014, w_056_491);
  nand2 I060_294(w_060_294, w_027_113, w_034_005);
  or2  I060_296(w_060_296, w_008_524, w_049_065);
  and2 I060_299(w_060_299, w_007_204, w_039_372);
  nand2 I060_300(w_060_300, w_045_161, w_014_028);
  not1 I060_305(w_060_305, w_033_216);
  nand2 I060_308(w_060_308, w_034_039, w_036_161);
  not1 I060_310(w_060_310, w_021_155);
  not1 I060_313(w_060_313, w_033_312);
  not1 I060_323(w_060_323, w_053_094);
  not1 I060_324(w_060_324, w_045_189);
  nand2 I060_326(w_060_326, w_037_308, w_010_125);
  not1 I060_330(w_060_330, w_037_211);
  or2  I060_331(w_060_331, w_014_009, w_001_023);
  or2  I060_332(w_060_332, w_001_019, w_004_059);
  not1 I060_333(w_060_333, w_006_030);
  or2  I060_336(w_060_336, w_000_574, w_050_621);
  nand2 I060_338(w_060_338, w_047_148, w_042_332);
  and2 I060_341(w_060_341, w_050_199, w_019_004);
  and2 I060_343(w_060_343, w_023_095, w_003_011);
  not1 I060_344(w_060_344, w_019_019);
  and2 I060_354(w_060_354, w_020_590, w_011_152);
  not1 I060_355(w_060_355, w_019_009);
  and2 I060_359(w_060_359, w_007_274, w_028_251);
  not1 I060_365(w_060_365, w_003_083);
  or2  I060_366(w_060_366, w_026_343, w_012_163);
  not1 I060_372(w_060_372, w_034_007);
  and2 I060_381(w_060_381, w_021_196, w_056_224);
  nand2 I060_387(w_060_387, w_059_045, w_048_009);
  or2  I060_395(w_060_395, w_040_409, w_055_164);
  and2 I061_002(w_061_002, w_043_035, w_006_115);
  not1 I061_003(w_061_003, w_027_202);
  nand2 I061_004(w_061_004, w_056_615, w_045_390);
  nand2 I061_005(w_061_005, w_011_131, w_036_229);
  not1 I061_012(w_061_012, w_018_031);
  or2  I061_023(w_061_023, w_052_005, w_058_148);
  not1 I061_027(w_061_027, w_057_022);
  nand2 I061_028(w_061_028, w_009_101, w_048_016);
  and2 I061_029(w_061_029, w_036_318, w_044_021);
  nand2 I061_033(w_061_033, w_040_327, w_034_032);
  nand2 I061_042(w_061_042, w_053_101, w_032_089);
  or2  I061_046(w_061_046, w_053_144, w_013_428);
  nand2 I061_047(w_061_047, w_028_089, w_058_638);
  and2 I061_050(w_061_050, w_044_403, w_027_071);
  not1 I061_051(w_061_051, w_043_023);
  nand2 I061_052(w_061_052, w_035_001, w_028_098);
  and2 I061_056(w_061_056, w_040_554, w_051_225);
  nand2 I061_057(w_061_057, w_036_180, w_022_053);
  nand2 I061_058(w_061_058, w_006_009, w_030_330);
  nand2 I061_059(w_061_059, w_058_428, w_009_301);
  nand2 I061_061(w_061_061, w_048_014, w_026_684);
  nand2 I061_062(w_061_062, w_036_261, w_060_272);
  not1 I061_063(w_061_063, w_052_029);
  or2  I061_064(w_061_064, w_029_042, w_003_011);
  nand2 I061_065(w_061_065, w_010_711, w_033_231);
  not1 I061_066(w_061_066, w_032_211);
  or2  I061_073(w_061_073, w_012_267, w_009_302);
  or2  I061_082(w_061_082, w_018_006, w_060_088);
  or2  I061_084(w_061_084, w_009_493, w_031_148);
  not1 I061_088(w_061_088, w_030_372);
  nand2 I061_089(w_061_089, w_035_068, w_051_107);
  and2 I061_099(w_061_099, w_033_605, w_045_181);
  and2 I061_100(w_061_100, w_046_096, w_048_012);
  nand2 I061_101(w_061_101, w_058_033, w_003_060);
  nand2 I061_103(w_061_103, w_007_054, w_035_095);
  nand2 I061_105(w_061_105, w_047_201, w_033_711);
  or2  I061_106(w_061_106, w_005_068, w_039_395);
  nand2 I061_122(w_061_122, w_021_249, w_028_326);
  not1 I061_123(w_061_123, w_005_182);
  and2 I061_125(w_061_125, w_021_007, w_059_103);
  and2 I061_126(w_061_126, w_028_197, w_053_089);
  not1 I061_142(w_061_142, w_001_010);
  not1 I061_143(w_061_143, w_021_082);
  or2  I061_146(w_061_146, w_059_727, w_020_181);
  and2 I061_147(w_061_147, w_050_630, w_002_458);
  not1 I061_148(w_061_148, w_031_162);
  nand2 I061_157(w_061_157, w_014_016, w_013_546);
  nand2 I061_158(w_061_158, w_013_049, w_059_233);
  and2 I061_160(w_061_160, w_060_332, w_053_067);
  not1 I061_161(w_061_161, w_020_110);
  or2  I061_162(w_061_162, w_052_019, w_028_097);
  not1 I061_168(w_061_168, w_043_042);
  not1 I061_172(w_061_172, w_029_067);
  not1 I061_175(w_061_175, w_012_019);
  or2  I061_178(w_061_178, w_038_061, w_017_293);
  not1 I061_179(w_061_179, w_008_212);
  nand2 I061_182(w_061_182, w_009_513, w_031_557);
  and2 I061_184(w_061_184, w_042_252, w_004_486);
  or2  I061_188(w_061_188, w_056_532, w_035_118);
  not1 I061_192(w_061_192, w_012_235);
  nand2 I061_194(w_061_194, w_031_083, w_023_035);
  or2  I061_196(w_061_196, w_046_099, w_019_013);
  or2  I061_198(w_061_198, w_045_205, w_051_369);
  not1 I061_199(w_061_199, w_060_338);
  not1 I061_200(w_061_200, w_040_071);
  and2 I061_205(w_061_205, w_004_402, w_028_464);
  or2  I061_213(w_061_213, w_033_057, w_025_042);
  and2 I061_217(w_061_217, w_011_564, w_018_008);
  and2 I061_219(w_061_219, w_056_172, w_015_118);
  not1 I061_221(w_061_221, w_027_125);
  and2 I061_227(w_061_227, w_004_159, w_037_130);
  nand2 I061_230(w_061_230, w_006_183, w_024_068);
  or2  I061_240(w_061_240, w_020_167, w_023_137);
  or2  I061_241(w_061_241, w_055_076, w_035_056);
  not1 I061_242(w_061_242, w_028_038);
  nand2 I061_253(w_061_253, w_004_291, w_047_214);
  not1 I061_255(w_061_255, w_042_036);
  or2  I061_256(w_061_256, w_003_025, w_026_453);
  nand2 I061_257(w_061_257, w_040_065, w_028_483);
  not1 I061_260(w_061_260, w_060_141);
  not1 I061_264(w_061_264, w_058_635);
  nand2 I061_266(w_061_266, w_004_204, w_021_248);
  nand2 I061_270(w_061_270, w_009_032, w_003_036);
  and2 I061_271(w_061_271, w_003_053, w_001_035);
  nand2 I061_276(w_061_276, w_000_147, w_056_049);
  nand2 I061_277(w_061_277, w_048_000, w_019_019);
  nand2 I061_283(w_061_283, w_028_543, w_006_165);
  nand2 I061_285(w_061_285, w_051_210, w_027_131);
  not1 I061_287(w_061_287, w_031_026);
  not1 I061_294(w_061_294, w_004_138);
  not1 I061_296(w_061_296, w_036_404);
  not1 I061_298(w_061_298, w_003_044);
  not1 I061_300(w_061_300, w_009_116);
  and2 I061_301(w_061_301, w_045_242, w_047_267);
  not1 I061_302(w_061_302, w_016_000);
  and2 I061_305(w_061_305, w_042_304, w_026_058);
  nand2 I061_306(w_061_306, w_039_039, w_021_188);
  nand2 I061_307(w_061_307, w_014_141, w_013_015);
  not1 I061_311(w_061_311, w_016_000);
  or2  I061_313(w_061_313, w_050_546, w_043_037);
  or2  I061_314(w_061_314, w_057_078, w_013_040);
  and2 I061_323(w_061_323, w_003_068, w_004_130);
  nand2 I061_326(w_061_326, w_004_372, w_028_321);
  nand2 I061_338(w_061_338, w_052_020, w_038_022);
  nand2 I061_343(w_061_343, w_016_008, w_049_341);
  not1 I061_356(w_061_356, w_018_028);
  and2 I061_357(w_061_357, w_033_631, w_013_583);
  nand2 I061_365(w_061_365, w_032_507, w_007_431);
  nand2 I061_374(w_061_374, w_044_384, w_016_003);
  nand2 I061_380(w_061_380, w_006_018, w_000_278);
  not1 I061_383(w_061_383, w_053_095);
  not1 I061_388(w_061_388, w_034_060);
  and2 I061_405(w_061_405, w_001_031, w_023_003);
  not1 I061_407(w_061_407, w_026_600);
  and2 I061_408(w_061_408, w_029_050, w_040_360);
  and2 I061_426(w_061_426, w_023_136, w_011_515);
  not1 I061_434(w_061_434, w_028_012);
  and2 I061_437(w_061_437, w_036_080, w_058_086);
  or2  I061_440(w_061_440, w_057_010, w_037_010);
  nand2 I061_443(w_061_443, w_006_013, w_000_780);
  not1 I061_452(w_061_452, w_024_478);
  not1 I061_464(w_061_464, w_010_057);
  or2  I061_465(w_061_465, w_050_148, w_021_033);
  and2 I061_467(w_061_467, w_024_164, w_025_242);
  and2 I061_472(w_061_472, w_007_199, w_026_274);
  or2  I061_473(w_061_473, w_027_157, w_050_024);
  or2  I061_477(w_061_477, w_002_560, w_016_007);
  nand2 I061_485(w_061_487, w_061_486, w_034_015);
  not1 I061_486(w_061_488, w_061_487);
  and2 I061_487(w_061_489, w_009_610, w_061_488);
  not1 I061_488(w_061_486, w_061_489);
  or2  I062_000(w_062_000, w_031_002, w_020_122);
  and2 I062_003(w_062_003, w_048_007, w_014_122);
  or2  I062_009(w_062_009, w_018_003, w_025_152);
  not1 I062_013(w_062_013, w_034_073);
  and2 I062_017(w_062_017, w_028_185, w_024_243);
  or2  I062_027(w_062_027, w_028_204, w_012_088);
  and2 I062_030(w_062_030, w_061_161, w_047_230);
  and2 I062_057(w_062_057, w_046_236, w_053_055);
  nand2 I062_058(w_062_058, w_031_182, w_044_666);
  or2  I062_060(w_062_060, w_030_119, w_060_003);
  and2 I062_081(w_062_081, w_037_031, w_046_323);
  nand2 I062_083(w_062_083, w_004_435, w_039_005);
  or2  I062_088(w_062_088, w_026_070, w_008_142);
  not1 I062_089(w_062_089, w_055_022);
  or2  I062_093(w_062_093, w_029_015, w_024_373);
  and2 I062_096(w_062_096, w_052_031, w_049_292);
  nand2 I062_099(w_062_099, w_019_001, w_040_425);
  nand2 I062_100(w_062_100, w_007_187, w_028_069);
  and2 I062_116(w_062_116, w_020_512, w_025_064);
  nand2 I062_125(w_062_125, w_050_071, w_058_162);
  nand2 I062_128(w_062_128, w_049_236, w_036_126);
  or2  I062_131(w_062_131, w_032_053, w_026_051);
  and2 I062_132(w_062_132, w_018_037, w_013_344);
  or2  I062_134(w_062_134, w_021_187, w_058_254);
  not1 I062_135(w_062_135, w_033_380);
  nand2 I062_138(w_062_138, w_052_028, w_053_053);
  not1 I062_140(w_062_140, w_011_315);
  or2  I062_144(w_062_144, w_045_023, w_036_274);
  and2 I062_149(w_062_149, w_020_489, w_008_331);
  or2  I062_151(w_062_151, w_030_261, w_012_071);
  nand2 I062_157(w_062_157, w_046_494, w_044_127);
  and2 I062_159(w_062_159, w_053_136, w_021_158);
  and2 I062_162(w_062_162, w_041_257, w_036_245);
  or2  I062_164(w_062_164, w_020_586, w_054_176);
  nand2 I062_168(w_062_168, w_010_769, w_031_009);
  not1 I062_173(w_062_173, w_055_018);
  or2  I062_177(w_062_177, w_003_030, w_042_310);
  or2  I062_178(w_062_178, w_037_207, w_056_119);
  not1 I062_185(w_062_185, w_043_025);
  not1 I062_194(w_062_194, w_052_040);
  and2 I062_206(w_062_206, w_057_230, w_045_109);
  or2  I062_208(w_062_208, w_046_452, w_031_119);
  not1 I062_211(w_062_211, w_025_063);
  and2 I062_220(w_062_220, w_050_164, w_046_013);
  not1 I062_224(w_062_224, w_004_031);
  not1 I062_229(w_062_229, w_056_505);
  not1 I062_239(w_062_239, w_059_596);
  and2 I062_241(w_062_241, w_000_185, w_055_243);
  not1 I062_245(w_062_245, w_034_037);
  not1 I062_249(w_062_249, w_001_031);
  nand2 I062_250(w_062_250, w_056_020, w_000_192);
  and2 I062_251(w_062_251, w_041_073, w_048_014);
  not1 I062_253(w_062_253, w_052_022);
  not1 I062_259(w_062_259, w_009_591);
  and2 I062_264(w_062_264, w_031_588, w_043_033);
  nand2 I062_268(w_062_268, w_021_017, w_049_070);
  or2  I062_273(w_062_273, w_055_337, w_028_284);
  nand2 I062_280(w_062_280, w_011_366, w_040_357);
  and2 I062_282(w_062_282, w_053_005, w_051_172);
  nand2 I062_305(w_062_305, w_014_002, w_029_105);
  not1 I062_307(w_062_307, w_007_017);
  not1 I062_308(w_062_308, w_033_029);
  and2 I062_311(w_062_311, w_022_145, w_057_279);
  and2 I062_313(w_062_313, w_055_142, w_008_576);
  nand2 I062_316(w_062_316, w_028_068, w_042_012);
  nand2 I062_329(w_062_329, w_021_083, w_021_082);
  nand2 I062_330(w_062_330, w_030_013, w_008_352);
  and2 I062_338(w_062_338, w_033_127, w_037_236);
  and2 I062_342(w_062_342, w_017_245, w_028_228);
  nand2 I062_349(w_062_349, w_004_344, w_000_329);
  or2  I062_352(w_062_352, w_048_019, w_040_515);
  not1 I062_355(w_062_355, w_005_110);
  nand2 I062_362(w_062_362, w_013_582, w_013_203);
  nand2 I062_370(w_062_370, w_033_157, w_055_090);
  not1 I062_371(w_062_371, w_013_121);
  and2 I062_377(w_062_377, w_006_220, w_050_138);
  or2  I062_378(w_062_378, w_057_053, w_022_183);
  or2  I062_380(w_062_380, w_043_011, w_021_210);
  not1 I062_384(w_062_384, w_019_002);
  nand2 I062_390(w_062_390, w_008_692, w_021_270);
  or2  I062_401(w_062_401, w_036_231, w_042_039);
  nand2 I062_406(w_062_406, w_030_008, w_019_011);
  and2 I062_430(w_062_430, w_037_233, w_048_010);
  and2 I062_435(w_062_435, w_002_012, w_014_116);
  and2 I062_440(w_062_440, w_059_313, w_017_103);
  and2 I062_455(w_062_455, w_050_222, w_047_280);
  or2  I062_458(w_062_458, w_052_014, w_002_421);
  and2 I062_465(w_062_465, w_016_001, w_036_266);
  not1 I062_473(w_062_473, w_049_268);
  or2  I062_483(w_062_483, w_026_023, w_014_282);
  and2 I062_484(w_062_484, w_006_103, w_020_460);
  not1 I062_503(w_062_503, w_056_082);
  not1 I062_508(w_062_508, w_023_025);
  or2  I062_511(w_062_511, w_052_005, w_010_270);
  and2 I062_512(w_062_512, w_001_002, w_018_007);
  or2  I062_513(w_062_513, w_011_224, w_028_228);
  nand2 I062_516(w_062_516, w_025_099, w_045_144);
  and2 I062_517(w_062_517, w_016_002, w_038_138);
  not1 I062_518(w_062_518, w_004_402);
  or2  I062_526(w_062_526, w_057_107, w_031_588);
  not1 I062_535(w_062_535, w_017_124);
  or2  I062_539(w_062_539, w_036_173, w_059_239);
  nand2 I062_540(w_062_540, w_054_145, w_049_005);
  and2 I062_544(w_062_544, w_013_232, w_005_124);
  not1 I062_546(w_062_546, w_020_172);
  or2  I062_549(w_062_549, w_020_398, w_057_019);
  nand2 I062_554(w_062_554, w_027_192, w_053_112);
  not1 I062_586(w_062_586, w_045_289);
  and2 I062_591(w_062_591, w_045_386, w_005_155);
  nand2 I062_593(w_062_593, w_041_244, w_003_071);
  and2 I062_598(w_062_598, w_019_008, w_023_060);
  and2 I062_606(w_062_606, w_044_628, w_056_661);
  and2 I062_607(w_062_607, w_019_016, w_037_003);
  or2  I062_612(w_062_612, w_010_148, w_031_016);
  and2 I062_628(w_062_628, w_058_655, w_018_006);
  not1 I062_633(w_062_633, w_008_661);
  or2  I062_643(w_062_643, w_013_030, w_012_226);
  nand2 I062_653(w_062_653, w_044_473, w_030_020);
  not1 I062_661(w_062_661, w_037_310);
  and2 I062_666(w_062_666, w_027_173, w_028_132);
  nand2 I062_670(w_062_670, w_014_081, w_049_036);
  and2 I062_672(w_062_672, w_045_345, w_059_315);
  not1 I062_673(w_062_673, w_050_532);
  nand2 I062_677(w_062_677, w_019_014, w_038_093);
  or2  I062_689(w_062_689, w_045_366, w_016_001);
  or2  I062_696(w_062_696, w_053_093, w_057_063);
  not1 I062_697(w_062_697, w_042_433);
  and2 I062_704(w_062_704, w_047_370, w_059_633);
  and2 I062_718(w_062_718, w_016_002, w_019_009);
  nand2 I062_731(w_062_731, w_024_024, w_002_074);
  not1 I062_732(w_062_732, w_053_087);
  not1 I062_734(w_062_734, w_003_059);
  not1 I062_739(w_062_739, w_008_653);
  and2 I062_745(w_062_745, w_047_248, w_022_188);
  and2 I062_761(w_062_761, w_034_032, w_050_267);
  and2 I062_768(w_062_768, w_023_000, w_017_264);
  or2  I062_772(w_062_772, w_050_032, w_033_629);
  not1 I062_776(w_062_776, w_001_006);
  nand2 I062_784(w_062_784, w_052_037, w_040_252);
  and2 I062_785(w_062_785, w_047_268, w_020_004);
  and2 I062_796(w_062_796, w_025_056, w_033_560);
  nand2 I063_002(w_063_002, w_048_014, w_003_031);
  nand2 I063_003(w_063_003, w_021_101, w_030_180);
  and2 I063_004(w_063_004, w_028_440, w_044_046);
  or2  I063_005(w_063_005, w_059_482, w_027_012);
  nand2 I063_006(w_063_006, w_041_489, w_019_003);
  not1 I063_008(w_063_008, w_044_487);
  and2 I063_009(w_063_009, w_047_229, w_057_243);
  and2 I063_010(w_063_010, w_022_365, w_044_033);
  or2  I063_014(w_063_014, w_010_211, w_054_088);
  not1 I063_018(w_063_018, w_001_001);
  or2  I063_019(w_063_019, w_030_223, w_055_156);
  nand2 I063_024(w_063_024, w_008_127, w_042_157);
  not1 I063_025(w_063_025, w_049_079);
  not1 I063_026(w_063_026, w_011_056);
  not1 I063_027(w_063_027, w_032_213);
  nand2 I063_029(w_063_029, w_049_207, w_042_325);
  and2 I063_034(w_063_034, w_044_046, w_061_253);
  nand2 I063_035(w_063_035, w_025_024, w_042_319);
  nand2 I063_036(w_063_036, w_024_030, w_019_012);
  not1 I063_045(w_063_045, w_012_027);
  and2 I063_047(w_063_047, w_044_022, w_032_285);
  and2 I063_050(w_063_050, w_029_001, w_058_467);
  or2  I063_052(w_063_052, w_062_132, w_044_026);
  and2 I063_058(w_063_058, w_052_005, w_014_142);
  and2 I063_059(w_063_059, w_056_314, w_059_554);
  and2 I063_062(w_063_062, w_042_318, w_019_011);
  or2  I063_063(w_063_063, w_046_037, w_040_568);
  or2  I063_064(w_063_064, w_048_004, w_029_021);
  not1 I063_066(w_063_066, w_054_141);
  and2 I063_072(w_063_072, w_043_033, w_020_409);
  not1 I063_073(w_063_073, w_053_139);
  and2 I063_076(w_063_076, w_047_383, w_039_656);
  nand2 I063_082(w_063_082, w_007_127, w_049_372);
  and2 I063_083(w_063_083, w_025_051, w_006_177);
  or2  I063_084(w_063_084, w_026_520, w_018_010);
  nand2 I063_085(w_063_085, w_023_108, w_019_016);
  and2 I063_086(w_063_086, w_005_017, w_041_463);
  or2  I063_088(w_063_088, w_047_220, w_006_107);
  or2  I063_089(w_063_089, w_029_036, w_049_232);
  and2 I063_090(w_063_090, w_045_268, w_039_240);
  nand2 I063_093(w_063_093, w_015_070, w_029_033);
  and2 I063_094(w_063_094, w_050_237, w_027_202);
  or2  I063_101(w_063_101, w_000_163, w_008_014);
  and2 I063_104(w_063_104, w_037_141, w_029_114);
  not1 I063_107(w_063_107, w_039_427);
  or2  I063_108(w_063_108, w_047_407, w_048_017);
  nand2 I063_109(w_063_109, w_047_080, w_013_063);
  not1 I063_110(w_063_110, w_014_046);
  nand2 I063_111(w_063_111, w_050_036, w_038_087);
  not1 I063_113(w_063_113, w_019_016);
  and2 I063_114(w_063_114, w_034_011, w_056_017);
  or2  I063_115(w_063_115, w_038_365, w_011_066);
  nand2 I063_120(w_063_120, w_014_233, w_030_199);
  or2  I063_121(w_063_121, w_023_073, w_016_002);
  nand2 I063_123(w_063_123, w_018_040, w_020_394);
  not1 I063_128(w_063_128, w_012_076);
  nand2 I063_133(w_063_133, w_052_037, w_042_222);
  nand2 I063_139(w_063_139, w_051_120, w_012_256);
  and2 I063_142(w_063_142, w_042_056, w_028_078);
  not1 I063_149(w_063_149, w_041_627);
  nand2 I063_153(w_063_153, w_050_211, w_020_272);
  or2  I063_155(w_063_155, w_042_113, w_041_117);
  nand2 I063_156(w_063_156, w_028_171, w_006_044);
  and2 I063_160(w_063_160, w_012_198, w_022_378);
  and2 I063_166(w_063_166, w_042_148, w_059_005);
  or2  I063_173(w_063_173, w_015_121, w_055_139);
  not1 I063_175(w_063_175, w_050_376);
  not1 I063_176(w_063_176, w_055_038);
  nand2 I063_177(w_063_177, w_053_082, w_040_164);
  and2 I063_178(w_063_178, w_018_026, w_026_275);
  not1 I063_179(w_063_179, w_032_504);
  or2  I063_180(w_063_180, w_036_020, w_057_083);
  not1 I063_181(w_063_181, w_011_592);
  nand2 I063_183(w_063_183, w_043_023, w_055_202);
  or2  I063_188(w_063_188, w_016_007, w_053_079);
  not1 I063_190(w_063_190, w_005_151);
  and2 I063_193(w_063_193, w_019_005, w_007_191);
  nand2 I063_194(w_063_194, w_012_026, w_043_003);
  or2  I063_197(w_063_197, w_020_146, w_034_002);
  or2  I063_198(w_063_198, w_030_177, w_014_111);
  and2 I063_208(w_063_208, w_046_267, w_044_598);
  nand2 I063_212(w_063_212, w_061_082, w_006_180);
  not1 I063_213(w_063_213, w_033_557);
  and2 I063_216(w_063_216, w_021_215, w_050_646);
  not1 I063_218(w_063_218, w_030_006);
  not1 I063_219(w_063_219, w_028_125);
  and2 I063_222(w_063_222, w_055_052, w_030_267);
  nand2 I063_223(w_063_223, w_044_632, w_057_239);
  not1 I063_224(w_063_224, w_054_425);
  and2 I063_225(w_063_225, w_006_039, w_054_026);
  not1 I063_226(w_063_226, w_010_420);
  or2  I063_227(w_063_227, w_050_646, w_041_531);
  or2  I063_228(w_063_228, w_061_052, w_028_505);
  or2  I063_229(w_063_229, w_020_455, w_015_096);
  not1 I063_233(w_063_233, w_062_598);
  or2  I063_238(w_063_238, w_005_072, w_037_253);
  not1 I063_244(w_063_244, w_017_103);
  or2  I063_245(w_063_245, w_053_093, w_001_021);
  nand2 I063_250(w_063_250, w_043_047, w_035_012);
  nand2 I063_251(w_063_251, w_021_032, w_055_187);
  nand2 I063_252(w_063_252, w_059_355, w_015_558);
  not1 I063_262(w_063_262, w_002_419);
  and2 I063_267(w_063_267, w_021_181, w_034_035);
  or2  I063_268(w_063_268, w_012_077, w_030_188);
  and2 I063_269(w_063_269, w_048_016, w_005_001);
  or2  I063_274(w_063_274, w_029_113, w_048_001);
  not1 I063_290(w_063_290, w_013_034);
  and2 I063_297(w_063_297, w_057_296, w_018_003);
  and2 I063_301(w_063_301, w_011_290, w_035_061);
  and2 I063_302(w_063_302, w_027_091, w_016_003);
  or2  I063_304(w_063_304, w_000_565, w_034_067);
  not1 I063_317(w_063_317, w_027_095);
  nand2 I063_319(w_063_319, w_050_584, w_005_153);
  or2  I063_326(w_063_326, w_026_114, w_027_199);
  and2 I063_341(w_063_341, w_033_017, w_027_020);
  nand2 I063_361(w_063_361, w_032_562, w_056_357);
  nand2 I063_366(w_063_366, w_026_699, w_050_543);
  nand2 I063_374(w_063_374, w_026_415, w_049_253);
  and2 I063_376(w_063_376, w_018_040, w_061_271);
  or2  I063_383(w_063_383, w_012_337, w_000_203);
  and2 I063_387(w_063_387, w_052_018, w_033_546);
  or2  I063_388(w_063_388, w_006_070, w_016_004);
  or2  I063_397(w_063_397, w_027_078, w_062_380);
  nand2 I063_400(w_063_400, w_032_099, w_040_123);
  not1 I063_402(w_063_402, w_021_025);
  and2 I063_410(w_063_410, w_022_181, w_015_208);
  not1 I063_415(w_063_415, w_057_246);
  not1 I063_417(w_063_417, w_008_320);
  not1 I063_418(w_063_418, w_016_002);
  nand2 I063_421(w_063_421, w_040_382, w_055_286);
  not1 I063_424(w_063_424, w_000_033);
  and2 I063_432(w_063_432, w_045_337, w_030_313);
  nand2 I063_438(w_063_438, w_020_407, w_002_076);
  or2  I063_445(w_063_445, w_046_121, w_058_366);
  and2 I063_450(w_063_450, w_055_085, w_035_015);
  or2  I063_456(w_063_456, w_040_298, w_019_006);
  nand2 I063_469(w_063_469, w_040_164, w_003_001);
  not1 I063_470(w_063_470, w_032_110);
  nand2 I063_483(w_063_483, w_015_166, w_018_040);
  or2  I063_503(w_063_503, w_054_170, w_042_092);
  not1 I063_504(w_063_504, w_018_037);
  nand2 I063_509(w_063_509, w_028_085, w_055_242);
  and2 I063_514(w_063_514, w_031_011, w_007_240);
  and2 I063_519(w_063_519, w_008_029, w_033_293);
  or2  I063_524(w_063_524, w_035_104, w_062_009);
  not1 I063_527(w_063_527, w_027_178);
  and2 I063_528(w_063_528, w_007_015, w_040_008);
  or2  I063_545(w_063_545, w_030_318, w_047_051);
  nand2 I063_547(w_063_547, w_039_680, w_012_181);
  and2 I064_004(w_064_004, w_025_154, w_063_470);
  or2  I064_005(w_064_005, w_016_001, w_000_541);
  not1 I064_009(w_064_009, w_062_305);
  not1 I064_010(w_064_010, w_011_364);
  not1 I064_012(w_064_012, w_026_082);
  nand2 I064_014(w_064_014, w_057_088, w_057_114);
  nand2 I064_018(w_064_018, w_063_528, w_052_013);
  and2 I064_020(w_064_020, w_023_149, w_055_215);
  nand2 I064_027(w_064_027, w_007_126, w_019_001);
  not1 I064_029(w_064_029, w_015_641);
  not1 I064_032(w_064_032, w_000_434);
  not1 I064_034(w_064_034, w_003_076);
  or2  I064_036(w_064_036, w_006_023, w_052_036);
  and2 I064_038(w_064_038, w_062_731, w_019_004);
  and2 I064_044(w_064_044, w_051_348, w_016_002);
  nand2 I064_049(w_064_049, w_017_616, w_003_030);
  not1 I064_052(w_064_052, w_055_015);
  and2 I064_055(w_064_055, w_045_198, w_056_434);
  nand2 I064_056(w_064_056, w_055_132, w_046_611);
  not1 I064_058(w_064_058, w_043_043);
  or2  I064_059(w_064_059, w_006_082, w_004_368);
  or2  I064_061(w_064_061, w_057_203, w_046_230);
  or2  I064_064(w_064_064, w_058_112, w_040_549);
  and2 I064_066(w_064_066, w_026_193, w_027_043);
  nand2 I064_069(w_064_069, w_042_113, w_058_164);
  not1 I064_070(w_064_070, w_047_279);
  not1 I064_072(w_064_072, w_037_314);
  or2  I064_074(w_064_074, w_014_175, w_017_434);
  and2 I064_077(w_064_077, w_009_072, w_063_402);
  nand2 I064_078(w_064_078, w_015_033, w_033_404);
  nand2 I064_080(w_064_080, w_002_347, w_034_055);
  or2  I064_081(w_064_081, w_037_147, w_041_104);
  and2 I064_082(w_064_082, w_009_533, w_046_580);
  and2 I064_086(w_064_086, w_040_027, w_045_284);
  nand2 I064_087(w_064_087, w_047_121, w_049_066);
  not1 I064_093(w_064_093, w_043_000);
  nand2 I064_094(w_064_094, w_032_287, w_058_304);
  or2  I064_097(w_064_097, w_023_052, w_015_051);
  nand2 I064_100(w_064_100, w_039_030, w_022_199);
  nand2 I064_103(w_064_103, w_031_315, w_003_025);
  or2  I064_106(w_064_106, w_037_302, w_005_125);
  nand2 I064_107(w_064_107, w_036_148, w_014_049);
  and2 I064_111(w_064_111, w_044_029, w_062_539);
  and2 I064_112(w_064_112, w_020_192, w_018_024);
  not1 I064_114(w_064_114, w_014_015);
  nand2 I064_115(w_064_115, w_050_305, w_052_014);
  not1 I064_118(w_064_118, w_043_031);
  and2 I064_121(w_064_121, w_024_207, w_003_044);
  not1 I064_125(w_064_125, w_044_312);
  not1 I064_127(w_064_127, w_009_293);
  and2 I064_130(w_064_130, w_063_153, w_034_041);
  not1 I064_133(w_064_133, w_041_041);
  and2 I064_134(w_064_134, w_057_007, w_030_287);
  and2 I064_135(w_064_135, w_039_040, w_048_011);
  or2  I064_136(w_064_136, w_059_567, w_026_663);
  and2 I064_140(w_064_140, w_030_250, w_052_027);
  not1 I064_142(w_064_142, w_057_095);
  not1 I064_143(w_064_143, w_024_116);
  not1 I064_150(w_064_150, w_057_220);
  not1 I064_153(w_064_153, w_010_616);
  not1 I064_154(w_064_154, w_010_095);
  nand2 I064_155(w_064_155, w_042_139, w_006_069);
  and2 I064_165(w_064_165, w_002_499, w_049_035);
  not1 I064_166(w_064_166, w_022_119);
  or2  I064_170(w_064_170, w_037_022, w_010_519);
  or2  I064_174(w_064_174, w_017_101, w_041_051);
  and2 I064_180(w_064_180, w_062_149, w_048_019);
  nand2 I064_182(w_064_182, w_052_045, w_027_103);
  nand2 I064_184(w_064_184, w_032_425, w_033_061);
  or2  I064_194(w_064_194, w_002_694, w_050_266);
  nand2 I064_197(w_064_197, w_048_012, w_011_016);
  not1 I064_202(w_064_202, w_057_229);
  and2 I064_205(w_064_205, w_009_623, w_054_283);
  and2 I064_207(w_064_207, w_040_505, w_022_272);
  and2 I064_214(w_064_214, w_033_629, w_025_163);
  nand2 I064_215(w_064_215, w_021_086, w_023_208);
  not1 I064_226(w_064_226, w_027_187);
  nand2 I064_228(w_064_228, w_015_135, w_031_434);
  or2  I064_229(w_064_229, w_053_098, w_021_043);
  nand2 I064_233(w_064_233, w_024_273, w_038_099);
  and2 I064_235(w_064_235, w_031_272, w_043_023);
  or2  I064_237(w_064_237, w_015_174, w_002_372);
  nand2 I064_241(w_064_241, w_050_488, w_024_109);
  or2  I064_253(w_064_253, w_051_348, w_007_096);
  not1 I064_255(w_064_255, w_015_055);
  and2 I064_256(w_064_256, w_019_009, w_025_035);
  and2 I064_265(w_064_265, w_047_158, w_028_117);
  nand2 I064_267(w_064_267, w_021_216, w_039_295);
  and2 I064_271(w_064_271, w_063_418, w_049_107);
  or2  I064_279(w_064_279, w_058_037, w_021_090);
  or2  I064_280(w_064_280, w_033_068, w_017_579);
  or2  I064_285(w_064_285, w_043_005, w_050_480);
  not1 I064_286(w_064_286, w_052_036);
  not1 I064_289(w_064_289, w_053_038);
  and2 I064_297(w_064_297, w_036_014, w_024_324);
  or2  I064_306(w_064_306, w_042_186, w_058_235);
  or2  I064_308(w_064_308, w_007_310, w_017_475);
  not1 I064_310(w_064_310, w_000_008);
  not1 I064_311(w_064_311, w_028_564);
  or2  I064_312(w_064_312, w_021_004, w_023_079);
  or2  I064_315(w_064_315, w_041_389, w_056_289);
  nand2 I064_324(w_064_324, w_010_289, w_012_327);
  not1 I064_327(w_064_327, w_010_181);
  or2  I064_328(w_064_328, w_041_476, w_025_116);
  not1 I064_329(w_064_329, w_061_003);
  nand2 I064_330(w_064_330, w_055_294, w_002_262);
  and2 I064_335(w_064_335, w_000_100, w_018_001);
  or2  I064_338(w_064_338, w_020_131, w_001_013);
  not1 I064_339(w_064_339, w_034_054);
  and2 I064_345(w_064_345, w_043_011, w_056_655);
  or2  I065_000(w_065_000, w_016_005, w_058_282);
  or2  I065_010(w_065_010, w_056_528, w_063_113);
  and2 I065_012(w_065_012, w_036_121, w_040_699);
  not1 I065_015(w_065_015, w_027_164);
  not1 I065_016(w_065_016, w_019_014);
  and2 I065_026(w_065_026, w_050_234, w_013_399);
  or2  I065_028(w_065_028, w_020_441, w_010_185);
  and2 I065_031(w_065_031, w_046_176, w_051_248);
  not1 I065_032(w_065_032, w_033_009);
  and2 I065_038(w_065_038, w_034_034, w_046_279);
  not1 I065_040(w_065_040, w_050_004);
  nand2 I065_043(w_065_043, w_060_003, w_043_001);
  or2  I065_046(w_065_046, w_035_021, w_050_520);
  nand2 I065_056(w_065_056, w_004_399, w_031_082);
  not1 I065_058(w_065_058, w_054_440);
  nand2 I065_059(w_065_059, w_035_076, w_047_224);
  and2 I065_060(w_065_060, w_059_328, w_054_228);
  or2  I065_063(w_065_063, w_042_252, w_026_045);
  and2 I065_066(w_065_066, w_020_240, w_042_165);
  and2 I065_069(w_065_069, w_058_453, w_056_071);
  not1 I065_074(w_065_074, w_054_084);
  nand2 I065_075(w_065_075, w_021_026, w_004_236);
  and2 I065_084(w_065_084, w_037_195, w_003_043);
  nand2 I065_086(w_065_086, w_034_008, w_023_033);
  nand2 I065_087(w_065_087, w_025_112, w_016_005);
  nand2 I065_095(w_065_095, w_048_009, w_054_176);
  and2 I065_097(w_065_097, w_008_291, w_064_327);
  not1 I065_098(w_065_098, w_009_402);
  and2 I065_107(w_065_107, w_052_039, w_042_414);
  or2  I065_117(w_065_117, w_005_180, w_030_155);
  or2  I065_126(w_065_126, w_015_188, w_020_114);
  not1 I065_132(w_065_132, w_012_019);
  or2  I065_136(w_065_136, w_036_073, w_003_052);
  or2  I065_144(w_065_144, w_047_047, w_021_105);
  not1 I065_152(w_065_152, w_049_281);
  and2 I065_165(w_065_165, w_000_047, w_058_503);
  not1 I065_172(w_065_172, w_045_182);
  nand2 I065_174(w_065_174, w_051_052, w_035_004);
  and2 I065_181(w_065_181, w_051_063, w_017_597);
  or2  I065_185(w_065_185, w_055_129, w_046_631);
  or2  I065_214(w_065_214, w_042_260, w_011_208);
  nand2 I065_218(w_065_218, w_053_014, w_016_007);
  nand2 I065_228(w_065_228, w_003_067, w_021_099);
  or2  I065_244(w_065_244, w_005_072, w_020_236);
  not1 I065_246(w_065_246, w_054_521);
  not1 I065_248(w_065_248, w_039_352);
  not1 I065_250(w_065_250, w_019_012);
  nand2 I065_253(w_065_253, w_051_138, w_032_098);
  and2 I065_256(w_065_256, w_064_064, w_008_407);
  or2  I065_259(w_065_259, w_052_012, w_009_512);
  not1 I065_263(w_065_263, w_005_197);
  or2  I065_270(w_065_270, w_010_770, w_058_132);
  nand2 I065_272(w_065_272, w_006_028, w_002_228);
  nand2 I065_275(w_065_275, w_031_315, w_037_218);
  or2  I065_280(w_065_280, w_002_468, w_029_061);
  not1 I065_285(w_065_285, w_051_090);
  or2  I065_295(w_065_295, w_018_034, w_028_014);
  not1 I065_296(w_065_296, w_029_054);
  and2 I065_304(w_065_304, w_019_008, w_052_045);
  nand2 I065_307(w_065_307, w_012_115, w_062_135);
  and2 I065_311(w_065_311, w_055_123, w_004_197);
  or2  I065_316(w_065_316, w_015_187, w_044_082);
  and2 I065_320(w_065_320, w_020_554, w_033_675);
  nand2 I065_327(w_065_327, w_042_437, w_049_256);
  not1 I065_333(w_065_333, w_019_011);
  or2  I065_338(w_065_338, w_063_290, w_021_044);
  not1 I065_342(w_065_342, w_039_182);
  or2  I065_343(w_065_343, w_059_089, w_056_058);
  and2 I065_344(w_065_344, w_011_268, w_031_009);
  and2 I065_348(w_065_348, w_020_072, w_053_116);
  not1 I065_359(w_065_359, w_032_169);
  and2 I065_361(w_065_361, w_059_196, w_041_062);
  not1 I065_363(w_065_363, w_014_132);
  not1 I065_372(w_065_372, w_001_014);
  or2  I065_381(w_065_381, w_057_262, w_042_057);
  nand2 I065_386(w_065_386, w_041_525, w_056_022);
  not1 I065_387(w_065_387, w_009_042);
  and2 I065_389(w_065_389, w_014_197, w_048_005);
  nand2 I065_393(w_065_393, w_015_570, w_053_021);
  or2  I065_407(w_065_407, w_049_079, w_043_045);
  or2  I065_411(w_065_411, w_002_121, w_008_398);
  or2  I065_425(w_065_425, w_039_380, w_031_206);
  or2  I065_426(w_065_426, w_055_108, w_034_030);
  or2  I065_449(w_065_449, w_021_123, w_021_007);
  and2 I065_453(w_065_453, w_019_019, w_021_223);
  not1 I065_474(w_065_474, w_052_027);
  nand2 I065_496(w_065_496, w_062_697, w_002_711);
  and2 I065_499(w_065_499, w_041_054, w_029_001);
  and2 I065_507(w_065_507, w_055_191, w_046_483);
  or2  I065_512(w_065_512, w_049_322, w_051_203);
  nand2 I065_515(w_065_515, w_038_018, w_022_366);
  not1 I065_517(w_065_517, w_028_080);
  or2  I065_522(w_065_522, w_052_035, w_035_031);
  nand2 I065_537(w_065_537, w_012_058, w_006_061);
  or2  I065_542(w_065_542, w_010_358, w_024_244);
  and2 I065_543(w_065_543, w_037_055, w_041_457);
  and2 I065_547(w_065_547, w_061_029, w_036_302);
  nand2 I065_555(w_065_555, w_016_008, w_026_261);
  and2 I065_557(w_065_557, w_023_157, w_055_282);
  or2  I065_558(w_065_558, w_042_220, w_020_483);
  nand2 I065_563(w_065_563, w_016_000, w_011_081);
  nand2 I065_565(w_065_565, w_032_011, w_016_007);
  nand2 I065_569(w_065_569, w_019_015, w_063_326);
  and2 I065_572(w_065_572, w_033_272, w_051_141);
  nand2 I065_576(w_065_576, w_063_121, w_007_217);
  not1 I065_582(w_065_582, w_058_316);
  or2  I065_590(w_065_590, w_036_114, w_061_126);
  and2 I065_593(w_065_593, w_051_165, w_026_121);
  not1 I065_603(w_065_603, w_033_779);
  not1 I065_606(w_065_606, w_014_022);
  and2 I065_609(w_065_609, w_051_115, w_038_070);
  not1 I065_641(w_065_641, w_018_013);
  not1 I065_646(w_065_646, w_000_415);
  nand2 I065_654(w_065_654, w_017_576, w_020_210);
  or2  I065_658(w_065_658, w_038_591, w_058_454);
  or2  I065_666(w_065_666, w_004_244, w_056_702);
  not1 I065_668(w_065_668, w_049_164);
  nand2 I065_673(w_065_673, w_011_606, w_058_086);
  not1 I065_687(w_065_687, w_056_457);
  and2 I066_004(w_066_004, w_034_010, w_056_545);
  nand2 I066_007(w_066_007, w_014_181, w_020_379);
  and2 I066_011(w_066_011, w_028_275, w_063_082);
  and2 I066_013(w_066_013, w_043_020, w_010_369);
  not1 I066_017(w_066_017, w_011_605);
  nand2 I066_023(w_066_023, w_059_249, w_054_347);
  nand2 I066_025(w_066_025, w_051_260, w_057_200);
  nand2 I066_029(w_066_029, w_045_039, w_004_040);
  or2  I066_035(w_066_035, w_062_128, w_042_172);
  and2 I066_040(w_066_040, w_009_031, w_063_008);
  and2 I066_045(w_066_045, w_023_083, w_045_259);
  not1 I066_052(w_066_052, w_004_004);
  and2 I066_058(w_066_058, w_064_154, w_019_006);
  not1 I066_061(w_066_061, w_040_083);
  nand2 I066_063(w_066_063, w_005_198, w_050_247);
  not1 I066_064(w_066_064, w_053_061);
  or2  I066_072(w_066_072, w_015_208, w_001_029);
  nand2 I066_080(w_066_080, w_034_039, w_008_758);
  nand2 I066_084(w_066_084, w_056_645, w_048_018);
  nand2 I066_089(w_066_089, w_018_028, w_017_017);
  or2  I066_093(w_066_093, w_046_164, w_011_179);
  not1 I066_095(w_066_095, w_056_044);
  not1 I066_099(w_066_099, w_050_533);
  not1 I066_101(w_066_101, w_016_005);
  not1 I066_103(w_066_103, w_026_606);
  and2 I066_104(w_066_104, w_015_087, w_033_630);
  and2 I066_110(w_066_110, w_042_402, w_055_302);
  nand2 I066_111(w_066_111, w_022_068, w_043_028);
  or2  I066_112(w_066_112, w_055_337, w_025_019);
  not1 I066_115(w_066_115, w_061_033);
  not1 I066_118(w_066_118, w_045_334);
  nand2 I066_119(w_066_119, w_034_071, w_020_050);
  and2 I066_123(w_066_123, w_051_354, w_025_165);
  and2 I066_125(w_066_125, w_014_215, w_049_140);
  not1 I066_126(w_066_126, w_004_104);
  and2 I066_134(w_066_134, w_051_358, w_018_032);
  or2  I066_135(w_066_135, w_032_057, w_031_058);
  and2 I066_141(w_066_141, w_054_417, w_023_093);
  nand2 I066_147(w_066_147, w_039_079, w_015_100);
  nand2 I066_154(w_066_154, w_051_095, w_032_074);
  nand2 I066_170(w_066_170, w_021_270, w_045_304);
  not1 I066_181(w_066_181, w_010_486);
  and2 I066_182(w_066_182, w_042_104, w_024_099);
  or2  I066_185(w_066_185, w_006_099, w_041_116);
  nand2 I066_191(w_066_191, w_004_255, w_055_089);
  nand2 I066_202(w_066_202, w_057_002, w_028_206);
  not1 I066_216(w_066_216, w_048_011);
  or2  I066_224(w_066_224, w_023_011, w_062_670);
  and2 I066_234(w_066_234, w_005_204, w_065_272);
  nand2 I066_240(w_066_240, w_022_220, w_043_000);
  and2 I066_243(w_066_243, w_059_337, w_065_059);
  nand2 I066_246(w_066_246, w_043_022, w_060_131);
  not1 I066_273(w_066_273, w_009_481);
  or2  I066_276(w_066_276, w_043_021, w_015_374);
  or2  I066_281(w_066_281, w_038_256, w_059_236);
  or2  I066_290(w_066_290, w_063_076, w_047_040);
  not1 I066_293(w_066_293, w_050_500);
  not1 I066_315(w_066_315, w_029_085);
  and2 I066_319(w_066_319, w_053_156, w_043_012);
  nand2 I066_327(w_066_327, w_062_473, w_053_099);
  or2  I066_335(w_066_335, w_046_660, w_025_040);
  and2 I066_341(w_066_341, w_002_251, w_048_003);
  not1 I066_343(w_066_343, w_027_050);
  or2  I066_348(w_066_348, w_057_101, w_055_287);
  and2 I066_349(w_066_349, w_053_135, w_058_073);
  not1 I066_356(w_066_356, w_008_334);
  nand2 I066_370(w_066_370, w_061_472, w_046_575);
  not1 I066_372(w_066_372, w_004_295);
  not1 I066_376(w_066_376, w_038_397);
  and2 I066_378(w_066_378, w_002_610, w_007_102);
  and2 I066_385(w_066_385, w_031_202, w_009_417);
  and2 I066_402(w_066_402, w_064_330, w_022_039);
  and2 I066_403(w_066_403, w_064_106, w_030_210);
  nand2 I066_404(w_066_404, w_044_366, w_057_296);
  and2 I066_405(w_066_405, w_061_047, w_054_146);
  and2 I066_406(w_066_406, w_043_037, w_030_270);
  and2 I066_416(w_066_416, w_046_390, w_056_280);
  or2  I066_421(w_066_421, w_010_350, w_037_050);
  and2 I066_433(w_066_433, w_043_010, w_031_116);
  or2  I066_454(w_066_454, w_021_119, w_061_061);
  and2 I066_463(w_066_463, w_024_088, w_038_025);
  not1 I066_473(w_066_473, w_014_135);
  nand2 I066_476(w_066_476, w_007_166, w_012_002);
  and2 I066_482(w_066_482, w_063_108, w_040_693);
  not1 I066_489(w_066_489, w_035_056);
  or2  I066_493(w_066_493, w_047_273, w_009_152);
  not1 I066_503(w_066_503, w_062_027);
  nand2 I066_512(w_066_512, w_024_034, w_009_199);
  and2 I066_516(w_066_516, w_042_321, w_062_458);
  and2 I066_518(w_066_518, w_020_425, w_028_436);
  and2 I066_531(w_066_531, w_028_162, w_014_261);
  or2  I066_542(w_066_542, w_009_606, w_005_006);
  nand2 I066_544(w_066_544, w_023_142, w_022_384);
  or2  I066_555(w_066_555, w_063_179, w_057_243);
  and2 I066_556(w_066_556, w_059_002, w_024_064);
  nand2 I066_558(w_066_558, w_034_034, w_024_194);
  or2  I066_559(w_066_559, w_055_064, w_052_034);
  and2 I066_572(w_066_572, w_015_385, w_026_538);
  or2  I066_578(w_066_578, w_065_363, w_019_004);
  or2  I066_584(w_066_584, w_031_387, w_053_105);
  and2 I066_586(w_066_586, w_012_317, w_018_024);
  or2  I066_594(w_066_594, w_047_033, w_060_160);
  not1 I066_595(w_066_595, w_049_047);
  and2 I066_625(w_066_625, w_054_055, w_018_019);
  and2 I066_627(w_066_627, w_041_048, w_060_310);
  or2  I067_003(w_067_003, w_033_494, w_025_171);
  nand2 I067_005(w_067_005, w_039_054, w_019_017);
  and2 I067_007(w_067_007, w_000_593, w_040_017);
  nand2 I067_010(w_067_010, w_031_168, w_010_560);
  not1 I067_013(w_067_013, w_025_133);
  nand2 I067_020(w_067_020, w_052_036, w_013_214);
  and2 I067_021(w_067_021, w_020_072, w_000_008);
  not1 I067_024(w_067_024, w_055_114);
  nand2 I067_027(w_067_027, w_011_125, w_032_444);
  not1 I067_037(w_067_037, w_024_569);
  not1 I067_039(w_067_039, w_024_155);
  or2  I067_046(w_067_046, w_042_076, w_033_341);
  not1 I067_049(w_067_049, w_008_403);
  or2  I067_052(w_067_052, w_045_052, w_049_016);
  or2  I067_053(w_067_053, w_041_549, w_021_263);
  not1 I067_060(w_067_060, w_004_508);
  nand2 I067_062(w_067_062, w_002_526, w_027_072);
  or2  I067_069(w_067_069, w_005_005, w_033_380);
  nand2 I067_076(w_067_076, w_063_094, w_000_575);
  nand2 I067_083(w_067_083, w_026_597, w_042_323);
  not1 I067_094(w_067_094, w_015_552);
  or2  I067_099(w_067_099, w_065_069, w_016_003);
  or2  I067_101(w_067_101, w_054_240, w_025_000);
  and2 I067_104(w_067_104, w_023_043, w_040_012);
  or2  I067_111(w_067_111, w_047_232, w_011_015);
  or2  I067_113(w_067_113, w_044_261, w_032_042);
  or2  I067_119(w_067_119, w_058_673, w_040_639);
  nand2 I067_122(w_067_122, w_009_629, w_032_359);
  or2  I067_125(w_067_125, w_016_003, w_065_381);
  nand2 I067_126(w_067_126, w_056_255, w_013_053);
  not1 I067_133(w_067_133, w_019_016);
  nand2 I067_134(w_067_134, w_057_085, w_004_151);
  and2 I067_137(w_067_137, w_007_107, w_027_035);
  not1 I067_140(w_067_140, w_060_112);
  or2  I067_141(w_067_141, w_064_081, w_013_189);
  not1 I067_146(w_067_146, w_010_192);
  nand2 I067_150(w_067_150, w_027_041, w_028_437);
  or2  I067_154(w_067_154, w_003_019, w_009_083);
  not1 I067_156(w_067_156, w_016_000);
  nand2 I067_162(w_067_162, w_058_193, w_031_495);
  nand2 I067_163(w_067_163, w_065_668, w_002_505);
  nand2 I067_165(w_067_165, w_018_007, w_021_179);
  not1 I067_166(w_067_166, w_036_093);
  and2 I067_169(w_067_169, w_001_003, w_032_043);
  and2 I067_171(w_067_171, w_056_493, w_026_274);
  nand2 I067_175(w_067_175, w_057_262, w_065_244);
  or2  I067_196(w_067_196, w_036_101, w_053_067);
  and2 I067_199(w_067_199, w_019_009, w_039_537);
  not1 I067_201(w_067_201, w_064_127);
  nand2 I067_204(w_067_204, w_055_049, w_017_095);
  nand2 I067_206(w_067_206, w_017_080, w_027_156);
  not1 I067_211(w_067_211, w_039_005);
  not1 I067_213(w_067_213, w_010_085);
  and2 I067_224(w_067_224, w_060_058, w_003_011);
  nand2 I067_232(w_067_232, w_020_530, w_051_019);
  and2 I067_239(w_067_239, w_055_074, w_057_175);
  and2 I067_250(w_067_250, w_012_127, w_005_126);
  or2  I067_253(w_067_253, w_021_051, w_024_028);
  nand2 I067_254(w_067_254, w_032_033, w_041_100);
  nand2 I067_255(w_067_255, w_048_013, w_004_115);
  nand2 I067_263(w_067_263, w_055_014, w_053_106);
  and2 I067_266(w_067_266, w_028_274, w_052_046);
  and2 I067_270(w_067_270, w_028_299, w_024_299);
  and2 I067_273(w_067_273, w_011_215, w_003_036);
  or2  I067_275(w_067_275, w_005_196, w_057_112);
  nand2 I067_276(w_067_276, w_032_360, w_050_135);
  and2 I067_280(w_067_280, w_055_058, w_029_072);
  or2  I067_290(w_067_290, w_039_089, w_008_583);
  or2  I067_292(w_067_292, w_034_050, w_025_222);
  nand2 I067_297(w_067_297, w_030_102, w_030_006);
  and2 I067_302(w_067_302, w_001_002, w_055_116);
  or2  I067_305(w_067_305, w_025_305, w_000_266);
  or2  I067_316(w_067_316, w_026_146, w_011_083);
  or2  I067_318(w_067_318, w_065_342, w_039_401);
  and2 I067_326(w_067_326, w_043_044, w_053_155);
  nand2 I067_328(w_067_328, w_032_178, w_052_038);
  and2 I067_329(w_067_329, w_024_272, w_049_182);
  or2  I067_333(w_067_333, w_027_067, w_037_131);
  or2  I067_334(w_067_334, w_042_278, w_029_074);
  or2  I067_336(w_067_336, w_052_019, w_035_115);
  nand2 I067_342(w_067_342, w_051_075, w_010_395);
  and2 I067_343(w_067_343, w_045_319, w_013_013);
  nand2 I067_344(w_067_344, w_035_127, w_063_018);
  not1 I067_346(w_067_346, w_055_122);
  and2 I067_347(w_067_347, w_061_058, w_037_083);
  or2  I067_352(w_067_352, w_056_663, w_051_230);
  or2  I067_353(w_067_353, w_056_250, w_054_150);
  nand2 I067_356(w_067_356, w_045_336, w_045_170);
  nand2 I067_358(w_067_358, w_030_117, w_004_212);
  or2  I067_360(w_067_360, w_028_409, w_047_152);
  not1 I067_362(w_067_362, w_061_125);
  or2  I067_363(w_067_363, w_056_070, w_036_191);
  and2 I067_371(w_067_371, w_063_252, w_016_007);
  or2  I067_373(w_067_373, w_023_176, w_038_358);
  not1 I067_374(w_067_374, w_000_406);
  and2 I067_381(w_067_381, w_062_096, w_062_338);
  or2  I067_382(w_067_382, w_059_174, w_066_017);
  nand2 I067_383(w_067_383, w_006_227, w_061_106);
  not1 I067_390(w_067_390, w_057_285);
  not1 I067_395(w_067_395, w_051_348);
  and2 I068_000(w_068_000, w_067_346, w_034_070);
  and2 I068_001(w_068_001, w_020_426, w_009_115);
  and2 I068_008(w_068_008, w_041_243, w_022_300);
  nand2 I068_009(w_068_009, w_014_192, w_032_364);
  nand2 I068_011(w_068_011, w_046_024, w_057_210);
  and2 I068_012(w_068_012, w_006_100, w_015_252);
  not1 I068_024(w_068_024, w_006_027);
  not1 I068_030(w_068_030, w_038_503);
  or2  I068_041(w_068_041, w_020_118, w_017_048);
  nand2 I068_042(w_068_042, w_050_064, w_023_093);
  nand2 I068_052(w_068_052, w_062_677, w_007_394);
  nand2 I068_056(w_068_056, w_060_266, w_059_616);
  and2 I068_060(w_068_060, w_008_040, w_013_541);
  and2 I068_062(w_068_062, w_002_022, w_016_004);
  and2 I068_069(w_068_069, w_033_622, w_052_031);
  not1 I068_070(w_068_070, w_067_266);
  nand2 I068_074(w_068_074, w_002_024, w_029_042);
  nand2 I068_075(w_068_075, w_041_412, w_022_330);
  and2 I068_076(w_068_076, w_063_002, w_021_007);
  nand2 I068_079(w_068_079, w_041_496, w_033_355);
  or2  I068_080(w_068_080, w_049_313, w_045_326);
  or2  I068_081(w_068_081, w_045_379, w_053_093);
  and2 I068_082(w_068_082, w_022_304, w_002_015);
  and2 I068_083(w_068_083, w_059_683, w_065_425);
  not1 I068_084(w_068_084, w_036_125);
  not1 I068_086(w_068_086, w_045_228);
  nand2 I068_092(w_068_092, w_040_520, w_029_105);
  nand2 I068_094(w_068_094, w_035_077, w_063_009);
  nand2 I068_095(w_068_095, w_035_108, w_030_374);
  nand2 I068_098(w_068_098, w_042_343, w_038_322);
  or2  I068_101(w_068_101, w_059_637, w_009_044);
  and2 I068_102(w_068_102, w_044_013, w_011_542);
  or2  I068_106(w_068_106, w_064_228, w_067_003);
  and2 I068_113(w_068_113, w_024_283, w_023_096);
  or2  I068_114(w_068_114, w_027_122, w_000_293);
  and2 I068_124(w_068_124, w_003_083, w_056_509);
  not1 I068_125(w_068_125, w_022_003);
  and2 I068_131(w_068_131, w_033_604, w_000_258);
  or2  I068_133(w_068_133, w_035_127, w_008_418);
  nand2 I068_136(w_068_136, w_052_008, w_054_346);
  nand2 I068_138(w_068_138, w_045_180, w_005_041);
  not1 I068_139(w_068_139, w_055_309);
  not1 I068_153(w_068_153, w_016_002);
  nand2 I068_167(w_068_167, w_044_093, w_010_126);
  or2  I068_170(w_068_170, w_006_002, w_049_045);
  and2 I068_174(w_068_174, w_026_060, w_001_003);
  and2 I068_176(w_068_176, w_061_142, w_017_252);
  and2 I068_181(w_068_181, w_013_074, w_059_724);
  not1 I068_182(w_068_182, w_039_170);
  and2 I068_183(w_068_183, w_064_082, w_064_237);
  or2  I068_192(w_068_192, w_001_013, w_001_025);
  and2 I068_194(w_068_194, w_039_318, w_008_439);
  or2  I068_200(w_068_200, w_050_415, w_022_051);
  and2 I068_204(w_068_204, w_013_543, w_015_045);
  not1 I068_206(w_068_206, w_017_102);
  and2 I068_209(w_068_209, w_043_015, w_049_018);
  not1 I068_210(w_068_210, w_027_183);
  and2 I068_213(w_068_213, w_031_012, w_033_590);
  nand2 I068_221(w_068_221, w_052_027, w_051_233);
  nand2 I068_224(w_068_224, w_061_277, w_033_449);
  or2  I068_225(w_068_225, w_044_573, w_039_203);
  or2  I068_226(w_068_226, w_058_568, w_034_069);
  or2  I068_231(w_068_231, w_067_253, w_002_073);
  not1 I068_237(w_068_237, w_041_409);
  and2 I068_242(w_068_242, w_065_012, w_032_546);
  and2 I068_246(w_068_246, w_051_061, w_012_087);
  nand2 I068_249(w_068_249, w_012_152, w_021_222);
  and2 I068_250(w_068_250, w_058_570, w_059_209);
  or2  I068_260(w_068_260, w_030_341, w_028_170);
  or2  I068_265(w_068_265, w_051_367, w_035_019);
  and2 I068_267(w_068_267, w_046_137, w_008_093);
  nand2 I068_268(w_068_268, w_008_020, w_038_115);
  or2  I068_275(w_068_275, w_014_173, w_058_134);
  and2 I068_276(w_068_276, w_021_145, w_028_045);
  nand2 I068_280(w_068_280, w_006_035, w_030_012);
  and2 I068_283(w_068_283, w_025_049, w_000_314);
  not1 I068_295(w_068_295, w_026_483);
  or2  I068_298(w_068_298, w_004_126, w_049_309);
  and2 I068_301(w_068_301, w_027_153, w_039_030);
  or2  I068_304(w_068_304, w_030_248, w_014_234);
  and2 I068_306(w_068_306, w_051_069, w_058_136);
  and2 I068_307(w_068_307, w_030_379, w_016_003);
  or2  I068_308(w_068_308, w_046_106, w_034_013);
  or2  I068_309(w_068_309, w_062_672, w_016_005);
  and2 I068_321(w_068_321, w_038_164, w_027_019);
  and2 I068_322(w_068_322, w_019_010, w_053_065);
  and2 I068_323(w_068_323, w_000_590, w_050_031);
  not1 I068_328(w_068_328, w_003_053);
  and2 I068_334(w_068_334, w_007_128, w_051_370);
  or2  I068_337(w_068_337, w_067_119, w_023_201);
  or2  I068_340(w_068_340, w_024_026, w_061_383);
  and2 I068_342(w_068_342, w_016_008, w_021_021);
  nand2 I068_344(w_068_344, w_046_196, w_064_107);
  and2 I068_346(w_068_346, w_056_507, w_035_030);
  and2 I068_348(w_068_348, w_056_303, w_001_033);
  nand2 I068_349(w_068_349, w_063_317, w_063_063);
  or2  I068_352(w_068_352, w_014_004, w_065_087);
  or2  I068_357(w_068_357, w_025_123, w_052_027);
  nand2 I068_360(w_068_360, w_012_007, w_010_275);
  or2  I068_361(w_068_361, w_014_002, w_039_064);
  not1 I069_001(w_069_001, w_023_012);
  nand2 I069_003(w_069_003, w_024_144, w_047_325);
  nand2 I069_005(w_069_005, w_009_545, w_027_202);
  or2  I069_009(w_069_009, w_017_121, w_053_073);
  and2 I069_014(w_069_014, w_063_064, w_066_404);
  and2 I069_016(w_069_016, w_038_512, w_054_102);
  nand2 I069_022(w_069_022, w_003_003, w_032_120);
  and2 I069_023(w_069_023, w_022_236, w_068_125);
  not1 I069_025(w_069_025, w_067_027);
  or2  I069_028(w_069_028, w_054_588, w_012_338);
  nand2 I069_029(w_069_029, w_045_049, w_012_287);
  and2 I069_033(w_069_033, w_058_404, w_057_145);
  nand2 I069_034(w_069_034, w_024_000, w_002_052);
  not1 I069_038(w_069_038, w_018_016);
  not1 I069_039(w_069_039, w_022_013);
  nand2 I069_042(w_069_042, w_019_017, w_037_066);
  not1 I069_048(w_069_048, w_020_561);
  nand2 I069_049(w_069_049, w_028_523, w_021_137);
  nand2 I069_053(w_069_053, w_061_146, w_066_454);
  or2  I069_055(w_069_055, w_041_275, w_009_140);
  nand2 I069_060(w_069_060, w_023_011, w_002_605);
  nand2 I069_063(w_069_063, w_014_074, w_011_232);
  not1 I069_064(w_069_064, w_009_123);
  and2 I069_065(w_069_065, w_017_013, w_038_467);
  nand2 I069_067(w_069_067, w_000_725, w_020_474);
  or2  I069_068(w_069_068, w_050_317, w_013_053);
  and2 I069_071(w_069_071, w_064_094, w_034_008);
  nand2 I069_075(w_069_075, w_028_135, w_014_153);
  not1 I069_076(w_069_076, w_066_555);
  or2  I069_077(w_069_077, w_063_229, w_031_162);
  or2  I069_078(w_069_078, w_067_206, w_020_436);
  nand2 I069_080(w_069_080, w_009_627, w_006_120);
  not1 I069_081(w_069_081, w_005_053);
  nand2 I069_087(w_069_087, w_033_437, w_060_114);
  nand2 I069_088(w_069_088, w_036_408, w_041_113);
  nand2 I069_089(w_069_089, w_042_026, w_015_546);
  nand2 I069_091(w_069_091, w_004_484, w_046_699);
  nand2 I069_093(w_069_093, w_001_018, w_022_283);
  not1 I069_096(w_069_096, w_046_100);
  not1 I069_097(w_069_097, w_058_534);
  and2 I069_104(w_069_104, w_026_541, w_062_732);
  and2 I069_105(w_069_105, w_020_543, w_005_159);
  and2 I069_107(w_069_107, w_035_098, w_013_297);
  or2  I069_110(w_069_110, w_021_141, w_046_637);
  and2 I069_117(w_069_117, w_008_407, w_063_093);
  or2  I069_120(w_069_120, w_066_403, w_052_005);
  or2  I069_125(w_069_125, w_057_147, w_028_228);
  and2 I069_128(w_069_128, w_067_020, w_004_236);
  or2  I069_140(w_069_140, w_057_124, w_006_128);
  nand2 I069_141(w_069_141, w_010_511, w_065_393);
  and2 I069_143(w_069_143, w_066_378, w_064_205);
  and2 I069_144(w_069_144, w_034_038, w_024_482);
  or2  I069_145(w_069_145, w_058_095, w_060_081);
  and2 I069_146(w_069_146, w_062_338, w_038_260);
  not1 I069_153(w_069_153, w_009_046);
  not1 I069_157(w_069_157, w_037_232);
  nand2 I069_158(w_069_158, w_058_005, w_048_006);
  not1 I069_159(w_069_159, w_020_264);
  and2 I069_165(w_069_165, w_016_008, w_055_220);
  and2 I069_167(w_069_167, w_047_458, w_055_064);
  and2 I069_168(w_069_168, w_056_736, w_043_001);
  nand2 I069_171(w_069_171, w_051_380, w_041_541);
  or2  I069_173(w_069_173, w_014_119, w_005_237);
  or2  I069_174(w_069_174, w_052_012, w_052_025);
  not1 I069_176(w_069_176, w_021_068);
  not1 I069_177(w_069_177, w_064_235);
  and2 I069_181(w_069_181, w_025_036, w_065_361);
  and2 I069_182(w_069_182, w_062_540, w_032_247);
  nand2 I069_185(w_069_185, w_007_193, w_042_081);
  and2 I069_188(w_069_188, w_052_035, w_050_141);
  nand2 I069_191(w_069_191, w_032_207, w_054_104);
  nand2 I069_192(w_069_192, w_061_122, w_035_010);
  nand2 I069_194(w_069_194, w_062_718, w_050_138);
  or2  I069_197(w_069_197, w_062_144, w_005_309);
  not1 I069_199(w_069_199, w_028_006);
  nand2 I069_202(w_069_202, w_002_202, w_062_371);
  and2 I069_207(w_069_207, w_068_213, w_024_482);
  nand2 I069_209(w_069_209, w_011_231, w_047_031);
  or2  I069_213(w_069_213, w_007_473, w_023_151);
  and2 I069_218(w_069_218, w_027_062, w_062_633);
  and2 I069_223(w_069_223, w_000_375, w_046_377);
  or2  I069_225(w_069_225, w_011_099, w_067_134);
  nand2 I069_226(w_069_226, w_028_129, w_059_135);
  or2  I069_227(w_069_227, w_047_188, w_068_138);
  and2 I069_228(w_069_228, w_058_379, w_047_248);
  or2  I069_230(w_069_230, w_039_550, w_011_624);
  and2 I069_232(w_069_232, w_005_277, w_063_036);
  and2 I069_236(w_069_236, w_057_068, w_035_024);
  and2 I069_237(w_069_237, w_057_105, w_017_366);
  nand2 I069_241(w_069_241, w_034_062, w_055_084);
  not1 I069_242(w_069_242, w_039_377);
  or2  I069_245(w_069_245, w_030_252, w_002_159);
  nand2 I069_254(w_069_254, w_038_123, w_046_390);
  and2 I069_259(w_069_259, w_029_092, w_021_005);
  or2  I069_260(w_069_260, w_032_269, w_043_047);
  not1 I069_265(w_069_265, w_030_307);
  nand2 I070_000(w_070_000, w_027_000, w_023_175);
  or2  I070_004(w_070_004, w_066_004, w_060_333);
  not1 I070_006(w_070_006, w_015_272);
  nand2 I070_007(w_070_007, w_068_124, w_046_240);
  or2  I070_008(w_070_008, w_029_018, w_050_242);
  or2  I070_009(w_070_009, w_001_000, w_065_304);
  and2 I070_010(w_070_010, w_032_575, w_035_022);
  or2  I070_014(w_070_014, w_021_273, w_027_111);
  or2  I070_018(w_070_018, w_067_166, w_041_661);
  not1 I070_019(w_070_019, w_069_218);
  or2  I070_021(w_070_021, w_018_011, w_012_267);
  not1 I070_027(w_070_027, w_032_030);
  nand2 I070_028(w_070_028, w_051_268, w_023_031);
  not1 I070_031(w_070_031, w_068_008);
  and2 I070_033(w_070_033, w_016_004, w_034_031);
  or2  I070_035(w_070_035, w_060_278, w_036_239);
  nand2 I070_041(w_070_041, w_014_022, w_042_110);
  or2  I070_044(w_070_044, w_006_012, w_017_426);
  or2  I070_050(w_070_050, w_046_443, w_038_505);
  and2 I070_056(w_070_056, w_005_229, w_001_020);
  or2  I070_060(w_070_060, w_059_578, w_066_454);
  or2  I070_069(w_070_069, w_028_060, w_040_234);
  and2 I070_071(w_070_071, w_001_002, w_021_116);
  and2 I070_080(w_070_080, w_056_119, w_039_536);
  or2  I070_083(w_070_083, w_042_109, w_055_040);
  and2 I070_084(w_070_084, w_047_054, w_059_600);
  nand2 I070_089(w_070_089, w_000_426, w_051_318);
  or2  I070_096(w_070_096, w_018_020, w_055_041);
  nand2 I070_100(w_070_100, w_034_000, w_017_116);
  nand2 I070_104(w_070_104, w_061_242, w_056_009);
  or2  I070_108(w_070_108, w_011_003, w_009_100);
  nand2 I070_109(w_070_109, w_041_340, w_004_199);
  and2 I070_112(w_070_112, w_066_542, w_067_204);
  or2  I070_117(w_070_117, w_028_488, w_006_001);
  and2 I070_121(w_070_121, w_029_087, w_023_132);
  or2  I070_123(w_070_123, w_055_029, w_032_575);
  and2 I070_142(w_070_142, w_041_079, w_007_170);
  not1 I070_143(w_070_143, w_028_130);
  not1 I070_148(w_070_148, w_013_422);
  nand2 I070_155(w_070_155, w_008_587, w_056_094);
  not1 I070_158(w_070_158, w_003_019);
  nand2 I070_161(w_070_161, w_006_142, w_028_567);
  or2  I070_170(w_070_170, w_039_329, w_050_514);
  or2  I070_173(w_070_173, w_023_078, w_001_032);
  nand2 I070_174(w_070_174, w_017_280, w_064_004);
  or2  I070_175(w_070_175, w_028_521, w_030_263);
  or2  I070_179(w_070_179, w_025_102, w_051_113);
  or2  I070_185(w_070_185, w_068_192, w_052_004);
  not1 I070_190(w_070_190, w_038_033);
  or2  I070_191(w_070_191, w_040_309, w_027_143);
  not1 I070_192(w_070_192, w_038_454);
  or2  I070_199(w_070_199, w_047_191, w_049_121);
  or2  I070_205(w_070_205, w_011_634, w_016_005);
  nand2 I070_209(w_070_209, w_010_437, w_027_168);
  and2 I070_210(w_070_210, w_064_297, w_066_370);
  and2 I070_213(w_070_213, w_003_002, w_022_089);
  or2  I070_216(w_070_216, w_055_074, w_033_391);
  or2  I070_220(w_070_220, w_012_040, w_049_110);
  or2  I070_232(w_070_232, w_005_116, w_010_134);
  or2  I070_253(w_070_253, w_047_113, w_050_080);
  not1 I070_256(w_070_256, w_014_127);
  or2  I070_270(w_070_270, w_052_009, w_056_012);
  not1 I070_271(w_070_271, w_060_176);
  or2  I070_280(w_070_280, w_059_012, w_052_002);
  and2 I070_287(w_070_287, w_004_263, w_028_474);
  nand2 I070_289(w_070_289, w_015_045, w_057_025);
  and2 I070_292(w_070_292, w_013_453, w_014_295);
  or2  I070_293(w_070_293, w_003_050, w_044_403);
  and2 I070_294(w_070_294, w_064_136, w_063_111);
  or2  I070_325(w_070_325, w_038_021, w_042_317);
  nand2 I070_327(w_070_327, w_006_075, w_063_034);
  nand2 I070_329(w_070_329, w_042_358, w_066_072);
  and2 I070_330(w_070_330, w_013_455, w_058_541);
  or2  I070_359(w_070_359, w_042_384, w_040_623);
  not1 I070_365(w_070_365, w_052_014);
  nand2 I070_381(w_070_381, w_015_401, w_035_069);
  or2  I070_384(w_070_384, w_058_459, w_057_236);
  nand2 I070_386(w_070_386, w_022_136, w_042_215);
  and2 I070_389(w_070_389, w_011_044, w_044_014);
  not1 I070_390(w_070_390, w_001_034);
  nand2 I070_396(w_070_396, w_042_071, w_034_017);
  or2  I070_404(w_070_404, w_050_120, w_036_386);
  and2 I070_408(w_070_408, w_062_241, w_031_346);
  and2 I070_412(w_070_412, w_060_254, w_056_567);
  and2 I070_424(w_070_424, w_034_060, w_020_091);
  or2  I070_435(w_070_435, w_038_111, w_061_046);
  nand2 I070_437(w_070_437, w_039_197, w_064_241);
  not1 I070_444(w_070_444, w_037_013);
  and2 I070_453(w_070_453, w_045_401, w_012_142);
  nand2 I070_455(w_070_455, w_014_248, w_010_364);
  nand2 I070_459(w_070_459, w_041_036, w_050_046);
  nand2 I070_465(w_070_465, w_045_225, w_026_296);
  nand2 I070_468(w_070_468, w_019_014, w_019_013);
  nand2 I070_471(w_070_471, w_063_160, w_032_191);
  nand2 I070_473(w_070_473, w_064_044, w_057_258);
  nand2 I070_476(w_070_476, w_029_050, w_063_274);
  or2  I070_478(w_070_478, w_020_257, w_061_405);
  nand2 I070_480(w_070_480, w_034_042, w_028_069);
  or2  I070_482(w_070_482, w_051_117, w_033_335);
  and2 I070_486(w_070_486, w_034_008, w_029_094);
  not1 I070_488(w_070_488, w_039_667);
  or2  I070_489(w_070_489, w_063_052, w_066_104);
  nand2 I070_496(w_070_496, w_037_343, w_039_155);
  or2  I070_499(w_070_499, w_012_059, w_020_057);
  nand2 I070_505(w_070_505, w_066_191, w_055_227);
  and2 I070_508(w_070_508, w_030_089, w_022_035);
  and2 I070_510(w_070_510, w_067_334, w_004_059);
  or2  I070_515(w_070_515, w_063_064, w_031_093);
  or2  I070_530(w_070_530, w_026_449, w_031_026);
  not1 I070_542(w_070_542, w_052_031);
  or2  I070_548(w_070_548, w_005_207, w_044_534);
  or2  I070_563(w_070_563, w_030_265, w_068_056);
  not1 I070_568(w_070_568, w_007_276);
  and2 I070_572(w_070_572, w_054_068, w_013_541);
  and2 I070_573(w_070_573, w_047_021, w_033_453);
  not1 I070_579(w_070_579, w_042_024);
  nand2 I071_000(w_071_000, w_036_043, w_055_076);
  not1 I071_001(w_071_001, w_048_011);
  not1 I071_014(w_071_014, w_022_123);
  not1 I071_018(w_071_018, w_041_055);
  and2 I071_020(w_071_020, w_018_039, w_066_356);
  or2  I071_022(w_071_022, w_039_421, w_068_095);
  and2 I071_026(w_071_026, w_021_143, w_019_016);
  or2  I071_029(w_071_029, w_059_459, w_030_378);
  and2 I071_031(w_071_031, w_064_253, w_055_051);
  and2 I071_034(w_071_034, w_050_016, w_018_029);
  nand2 I071_038(w_071_038, w_040_174, w_063_133);
  nand2 I071_045(w_071_045, w_011_594, w_042_109);
  or2  I071_047(w_071_047, w_044_657, w_047_283);
  or2  I071_048(w_071_048, w_020_165, w_007_303);
  or2  I071_052(w_071_052, w_050_446, w_009_550);
  and2 I071_055(w_071_055, w_034_040, w_032_065);
  or2  I071_056(w_071_056, w_059_258, w_055_030);
  or2  I071_058(w_071_058, w_049_280, w_011_167);
  or2  I071_063(w_071_063, w_016_006, w_033_705);
  nand2 I071_066(w_071_066, w_062_739, w_022_093);
  not1 I071_075(w_071_075, w_024_118);
  nand2 I071_076(w_071_076, w_030_151, w_063_014);
  nand2 I071_082(w_071_082, w_007_029, w_030_313);
  nand2 I071_084(w_071_084, w_063_128, w_027_019);
  not1 I071_085(w_071_085, w_023_063);
  nand2 I071_091(w_071_091, w_049_060, w_064_324);
  and2 I071_093(w_071_093, w_049_362, w_010_425);
  or2  I071_094(w_071_094, w_044_366, w_048_009);
  not1 I071_095(w_071_095, w_046_318);
  not1 I071_096(w_071_096, w_051_353);
  and2 I071_097(w_071_097, w_061_158, w_038_298);
  or2  I071_099(w_071_099, w_043_038, w_063_226);
  or2  I071_100(w_071_100, w_040_017, w_034_052);
  nand2 I071_102(w_071_102, w_061_276, w_038_458);
  or2  I071_104(w_071_104, w_069_005, w_043_004);
  nand2 I071_105(w_071_105, w_036_160, w_030_074);
  and2 I071_107(w_071_107, w_003_011, w_007_217);
  or2  I071_109(w_071_109, w_002_330, w_049_220);
  nand2 I071_113(w_071_113, w_030_076, w_008_226);
  not1 I071_121(w_071_121, w_042_327);
  and2 I071_124(w_071_124, w_058_161, w_045_009);
  not1 I071_129(w_071_129, w_040_479);
  not1 I071_138(w_071_138, w_024_218);
  nand2 I071_143(w_071_143, w_022_256, w_039_076);
  or2  I071_144(w_071_144, w_006_248, w_059_260);
  or2  I071_145(w_071_145, w_043_046, w_030_275);
  or2  I071_147(w_071_147, w_022_125, w_028_415);
  not1 I071_148(w_071_148, w_012_322);
  or2  I071_151(w_071_151, w_035_118, w_035_073);
  not1 I071_154(w_071_154, w_022_369);
  and2 I071_155(w_071_155, w_035_076, w_023_034);
  and2 I071_171(w_071_171, w_035_059, w_050_117);
  nand2 I071_173(w_071_173, w_009_268, w_054_199);
  and2 I071_176(w_071_176, w_013_317, w_009_026);
  and2 I071_188(w_071_188, w_014_015, w_012_237);
  and2 I071_205(w_071_205, w_053_018, w_028_088);
  and2 I071_206(w_071_206, w_030_148, w_068_183);
  or2  I071_209(w_071_209, w_050_259, w_067_039);
  or2  I071_213(w_071_213, w_063_514, w_038_121);
  not1 I071_217(w_071_217, w_048_008);
  and2 I071_227(w_071_227, w_068_283, w_011_149);
  nand2 I071_247(w_071_247, w_061_313, w_007_093);
  or2  I071_250(w_071_250, w_018_042, w_070_563);
  or2  I071_252(w_071_252, w_023_070, w_019_013);
  or2  I071_257(w_071_257, w_016_004, w_063_216);
  not1 I071_260(w_071_260, w_012_235);
  nand2 I071_261(w_071_261, w_061_343, w_042_288);
  or2  I071_265(w_071_265, w_061_440, w_039_095);
  nand2 I071_267(w_071_267, w_011_367, w_021_097);
  not1 I071_270(w_071_270, w_059_200);
  nand2 I071_276(w_071_276, w_068_176, w_035_073);
  nand2 I071_277(w_071_277, w_023_093, w_059_647);
  or2  I071_281(w_071_281, w_023_031, w_061_028);
  nand2 I071_284(w_071_284, w_050_427, w_043_012);
  and2 I071_289(w_071_289, w_022_152, w_052_013);
  nand2 I071_294(w_071_294, w_038_067, w_012_075);
  not1 I071_299(w_071_299, w_035_070);
  or2  I071_300(w_071_300, w_006_061, w_044_022);
  and2 I071_302(w_071_302, w_040_013, w_046_630);
  and2 I071_303(w_071_303, w_003_065, w_008_114);
  or2  I071_304(w_071_304, w_043_006, w_030_318);
  and2 I071_305(w_071_305, w_070_112, w_020_124);
  nand2 I071_312(w_071_312, w_056_623, w_047_237);
  or2  I071_315(w_071_315, w_025_141, w_041_647);
  and2 I071_316(w_071_316, w_016_001, w_026_535);
  or2  I071_317(w_071_317, w_050_611, w_066_216);
  nand2 I071_322(w_071_322, w_001_003, w_052_018);
  not1 I072_000(w_072_000, w_040_043);
  not1 I072_001(w_072_001, w_036_083);
  nand2 I072_003(w_072_003, w_014_162, w_038_285);
  not1 I072_005(w_072_005, w_026_322);
  or2  I072_012(w_072_012, w_070_359, w_064_112);
  and2 I072_017(w_072_017, w_048_011, w_031_020);
  and2 I072_020(w_072_020, w_056_400, w_068_011);
  not1 I072_021(w_072_021, w_046_110);
  not1 I072_024(w_072_024, w_000_652);
  or2  I072_034(w_072_034, w_066_170, w_031_156);
  and2 I072_043(w_072_043, w_028_578, w_035_068);
  and2 I072_047(w_072_047, w_011_118, w_059_321);
  or2  I072_048(w_072_048, w_015_099, w_047_207);
  nand2 I072_051(w_072_051, w_056_490, w_011_191);
  not1 I072_052(w_072_052, w_039_032);
  nand2 I072_053(w_072_053, w_048_005, w_008_089);
  not1 I072_054(w_072_054, w_019_013);
  nand2 I072_057(w_072_057, w_022_026, w_004_170);
  and2 I072_058(w_072_058, w_060_257, w_055_097);
  not1 I072_059(w_072_059, w_022_065);
  or2  I072_060(w_072_060, w_015_261, w_002_152);
  nand2 I072_061(w_072_061, w_037_015, w_028_490);
  or2  I072_064(w_072_064, w_060_049, w_065_641);
  not1 I072_067(w_072_067, w_048_016);
  nand2 I072_070(w_072_070, w_022_088, w_036_247);
  nand2 I072_082(w_072_082, w_044_419, w_025_032);
  and2 I072_084(w_072_084, w_044_518, w_065_117);
  not1 I072_090(w_072_090, w_050_069);
  not1 I072_092(w_072_092, w_040_106);
  not1 I072_095(w_072_095, w_042_195);
  not1 I072_096(w_072_096, w_032_148);
  not1 I072_097(w_072_097, w_036_350);
  not1 I072_098(w_072_098, w_013_172);
  and2 I072_101(w_072_101, w_026_670, w_031_165);
  not1 I072_102(w_072_102, w_049_267);
  or2  I072_103(w_072_103, w_024_517, w_060_026);
  nand2 I072_106(w_072_106, w_059_157, w_023_114);
  nand2 I072_107(w_072_107, w_004_288, w_027_117);
  or2  I072_111(w_072_111, w_013_064, w_022_132);
  not1 I072_113(w_072_113, w_008_130);
  or2  I072_114(w_072_114, w_070_148, w_022_123);
  not1 I072_116(w_072_116, w_001_002);
  not1 I072_120(w_072_120, w_002_078);
  nand2 I072_122(w_072_122, w_006_087, w_046_425);
  nand2 I072_123(w_072_123, w_047_215, w_026_160);
  or2  I072_129(w_072_129, w_062_311, w_028_462);
  not1 I072_130(w_072_130, w_055_276);
  or2  I072_131(w_072_131, w_049_271, w_048_018);
  not1 I072_134(w_072_134, w_034_018);
  nand2 I072_135(w_072_135, w_010_571, w_019_004);
  or2  I072_137(w_072_137, w_004_502, w_058_085);
  nand2 I072_143(w_072_143, w_002_301, w_037_172);
  nand2 I072_144(w_072_144, w_059_017, w_030_053);
  nand2 I072_149(w_072_149, w_052_019, w_040_149);
  and2 I072_152(w_072_152, w_059_555, w_035_063);
  nand2 I072_156(w_072_156, w_019_019, w_033_253);
  and2 I072_157(w_072_157, w_041_403, w_066_147);
  nand2 I072_161(w_072_161, w_015_559, w_003_061);
  and2 I072_163(w_072_163, w_067_162, w_041_037);
  or2  I072_165(w_072_165, w_063_156, w_032_044);
  nand2 I072_167(w_072_167, w_013_071, w_062_280);
  or2  I072_169(w_072_169, w_067_263, w_022_206);
  or2  I072_171(w_072_171, w_057_013, w_070_056);
  or2  I072_172(w_072_172, w_031_101, w_009_169);
  nand2 I072_175(w_072_175, w_065_010, w_071_100);
  and2 I072_177(w_072_177, w_061_357, w_053_062);
  or2  I072_178(w_072_178, w_007_427, w_026_648);
  and2 I072_184(w_072_184, w_018_008, w_037_293);
  and2 I072_186(w_072_186, w_060_225, w_023_007);
  nand2 I072_187(w_072_187, w_060_222, w_022_206);
  or2  I072_190(w_072_190, w_054_151, w_061_296);
  not1 I072_195(w_072_195, w_042_185);
  or2  I072_199(w_072_199, w_007_189, w_058_082);
  or2  I072_201(w_072_201, w_011_086, w_002_070);
  not1 I072_208(w_072_208, w_005_092);
  not1 I072_215(w_072_215, w_037_225);
  nand2 I072_232(w_072_232, w_029_051, w_035_066);
  or2  I072_235(w_072_235, w_002_503, w_016_001);
  not1 I072_242(w_072_242, w_007_147);
  not1 I072_260(w_072_260, w_071_095);
  or2  I072_266(w_072_266, w_018_010, w_046_023);
  and2 I072_272(w_072_272, w_004_345, w_069_265);
  not1 I072_278(w_072_278, w_021_147);
  not1 I072_288(w_072_288, w_025_032);
  nand2 I072_289(w_072_289, w_030_332, w_017_319);
  not1 I072_292(w_072_292, w_008_107);
  nand2 I072_295(w_072_295, w_068_076, w_068_357);
  or2  I073_000(w_073_000, w_033_505, w_060_164);
  or2  I073_003(w_073_003, w_032_438, w_072_143);
  or2  I073_009(w_073_009, w_043_009, w_044_367);
  nand2 I073_016(w_073_016, w_067_101, w_018_008);
  and2 I073_017(w_073_017, w_046_619, w_020_076);
  and2 I073_018(w_073_018, w_012_141, w_065_673);
  or2  I073_020(w_073_020, w_010_419, w_026_169);
  nand2 I073_026(w_073_026, w_015_014, w_019_005);
  or2  I073_034(w_073_034, w_036_162, w_053_110);
  and2 I073_037(w_073_037, w_028_012, w_010_632);
  nand2 I073_040(w_073_040, w_048_007, w_007_117);
  nand2 I073_041(w_073_041, w_045_300, w_019_013);
  not1 I073_042(w_073_042, w_043_020);
  or2  I073_043(w_073_043, w_065_270, w_050_408);
  not1 I073_044(w_073_044, w_062_772);
  nand2 I073_049(w_073_049, w_016_006, w_042_356);
  nand2 I073_052(w_073_052, w_033_142, w_070_465);
  nand2 I073_053(w_073_053, w_071_147, w_071_270);
  and2 I073_055(w_073_055, w_030_295, w_068_114);
  and2 I073_068(w_073_068, w_006_068, w_008_175);
  not1 I073_071(w_073_071, w_066_473);
  or2  I073_085(w_073_085, w_052_043, w_066_482);
  and2 I073_088(w_073_088, w_072_242, w_063_083);
  not1 I073_090(w_073_090, w_007_198);
  nand2 I073_095(w_073_095, w_030_076, w_032_160);
  or2  I073_101(w_073_101, w_000_574, w_016_002);
  nand2 I073_114(w_073_114, w_038_317, w_061_056);
  not1 I073_117(w_073_117, w_011_332);
  or2  I073_130(w_073_130, w_045_007, w_017_034);
  or2  I073_139(w_073_139, w_048_012, w_062_173);
  nand2 I073_143(w_073_143, w_058_469, w_014_179);
  or2  I073_150(w_073_150, w_030_104, w_031_555);
  or2  I073_169(w_073_169, w_058_425, w_009_248);
  not1 I073_175(w_073_175, w_003_031);
  not1 I073_183(w_073_183, w_035_050);
  nand2 I073_196(w_073_196, w_009_603, w_042_186);
  nand2 I073_198(w_073_198, w_070_170, w_053_152);
  and2 I073_200(w_073_200, w_049_104, w_003_068);
  and2 I073_203(w_073_203, w_033_057, w_072_054);
  or2  I073_204(w_073_204, w_066_185, w_031_150);
  nand2 I073_209(w_073_209, w_014_073, w_047_051);
  and2 I073_219(w_073_219, w_058_594, w_060_365);
  nand2 I073_224(w_073_224, w_023_078, w_046_057);
  or2  I073_245(w_073_245, w_072_111, w_052_017);
  not1 I073_252(w_073_252, w_051_303);
  or2  I073_253(w_073_253, w_000_263, w_018_004);
  and2 I073_258(w_073_258, w_023_045, w_045_381);
  not1 I073_262(w_073_262, w_019_000);
  not1 I073_284(w_073_284, w_024_209);
  or2  I073_299(w_073_299, w_022_021, w_002_034);
  nand2 I073_326(w_073_326, w_043_007, w_036_386);
  nand2 I073_347(w_073_347, w_039_187, w_063_027);
  or2  I073_363(w_073_363, w_070_123, w_055_000);
  or2  I073_374(w_073_374, w_053_054, w_057_100);
  nand2 I073_379(w_073_379, w_040_409, w_017_260);
  nand2 I073_382(w_073_382, w_018_017, w_042_103);
  nand2 I073_402(w_073_402, w_026_125, w_035_127);
  nand2 I073_404(w_073_404, w_064_335, w_009_325);
  or2  I073_407(w_073_407, w_057_056, w_037_075);
  and2 I073_413(w_073_413, w_040_463, w_032_290);
  or2  I073_419(w_073_419, w_004_199, w_021_021);
  and2 I073_422(w_073_422, w_049_246, w_043_046);
  nand2 I073_428(w_073_428, w_013_529, w_032_151);
  and2 I073_439(w_073_439, w_026_711, w_007_318);
  not1 I073_443(w_073_443, w_043_024);
  nand2 I073_457(w_073_457, w_046_397, w_049_006);
  nand2 I073_463(w_073_463, w_028_304, w_018_007);
  not1 I073_474(w_073_474, w_044_223);
  or2  I073_484(w_073_484, w_057_063, w_015_336);
  or2  I073_489(w_073_489, w_001_013, w_012_201);
  nand2 I073_492(w_073_492, w_029_076, w_002_507);
  nand2 I073_493(w_073_493, w_052_034, w_058_536);
  or2  I073_499(w_073_499, w_057_097, w_056_069);
  not1 I073_503(w_073_503, w_070_050);
  nand2 I073_507(w_073_507, w_062_455, w_008_483);
  and2 I073_512(w_073_512, w_020_400, w_027_020);
  or2  I073_514(w_073_514, w_021_271, w_003_020);
  and2 I073_516(w_073_516, w_035_107, w_024_044);
  nand2 I073_526(w_073_526, w_033_259, w_072_021);
  or2  I073_537(w_073_537, w_041_220, w_062_208);
  nand2 I073_540(w_073_540, w_005_035, w_057_215);
  nand2 I073_554(w_073_554, w_024_216, w_035_006);
  or2  I073_569(w_073_569, w_039_424, w_051_137);
  and2 I073_592(w_073_592, w_005_161, w_053_079);
  nand2 I073_601(w_073_601, w_033_076, w_004_061);
  or2  I073_602(w_073_602, w_007_241, w_055_104);
  not1 I073_605(w_073_605, w_017_408);
  or2  I073_613(w_073_613, w_012_017, w_001_001);
  nand2 I073_621(w_073_621, w_070_031, w_039_621);
  and2 I073_624(w_073_624, w_013_066, w_023_112);
  not1 I073_627(w_073_627, w_049_074);
  not1 I073_632(w_073_632, w_024_434);
  nand2 I073_634(w_073_634, w_004_240, w_017_200);
  not1 I073_649(w_073_649, w_069_197);
  not1 I073_675(w_073_675, w_005_032);
  nand2 I073_687(w_073_687, w_025_021, w_056_525);
  not1 I073_688(w_073_688, w_018_032);
  nand2 I073_691(w_073_691, w_062_081, w_013_153);
  or2  I073_697(w_073_697, w_058_479, w_056_267);
  nand2 I073_714(w_073_714, w_069_075, w_022_337);
  and2 I073_715(w_073_715, w_048_012, w_012_182);
  or2  I073_717(w_073_717, w_016_008, w_010_269);
  not1 I073_722(w_073_722, w_009_602);
  or2  I073_734(w_073_734, w_040_524, w_003_046);
  not1 I073_735(w_073_735, w_001_036);
  and2 I073_740(w_073_740, w_026_115, w_031_015);
  not1 I074_000(w_074_000, w_073_090);
  and2 I074_005(w_074_005, w_061_326, w_006_005);
  nand2 I074_009(w_074_009, w_053_131, w_004_363);
  nand2 I074_012(w_074_012, w_026_706, w_020_107);
  nand2 I074_014(w_074_014, w_051_235, w_013_530);
  or2  I074_023(w_074_023, w_020_139, w_066_202);
  nand2 I074_024(w_074_024, w_006_006, w_047_256);
  nand2 I074_030(w_074_030, w_006_134, w_072_114);
  nand2 I074_032(w_074_032, w_038_240, w_066_007);
  not1 I074_033(w_074_033, w_044_050);
  not1 I074_041(w_074_041, w_035_085);
  nand2 I074_044(w_074_044, w_023_134, w_063_006);
  or2  I074_045(w_074_045, w_031_021, w_007_065);
  and2 I074_046(w_074_046, w_014_280, w_066_578);
  or2  I074_052(w_074_052, w_024_316, w_052_017);
  not1 I074_070(w_074_070, w_008_034);
  or2  I074_077(w_074_077, w_050_008, w_023_166);
  not1 I074_081(w_074_081, w_045_296);
  nand2 I074_099(w_074_099, w_063_503, w_015_210);
  nand2 I074_100(w_074_100, w_071_109, w_065_295);
  and2 I074_104(w_074_104, w_023_079, w_016_000);
  or2  I074_105(w_074_105, w_069_165, w_064_286);
  and2 I074_107(w_074_107, w_014_067, w_064_038);
  not1 I074_108(w_074_108, w_053_090);
  and2 I074_111(w_074_111, w_065_449, w_016_007);
  or2  I074_114(w_074_114, w_015_557, w_013_092);
  not1 I074_117(w_074_117, w_033_244);
  not1 I074_124(w_074_124, w_055_104);
  and2 I074_127(w_074_127, w_058_647, w_034_006);
  nand2 I074_128(w_074_128, w_016_007, w_008_402);
  nand2 I074_141(w_074_141, w_018_021, w_021_072);
  not1 I074_144(w_074_144, w_071_317);
  nand2 I074_152(w_074_152, w_043_047, w_021_073);
  not1 I074_153(w_074_153, w_058_683);
  and2 I074_154(w_074_154, w_063_302, w_007_477);
  and2 I074_157(w_074_157, w_020_511, w_019_015);
  or2  I074_159(w_074_159, w_025_126, w_017_098);
  and2 I074_166(w_074_166, w_027_058, w_024_097);
  not1 I074_168(w_074_168, w_025_155);
  or2  I074_169(w_074_169, w_003_077, w_023_138);
  or2  I074_175(w_074_175, w_039_466, w_057_099);
  nand2 I074_176(w_074_176, w_006_152, w_050_123);
  and2 I074_177(w_074_177, w_066_093, w_002_358);
  or2  I074_179(w_074_179, w_041_228, w_011_322);
  or2  I074_182(w_074_182, w_073_363, w_058_645);
  or2  I074_184(w_074_184, w_027_173, w_017_135);
  nand2 I074_186(w_074_186, w_027_028, w_000_013);
  and2 I074_190(w_074_190, w_008_429, w_017_613);
  or2  I074_193(w_074_193, w_055_279, w_005_127);
  not1 I074_194(w_074_194, w_016_001);
  nand2 I074_196(w_074_196, w_006_183, w_002_312);
  nand2 I074_200(w_074_200, w_016_005, w_013_407);
  and2 I074_201(w_074_201, w_036_307, w_010_653);
  not1 I074_209(w_074_209, w_072_177);
  nand2 I074_210(w_074_210, w_032_121, w_027_130);
  and2 I074_215(w_074_215, w_046_389, w_035_114);
  or2  I074_218(w_074_218, w_006_100, w_021_000);
  not1 I074_221(w_074_221, w_071_322);
  not1 I074_227(w_074_227, w_071_261);
  nand2 I074_231(w_074_231, w_036_449, w_029_081);
  or2  I074_232(w_074_232, w_028_182, w_035_064);
  and2 I074_233(w_074_233, w_052_015, w_030_355);
  not1 I074_243(w_074_243, w_033_282);
  or2  I074_250(w_074_250, w_071_018, w_016_002);
  or2  I074_251(w_074_251, w_051_215, w_053_092);
  and2 I074_252(w_074_252, w_016_000, w_014_081);
  not1 I074_254(w_074_254, w_062_761);
  and2 I074_256(w_074_256, w_037_336, w_073_130);
  nand2 I074_258(w_074_258, w_013_064, w_045_245);
  nand2 I074_259(w_074_259, w_038_055, w_025_061);
  not1 I074_265(w_074_265, w_017_050);
  not1 I074_277(w_074_277, w_001_012);
  and2 I074_287(w_074_287, w_055_038, w_063_225);
  and2 I074_288(w_074_288, w_033_116, w_030_191);
  and2 I074_293(w_074_293, w_035_120, w_044_115);
  not1 I074_294(w_074_294, w_011_049);
  and2 I074_296(w_074_296, w_039_160, w_012_017);
  or2  I074_297(w_074_297, w_064_142, w_053_081);
  nand2 I074_300(w_074_300, w_052_030, w_070_010);
  not1 I074_303(w_074_303, w_025_123);
  and2 I074_309(w_074_309, w_033_026, w_069_192);
  not1 I074_313(w_074_313, w_004_444);
  or2  I074_317(w_074_317, w_061_477, w_006_017);
  or2  I074_320(w_074_320, w_016_007, w_007_240);
  and2 I074_321(w_074_321, w_046_194, w_024_481);
  and2 I074_322(w_074_322, w_059_354, w_002_025);
  or2  I074_327(w_074_327, w_026_297, w_071_138);
  nand2 I074_331(w_074_331, w_056_007, w_001_034);
  or2  I074_334(w_074_334, w_024_329, w_059_178);
  not1 I074_337(w_074_337, w_043_003);
  or2  I074_340(w_074_340, w_049_153, w_040_031);
  nand2 I074_342(w_074_342, w_048_003, w_047_021);
  not1 I074_343(w_074_343, w_021_037);
  and2 I074_344(w_074_344, w_043_022, w_027_148);
  nand2 I074_345(w_074_345, w_049_165, w_008_509);
  or2  I074_348(w_074_348, w_008_591, w_067_383);
  or2  I074_351(w_074_351, w_069_159, w_026_004);
  and2 I074_360(w_074_360, w_042_002, w_016_003);
  nand2 I074_363(w_074_363, w_025_056, w_068_000);
  and2 I074_370(w_074_370, w_004_039, w_060_189);
  and2 I074_374(w_074_374, w_024_277, w_026_305);
  nand2 I074_375(w_074_375, w_039_032, w_002_181);
  nand2 I075_000(w_075_000, w_045_389, w_049_347);
  nand2 I075_001(w_075_001, w_061_408, w_018_003);
  not1 I075_002(w_075_002, w_001_005);
  nand2 I075_005(w_075_005, w_064_286, w_058_696);
  not1 I075_007(w_075_007, w_037_096);
  and2 I075_009(w_075_009, w_043_034, w_063_064);
  and2 I075_010(w_075_010, w_003_010, w_067_013);
  not1 I075_011(w_075_011, w_029_113);
  nand2 I075_013(w_075_013, w_032_064, w_073_253);
  or2  I075_014(w_075_014, w_021_043, w_047_323);
  nand2 I075_016(w_075_016, w_027_165, w_067_381);
  or2  I075_018(w_075_018, w_012_187, w_011_071);
  and2 I075_019(w_075_019, w_031_281, w_011_013);
  not1 I075_020(w_075_020, w_022_202);
  nand2 I075_023(w_075_023, w_057_102, w_008_544);
  not1 I075_024(w_075_024, w_001_029);
  and2 I075_025(w_075_025, w_014_229, w_047_141);
  or2  I075_027(w_075_027, w_061_179, w_057_062);
  or2  I075_030(w_075_030, w_040_005, w_025_143);
  and2 I075_032(w_075_032, w_051_080, w_048_016);
  not1 I075_033(w_075_033, w_008_145);
  or2  I075_034(w_075_034, w_042_035, w_016_005);
  nand2 I075_037(w_075_037, w_036_182, w_017_341);
  and2 I075_039(w_075_039, w_055_036, w_063_050);
  or2  I075_043(w_075_043, w_050_021, w_001_020);
  not1 I075_044(w_075_044, w_018_039);
  or2  I075_045(w_075_045, w_049_012, w_047_155);
  and2 I075_046(w_075_046, w_027_145, w_061_255);
  not1 I075_047(w_075_047, w_057_000);
  not1 I075_049(w_075_049, w_055_239);
  or2  I075_050(w_075_050, w_062_194, w_027_006);
  nand2 I075_052(w_075_052, w_014_066, w_034_018);
  nand2 I075_053(w_075_053, w_062_250, w_037_071);
  not1 I075_054(w_075_054, w_052_026);
  nand2 I075_055(w_075_055, w_007_200, w_022_074);
  or2  I075_058(w_075_058, w_055_168, w_023_154);
  nand2 I075_061(w_075_061, w_020_054, w_015_675);
  or2  I075_062(w_075_062, w_022_017, w_074_104);
  not1 I075_063(w_075_063, w_053_108);
  not1 I075_065(w_075_065, w_025_021);
  and2 I075_067(w_075_067, w_000_154, w_016_005);
  not1 I075_069(w_075_069, w_069_068);
  nand2 I075_071(w_075_071, w_074_177, w_007_103);
  or2  I075_072(w_075_072, w_058_427, w_001_002);
  not1 I075_074(w_075_074, w_018_017);
  not1 I075_076(w_075_076, w_015_068);
  and2 I075_077(w_075_077, w_010_688, w_025_294);
  or2  I075_078(w_075_078, w_049_254, w_010_128);
  or2  I075_079(w_075_079, w_070_453, w_046_372);
  and2 I075_083(w_075_083, w_074_288, w_058_159);
  and2 I075_087(w_075_087, w_022_283, w_046_121);
  and2 I075_091(w_075_091, w_048_011, w_019_016);
  or2  I075_096(w_075_096, w_060_395, w_028_586);
  and2 I075_097(w_075_097, w_045_274, w_000_120);
  not1 I075_100(w_075_100, w_047_047);
  and2 I075_101(w_075_101, w_001_033, w_032_579);
  not1 I075_105(w_075_105, w_045_280);
  and2 I075_109(w_075_109, w_006_009, w_067_113);
  nand2 I075_111(w_075_111, w_012_004, w_026_608);
  nand2 I075_113(w_075_113, w_053_040, w_002_639);
  not1 I075_114(w_075_114, w_024_456);
  not1 I075_116(w_075_116, w_057_268);
  or2  I075_117(w_075_117, w_070_486, w_048_014);
  nand2 I075_118(w_075_118, w_066_125, w_018_035);
  or2  I075_120(w_075_120, w_062_168, w_041_676);
  or2  I075_127(w_075_127, w_067_141, w_044_139);
  or2  I075_128(w_075_128, w_061_066, w_009_006);
  or2  I075_132(w_075_132, w_017_066, w_032_160);
  nand2 I075_133(w_075_133, w_033_730, w_036_354);
  or2  I075_134(w_075_134, w_014_169, w_012_023);
  and2 I075_135(w_075_135, w_062_224, w_068_133);
  not1 I075_136(w_075_136, w_002_372);
  nand2 I075_137(w_075_137, w_066_080, w_043_033);
  and2 I075_138(w_075_138, w_036_052, w_035_003);
  and2 I075_139(w_075_139, w_044_019, w_004_128);
  and2 I075_140(w_075_140, w_018_032, w_069_209);
  and2 I075_141(w_075_141, w_058_135, w_025_186);
  nand2 I075_144(w_075_144, w_016_001, w_022_152);
  not1 I075_145(w_075_145, w_034_004);
  or2  I075_147(w_075_147, w_059_722, w_001_020);
  nand2 I075_148(w_075_148, w_011_026, w_001_013);
  and2 I075_152(w_075_152, w_057_150, w_060_299);
  nand2 I075_153(w_075_153, w_068_342, w_067_094);
  nand2 I075_155(w_075_155, w_047_040, w_000_293);
  or2  I075_157(w_075_159, w_065_174, w_075_158);
  or2  I075_158(w_075_160, w_051_196, w_075_159);
  and2 I075_159(w_075_161, w_075_160, w_005_107);
  or2  I075_160(w_075_158, w_050_226, w_075_161);
  not1 I076_014(w_076_014, w_069_158);
  nand2 I076_015(w_076_015, w_045_331, w_057_049);
  or2  I076_033(w_076_033, w_010_375, w_018_018);
  not1 I076_036(w_076_036, w_004_004);
  or2  I076_040(w_076_040, w_073_016, w_019_013);
  nand2 I076_043(w_076_043, w_001_010, w_073_175);
  not1 I076_046(w_076_046, w_007_000);
  not1 I076_050(w_076_050, w_038_148);
  not1 I076_052(w_076_052, w_067_250);
  or2  I076_060(w_076_060, w_061_257, w_034_062);
  nand2 I076_062(w_076_062, w_070_455, w_017_086);
  not1 I076_070(w_076_070, w_003_050);
  nand2 I076_072(w_076_072, w_004_293, w_030_168);
  and2 I076_074(w_076_074, w_053_149, w_027_151);
  and2 I076_087(w_076_087, w_030_252, w_059_507);
  not1 I076_091(w_076_091, w_041_298);
  or2  I076_098(w_076_098, w_023_114, w_047_177);
  or2  I076_099(w_076_099, w_036_314, w_050_385);
  and2 I076_102(w_076_102, w_062_178, w_034_054);
  or2  I076_104(w_076_104, w_041_037, w_037_300);
  not1 I076_107(w_076_107, w_023_060);
  and2 I076_108(w_076_108, w_062_378, w_042_409);
  and2 I076_111(w_076_111, w_068_092, w_053_047);
  not1 I076_115(w_076_115, w_032_418);
  and2 I076_130(w_076_130, w_047_263, w_009_035);
  and2 I076_134(w_076_134, w_011_373, w_041_102);
  and2 I076_136(w_076_136, w_040_312, w_052_031);
  nand2 I076_137(w_076_137, w_061_323, w_031_088);
  and2 I076_140(w_076_140, w_018_014, w_008_032);
  nand2 I076_145(w_076_145, w_060_324, w_052_007);
  not1 I076_157(w_076_157, w_020_370);
  or2  I076_158(w_076_158, w_062_776, w_052_041);
  nand2 I076_161(w_076_161, w_021_192, w_010_004);
  and2 I076_162(w_076_162, w_065_038, w_053_069);
  or2  I076_168(w_076_168, w_023_054, w_008_568);
  and2 I076_173(w_076_173, w_043_018, w_066_123);
  not1 I076_181(w_076_181, w_035_114);
  not1 I076_182(w_076_182, w_061_434);
  nand2 I076_183(w_076_183, w_062_131, w_069_194);
  or2  I076_197(w_076_197, w_058_224, w_012_075);
  nand2 I076_200(w_076_200, w_054_510, w_051_006);
  and2 I076_201(w_076_201, w_062_734, w_035_122);
  and2 I076_206(w_076_206, w_045_401, w_003_009);
  or2  I076_209(w_076_209, w_042_201, w_011_320);
  nand2 I076_210(w_076_210, w_062_796, w_022_138);
  and2 I076_218(w_076_218, w_000_614, w_057_061);
  and2 I076_220(w_076_220, w_049_411, w_000_783);
  not1 I076_221(w_076_221, w_031_179);
  or2  I076_233(w_076_233, w_031_188, w_060_033);
  not1 I076_237(w_076_237, w_037_188);
  or2  I076_240(w_076_240, w_046_532, w_046_143);
  or2  I076_241(w_076_241, w_003_049, w_073_697);
  and2 I076_255(w_076_255, w_016_006, w_038_495);
  not1 I076_258(w_076_258, w_016_006);
  nand2 I076_262(w_076_262, w_055_267, w_005_132);
  and2 I076_277(w_076_277, w_071_252, w_014_031);
  not1 I076_292(w_076_292, w_012_239);
  nand2 I076_294(w_076_294, w_027_125, w_062_017);
  not1 I076_295(w_076_295, w_019_008);
  not1 I076_296(w_076_296, w_032_526);
  and2 I076_300(w_076_300, w_027_111, w_062_093);
  and2 I076_311(w_076_311, w_008_659, w_057_241);
  and2 I076_319(w_076_319, w_075_109, w_049_171);
  not1 I076_321(w_076_321, w_038_489);
  not1 I076_326(w_076_326, w_001_008);
  nand2 I076_327(w_076_327, w_018_007, w_019_009);
  and2 I076_334(w_076_334, w_005_055, w_050_186);
  or2  I076_345(w_076_345, w_063_417, w_053_037);
  nand2 I076_347(w_076_347, w_043_020, w_033_111);
  nand2 I076_351(w_076_351, w_031_445, w_048_012);
  nand2 I076_362(w_076_362, w_031_556, w_022_380);
  nand2 I076_364(w_076_364, w_038_099, w_031_150);
  and2 I076_375(w_076_375, w_009_574, w_027_065);
  or2  I076_405(w_076_405, w_003_080, w_022_386);
  not1 I076_418(w_076_418, w_025_152);
  or2  I076_421(w_076_421, w_063_029, w_002_308);
  or2  I076_432(w_076_432, w_009_449, w_021_064);
  and2 I076_447(w_076_447, w_062_307, w_065_359);
  and2 I076_458(w_076_458, w_029_023, w_051_301);
  and2 I076_459(w_076_459, w_041_714, w_018_044);
  and2 I076_461(w_076_461, w_042_385, w_003_050);
  and2 I076_476(w_076_476, w_029_053, w_073_443);
  not1 I076_479(w_076_479, w_008_347);
  nand2 I076_489(w_076_489, w_031_120, w_039_152);
  or2  I076_492(w_076_494, w_070_548, w_076_493);
  nand2 I076_493(w_076_495, w_059_186, w_076_494);
  not1 I076_494(w_076_496, w_076_495);
  nand2 I076_495(w_076_497, w_076_496, w_040_225);
  nand2 I076_496(w_076_498, w_012_108, w_076_497);
  and2 I076_497(w_076_499, w_076_498, w_056_686);
  or2  I076_498(w_076_500, w_009_415, w_076_499);
  and2 I076_499(w_076_501, w_076_500, w_045_160);
  and2 I076_500(w_076_502, w_047_311, w_076_501);
  or2  I076_501(w_076_493, w_076_502, w_023_144);
  and2 I077_000(w_077_000, w_022_104, w_042_328);
  not1 I077_011(w_077_011, w_004_024);
  not1 I077_019(w_077_019, w_055_095);
  or2  I077_021(w_077_021, w_057_123, w_045_003);
  nand2 I077_022(w_077_022, w_020_098, w_038_147);
  and2 I077_026(w_077_026, w_002_460, w_001_019);
  and2 I077_029(w_077_029, w_074_023, w_027_054);
  not1 I077_032(w_077_032, w_047_038);
  and2 I077_035(w_077_035, w_054_502, w_010_060);
  not1 I077_039(w_077_039, w_009_000);
  nand2 I077_043(w_077_043, w_011_103, w_005_251);
  not1 I077_044(w_077_044, w_064_233);
  not1 I077_048(w_077_048, w_055_043);
  and2 I077_052(w_077_052, w_072_021, w_051_053);
  nand2 I077_054(w_077_054, w_009_432, w_021_216);
  or2  I077_057(w_077_057, w_023_123, w_023_076);
  not1 I077_058(w_077_058, w_015_332);
  or2  I077_060(w_077_060, w_035_085, w_058_253);
  nand2 I077_086(w_077_086, w_045_191, w_059_090);
  nand2 I077_089(w_077_089, w_040_660, w_066_273);
  not1 I077_091(w_077_091, w_041_016);
  not1 I077_099(w_077_099, w_062_185);
  nand2 I077_102(w_077_102, w_056_390, w_051_188);
  or2  I077_107(w_077_107, w_024_098, w_036_217);
  and2 I077_110(w_077_110, w_021_094, w_072_137);
  not1 I077_123(w_077_123, w_061_004);
  or2  I077_127(w_077_127, w_069_071, w_036_082);
  and2 I077_133(w_077_133, w_073_034, w_020_350);
  not1 I077_140(w_077_140, w_013_519);
  nand2 I077_150(w_077_150, w_073_407, w_033_613);
  or2  I077_151(w_077_151, w_022_155, w_031_145);
  not1 I077_152(w_077_152, w_027_117);
  and2 I077_165(w_077_165, w_071_076, w_068_301);
  and2 I077_166(w_077_166, w_069_087, w_017_425);
  nand2 I077_176(w_077_176, w_045_181, w_002_191);
  nand2 I077_178(w_077_178, w_003_053, w_019_007);
  nand2 I077_185(w_077_185, w_027_078, w_039_448);
  nand2 I077_209(w_077_209, w_044_681, w_053_132);
  not1 I077_210(w_077_210, w_065_056);
  or2  I077_223(w_077_223, w_034_067, w_042_066);
  nand2 I077_232(w_077_232, w_064_121, w_008_041);
  and2 I077_240(w_077_240, w_006_122, w_049_070);
  and2 I077_242(w_077_242, w_053_076, w_001_001);
  or2  I077_245(w_077_245, w_060_341, w_061_374);
  and2 I077_251(w_077_251, w_062_503, w_008_240);
  and2 I077_254(w_077_254, w_045_228, w_043_006);
  not1 I077_262(w_077_262, w_065_126);
  not1 I077_272(w_077_272, w_063_245);
  or2  I077_282(w_077_282, w_032_167, w_057_025);
  or2  I077_286(w_077_286, w_015_183, w_054_066);
  and2 I077_289(w_077_289, w_076_182, w_052_023);
  not1 I077_290(w_077_290, w_062_612);
  nand2 I077_292(w_077_292, w_063_025, w_025_007);
  or2  I077_310(w_077_310, w_031_107, w_058_555);
  not1 I077_313(w_077_313, w_076_197);
  or2  I077_315(w_077_315, w_040_193, w_043_017);
  or2  I077_321(w_077_321, w_061_162, w_074_024);
  and2 I077_344(w_077_344, w_007_081, w_017_256);
  or2  I077_361(w_077_361, w_025_134, w_013_462);
  not1 I077_372(w_077_372, w_023_087);
  nand2 I077_378(w_077_378, w_014_130, w_073_114);
  or2  I077_382(w_077_382, w_075_050, w_009_455);
  or2  I077_385(w_077_385, w_059_517, w_071_205);
  or2  I077_398(w_077_398, w_030_288, w_030_396);
  nand2 I077_401(w_077_401, w_015_165, w_007_235);
  not1 I077_409(w_077_409, w_023_035);
  not1 I077_412(w_077_412, w_032_180);
  and2 I077_420(w_077_420, w_019_012, w_065_572);
  nand2 I077_424(w_077_424, w_040_427, w_002_121);
  or2  I077_431(w_077_431, w_004_000, w_066_586);
  and2 I077_440(w_077_440, w_048_015, w_019_019);
  not1 I077_444(w_077_444, w_059_002);
  and2 I077_479(w_077_479, w_054_061, w_061_192);
  and2 I077_481(w_077_481, w_020_180, w_042_226);
  and2 I077_483(w_077_483, w_001_004, w_054_164);
  not1 I077_488(w_077_488, w_007_226);
  and2 I077_500(w_077_500, w_007_069, w_014_178);
  or2  I077_519(w_077_519, w_059_166, w_064_133);
  nand2 I077_522(w_077_522, w_052_034, w_073_040);
  nand2 I077_540(w_077_540, w_067_099, w_068_030);
  nand2 I077_551(w_077_551, w_064_308, w_009_129);
  or2  I077_552(w_077_552, w_070_270, w_034_021);
  and2 I077_558(w_077_558, w_062_512, w_053_091);
  or2  I077_560(w_077_560, w_023_157, w_039_173);
  or2  I077_577(w_077_577, w_068_210, w_036_272);
  not1 I077_586(w_077_586, w_002_441);
  and2 I077_590(w_077_590, w_030_021, w_017_043);
  nand2 I077_592(w_077_592, w_000_305, w_050_050);
  nand2 I077_597(w_077_597, w_019_007, w_053_041);
  or2  I077_601(w_077_601, w_028_536, w_007_337);
  or2  I077_610(w_077_610, w_059_183, w_064_100);
  or2  I077_619(w_077_619, w_042_162, w_074_317);
  or2  I077_626(w_077_626, w_001_034, w_026_630);
  not1 I077_629(w_077_631, w_077_630);
  nand2 I077_630(w_077_632, w_019_004, w_077_631);
  nand2 I077_631(w_077_633, w_064_265, w_077_632);
  and2 I077_632(w_077_634, w_077_633, w_047_045);
  nand2 I077_633(w_077_630, w_023_055, w_077_634);
  and2 I078_004(w_078_004, w_054_439, w_012_007);
  or2  I078_013(w_078_013, w_005_129, w_035_125);
  not1 I078_015(w_078_015, w_052_020);
  nand2 I078_016(w_078_016, w_006_199, w_051_330);
  nand2 I078_024(w_078_024, w_054_279, w_067_333);
  not1 I078_033(w_078_033, w_065_295);
  or2  I078_037(w_078_037, w_030_296, w_055_084);
  not1 I078_038(w_078_038, w_006_235);
  or2  I078_039(w_078_039, w_073_000, w_028_182);
  and2 I078_043(w_078_043, w_057_025, w_064_184);
  or2  I078_044(w_078_044, w_049_237, w_053_034);
  and2 I078_050(w_078_050, w_054_557, w_050_103);
  not1 I078_053(w_078_053, w_075_141);
  not1 I078_055(w_078_055, w_020_519);
  not1 I078_056(w_078_056, w_049_240);
  not1 I078_058(w_078_058, w_003_075);
  and2 I078_061(w_078_061, w_024_257, w_042_094);
  nand2 I078_063(w_078_063, w_077_289, w_008_435);
  not1 I078_070(w_078_070, w_059_455);
  and2 I078_078(w_078_078, w_029_108, w_019_015);
  or2  I078_080(w_078_080, w_059_439, w_031_008);
  nand2 I078_083(w_078_083, w_057_018, w_037_203);
  or2  I078_084(w_078_084, w_005_296, w_026_477);
  and2 I078_089(w_078_089, w_051_159, w_072_005);
  nand2 I078_093(w_078_093, w_067_352, w_058_090);
  not1 I078_101(w_078_101, w_026_508);
  or2  I078_102(w_078_102, w_059_052, w_009_013);
  and2 I078_103(w_078_103, w_038_144, w_070_006);
  not1 I078_104(w_078_104, w_055_078);
  or2  I078_106(w_078_106, w_066_463, w_061_199);
  not1 I078_112(w_078_112, w_038_501);
  nand2 I078_121(w_078_121, w_015_606, w_017_508);
  nand2 I078_122(w_078_122, w_070_096, w_057_028);
  and2 I078_130(w_078_130, w_050_024, w_068_306);
  not1 I078_142(w_078_142, w_036_327);
  not1 I078_144(w_078_144, w_014_094);
  not1 I078_145(w_078_145, w_059_340);
  and2 I078_149(w_078_149, w_042_155, w_027_024);
  or2  I078_150(w_078_150, w_036_257, w_011_011);
  and2 I078_152(w_078_152, w_063_086, w_012_108);
  or2  I078_166(w_078_166, w_008_709, w_064_306);
  or2  I078_168(w_078_168, w_075_132, w_043_006);
  or2  I078_169(w_078_169, w_028_058, w_044_201);
  nand2 I078_170(w_078_170, w_052_022, w_039_073);
  not1 I078_177(w_078_177, w_066_518);
  not1 I078_183(w_078_183, w_048_011);
  or2  I078_188(w_078_188, w_065_097, w_049_112);
  nand2 I078_195(w_078_195, w_064_094, w_061_473);
  and2 I078_200(w_078_200, w_058_274, w_002_039);
  and2 I078_208(w_078_208, w_032_309, w_006_132);
  not1 I078_213(w_078_213, w_071_093);
  nand2 I078_225(w_078_225, w_000_279, w_055_262);
  or2  I078_229(w_078_229, w_052_014, w_052_013);
  nand2 I078_230(w_078_230, w_032_228, w_050_037);
  nand2 I078_251(w_078_251, w_072_101, w_067_140);
  nand2 I078_306(w_078_306, w_038_297, w_000_265);
  or2  I078_318(w_078_318, w_032_092, w_044_209);
  or2  I078_329(w_078_329, w_074_277, w_031_026);
  and2 I078_345(w_078_345, w_025_265, w_039_600);
  nand2 I078_349(w_078_349, w_051_406, w_040_072);
  and2 I078_366(w_078_366, w_056_049, w_050_611);
  or2  I078_379(w_078_379, w_036_072, w_047_251);
  and2 I078_381(w_078_381, w_072_169, w_039_218);
  not1 I078_396(w_078_396, w_047_199);
  or2  I078_401(w_078_401, w_071_082, w_024_535);
  not1 I078_416(w_078_416, w_069_049);
  or2  I078_421(w_078_421, w_026_515, w_000_671);
  not1 I078_428(w_078_428, w_074_154);
  not1 I078_429(w_078_429, w_023_181);
  nand2 I078_434(w_078_434, w_064_115, w_054_098);
  and2 I078_441(w_078_441, w_014_286, w_028_090);
  nand2 I078_445(w_078_445, w_028_003, w_076_108);
  not1 I078_446(w_078_446, w_041_334);
  not1 I078_464(w_078_464, w_021_088);
  or2  I078_465(w_078_465, w_062_784, w_020_158);
  not1 I078_475(w_078_475, w_041_241);
  nand2 I078_497(w_078_497, w_031_596, w_002_321);
  not1 I078_511(w_078_511, w_069_174);
  or2  I078_514(w_078_514, w_047_155, w_020_049);
  not1 I078_520(w_078_520, w_009_395);
  nand2 I078_560(w_078_560, w_025_115, w_073_041);
  or2  I078_566(w_078_566, w_055_297, w_047_396);
  and2 I078_571(w_078_571, w_015_652, w_023_070);
  not1 I078_573(w_078_573, w_003_037);
  nand2 I078_588(w_078_588, w_049_101, w_010_187);
  and2 I078_597(w_078_597, w_058_602, w_072_113);
  nand2 I079_000(w_079_000, w_054_013, w_026_067);
  or2  I079_001(w_079_001, w_069_228, w_014_112);
  or2  I079_002(w_079_002, w_043_022, w_007_077);
  nand2 I079_003(w_079_003, w_018_041, w_035_057);
  and2 I079_004(w_079_004, w_025_081, w_049_024);
  not1 I079_005(w_079_005, w_076_476);
  nand2 I079_007(w_079_007, w_030_331, w_041_579);
  and2 I079_008(w_079_008, w_030_037, w_052_028);
  nand2 I079_010(w_079_010, w_007_033, w_029_096);
  nand2 I079_012(w_079_012, w_019_014, w_049_299);
  not1 I079_015(w_079_015, w_031_120);
  or2  I079_016(w_079_016, w_066_063, w_001_012);
  nand2 I079_017(w_079_017, w_063_190, w_007_340);
  not1 I079_018(w_079_018, w_035_055);
  nand2 I079_020(w_079_020, w_015_097, w_017_115);
  and2 I079_021(w_079_021, w_015_676, w_024_367);
  not1 I079_022(w_079_022, w_031_487);
  nand2 I079_023(w_079_023, w_018_015, w_046_334);
  not1 I079_024(w_079_024, w_030_097);
  and2 I079_025(w_079_025, w_075_101, w_076_334);
  and2 I079_027(w_079_027, w_060_300, w_019_015);
  and2 I079_028(w_079_028, w_009_166, w_031_092);
  not1 I079_029(w_079_029, w_062_131);
  or2  I079_030(w_079_030, w_055_066, w_060_216);
  and2 I079_031(w_079_031, w_065_343, w_047_362);
  not1 I079_033(w_079_033, w_028_113);
  and2 I079_035(w_079_035, w_045_001, w_017_529);
  and2 I079_036(w_079_036, w_020_103, w_059_538);
  or2  I079_037(w_079_037, w_035_028, w_053_048);
  or2  I079_038(w_079_038, w_040_592, w_046_248);
  not1 I079_039(w_079_039, w_041_496);
  or2  I079_040(w_079_040, w_070_396, w_009_364);
  or2  I079_041(w_079_041, w_004_309, w_049_397);
  not1 I079_043(w_079_043, w_037_234);
  nand2 I079_044(w_079_044, w_003_080, w_002_360);
  or2  I079_045(w_079_045, w_024_577, w_040_101);
  and2 I079_047(w_079_047, w_023_018, w_078_144);
  or2  I079_048(w_079_048, w_004_005, w_021_069);
  nand2 I079_050(w_079_050, w_064_226, w_038_196);
  and2 I079_051(w_079_051, w_039_505, w_043_047);
  not1 I079_052(w_079_052, w_059_559);
  not1 I079_053(w_079_053, w_012_047);
  not1 I079_054(w_079_054, w_011_634);
  or2  I079_055(w_079_055, w_078_379, w_037_021);
  not1 I079_056(w_079_056, w_012_136);
  and2 I079_057(w_079_057, w_070_060, w_056_058);
  or2  I079_058(w_079_058, w_030_317, w_011_396);
  or2  I079_059(w_079_059, w_052_000, w_007_389);
  nand2 I079_060(w_079_060, w_050_008, w_035_066);
  nand2 I079_062(w_079_062, w_020_088, w_042_309);
  or2  I080_003(w_080_003, w_073_526, w_032_097);
  not1 I080_007(w_080_007, w_065_032);
  and2 I080_011(w_080_011, w_015_011, w_017_022);
  not1 I080_013(w_080_013, w_035_035);
  nand2 I080_019(w_080_019, w_036_062, w_030_151);
  and2 I080_023(w_080_023, w_053_081, w_043_047);
  not1 I080_029(w_080_029, w_022_385);
  or2  I080_032(w_080_032, w_028_144, w_012_001);
  and2 I080_033(w_080_033, w_043_019, w_071_094);
  nand2 I080_044(w_080_044, w_076_326, w_059_444);
  or2  I080_052(w_080_052, w_051_208, w_026_683);
  or2  I080_053(w_080_053, w_012_004, w_074_201);
  or2  I080_054(w_080_054, w_079_062, w_023_152);
  or2  I080_063(w_080_063, w_064_255, w_050_406);
  not1 I080_065(w_080_065, w_016_006);
  or2  I080_076(w_080_076, w_024_305, w_046_525);
  not1 I080_079(w_080_079, w_009_340);
  not1 I080_080(w_080_080, w_022_083);
  or2  I080_085(w_080_085, w_022_111, w_031_366);
  or2  I080_086(w_080_086, w_061_298, w_019_008);
  and2 I080_096(w_080_096, w_049_003, w_009_423);
  or2  I080_098(w_080_098, w_058_123, w_062_440);
  not1 I080_113(w_080_113, w_016_008);
  and2 I080_118(w_080_118, w_018_019, w_071_317);
  nand2 I080_120(w_080_120, w_051_317, w_072_095);
  or2  I080_131(w_080_131, w_078_213, w_014_116);
  not1 I080_132(w_080_132, w_037_070);
  not1 I080_134(w_080_134, w_008_409);
  nand2 I080_138(w_080_138, w_010_059, w_010_260);
  and2 I080_153(w_080_153, w_048_018, w_007_339);
  or2  I080_154(w_080_154, w_042_312, w_004_125);
  and2 I080_158(w_080_158, w_042_286, w_033_660);
  not1 I080_159(w_080_159, w_039_231);
  nand2 I080_162(w_080_162, w_073_740, w_041_355);
  nand2 I080_171(w_080_171, w_078_429, w_047_155);
  not1 I080_173(w_080_173, w_075_114);
  and2 I080_176(w_080_176, w_074_259, w_073_252);
  not1 I080_182(w_080_182, w_028_550);
  nand2 I080_183(w_080_183, w_040_607, w_069_241);
  not1 I080_185(w_080_185, w_000_179);
  not1 I080_186(w_080_186, w_022_172);
  or2  I080_192(w_080_192, w_065_654, w_052_002);
  not1 I080_202(w_080_202, w_011_011);
  not1 I080_212(w_080_212, w_076_206);
  or2  I080_213(w_080_213, w_036_138, w_072_120);
  not1 I080_222(w_080_222, w_031_040);
  and2 I080_225(w_080_225, w_054_004, w_026_072);
  nand2 I080_230(w_080_230, w_044_521, w_013_160);
  not1 I080_231(w_080_231, w_077_558);
  nand2 I080_233(w_080_233, w_073_540, w_023_068);
  and2 I080_237(w_080_237, w_026_059, w_001_008);
  nand2 I080_238(w_080_238, w_079_000, w_009_375);
  not1 I080_245(w_080_245, w_001_008);
  or2  I080_249(w_080_249, w_076_489, w_070_117);
  nand2 I080_251(w_080_251, w_066_111, w_011_216);
  not1 I080_255(w_080_255, w_059_043);
  or2  I080_257(w_080_257, w_028_005, w_004_097);
  and2 I080_269(w_080_269, w_023_073, w_070_192);
  and2 I080_279(w_080_279, w_035_114, w_073_020);
  not1 I080_284(w_080_284, w_056_610);
  nand2 I080_287(w_080_287, w_037_338, w_056_120);
  or2  I080_289(w_080_289, w_026_045, w_044_048);
  or2  I080_290(w_080_290, w_051_095, w_048_000);
  nand2 I080_295(w_080_295, w_049_200, w_046_201);
  nand2 I080_303(w_080_303, w_063_218, w_016_003);
  or2  I080_311(w_080_311, w_025_205, w_075_014);
  and2 I080_313(w_080_313, w_074_169, w_043_012);
  or2  I080_319(w_080_319, w_031_566, w_030_318);
  nand2 I080_336(w_080_336, w_066_402, w_010_682);
  or2  I080_360(w_080_360, w_003_070, w_074_124);
  not1 I080_362(w_080_362, w_032_583);
  nand2 I080_369(w_080_369, w_012_072, w_079_044);
  or2  I080_389(w_080_389, w_035_111, w_032_345);
  nand2 I080_394(w_080_394, w_026_613, w_045_177);
  or2  I080_397(w_080_397, w_074_000, w_043_013);
  and2 I080_399(w_080_399, w_072_178, w_002_458);
  or2  I080_403(w_080_403, w_043_019, w_018_035);
  or2  I080_407(w_080_407, w_058_383, w_045_157);
  or2  I080_417(w_080_417, w_066_119, w_015_204);
  not1 I080_430(w_080_430, w_074_111);
  and2 I080_433(w_080_433, w_029_036, w_004_301);
  or2  I080_440(w_080_440, w_013_012, w_057_006);
  not1 I080_464(w_080_464, w_062_003);
  and2 I080_472(w_080_472, w_078_039, w_044_465);
  nand2 I080_476(w_080_476, w_052_008, w_039_035);
  not1 I080_477(w_080_477, w_064_153);
  or2  I080_478(w_080_478, w_055_339, w_042_152);
  and2 I080_481(w_080_481, w_057_073, w_013_269);
  nand2 I081_000(w_081_000, w_037_218, w_055_088);
  not1 I081_001(w_081_001, w_051_148);
  nand2 I081_002(w_081_002, w_004_045, w_062_099);
  or2  I081_003(w_081_003, w_000_475, w_053_071);
  and2 I081_004(w_081_004, w_070_280, w_045_050);
  not1 I081_005(w_081_005, w_039_478);
  or2  I081_006(w_081_006, w_045_149, w_004_289);
  or2  I081_007(w_081_007, w_041_408, w_010_759);
  not1 I081_008(w_081_008, w_077_522);
  or2  I081_009(w_081_009, w_000_277, w_008_322);
  nand2 I081_010(w_081_010, w_008_031, w_015_135);
  not1 I081_011(w_081_011, w_020_416);
  nand2 I081_012(w_081_012, w_072_278, w_046_037);
  nand2 I081_013(w_081_013, w_011_062, w_072_289);
  nand2 I081_014(w_081_014, w_033_197, w_057_036);
  nand2 I081_015(w_081_015, w_069_110, w_062_000);
  nand2 I081_016(w_081_016, w_005_003, w_002_651);
  and2 I081_017(w_081_017, w_017_116, w_035_127);
  nand2 I081_018(w_081_018, w_042_072, w_045_294);
  or2  I081_019(w_081_019, w_032_594, w_070_459);
  nand2 I081_020(w_081_020, w_036_088, w_042_059);
  and2 I081_021(w_081_021, w_012_294, w_078_149);
  or2  I081_022(w_081_022, w_037_068, w_036_046);
  or2  I082_003(w_082_003, w_012_215, w_008_742);
  nand2 I082_019(w_082_019, w_029_098, w_020_140);
  and2 I082_020(w_082_020, w_055_047, w_065_086);
  or2  I082_026(w_082_026, w_011_357, w_051_312);
  or2  I082_027(w_082_027, w_027_116, w_030_231);
  and2 I082_040(w_082_040, w_016_006, w_081_014);
  not1 I082_041(w_082_041, w_047_038);
  and2 I082_044(w_082_044, w_004_238, w_034_072);
  not1 I082_049(w_082_049, w_039_121);
  nand2 I082_051(w_082_051, w_052_035, w_067_302);
  not1 I082_053(w_082_053, w_075_079);
  and2 I082_058(w_082_058, w_026_082, w_069_016);
  and2 I082_059(w_082_059, w_031_030, w_054_114);
  and2 I082_066(w_082_066, w_041_246, w_044_169);
  not1 I082_069(w_082_069, w_059_431);
  nand2 I082_070(w_082_070, w_039_175, w_076_432);
  and2 I082_073(w_082_073, w_075_076, w_017_057);
  and2 I082_079(w_082_079, w_031_444, w_060_009);
  and2 I082_082(w_082_082, w_022_124, w_030_167);
  not1 I082_090(w_082_090, w_034_037);
  and2 I082_092(w_082_092, w_005_022, w_070_019);
  not1 I082_104(w_082_104, w_045_038);
  nand2 I082_106(w_082_106, w_014_187, w_025_178);
  or2  I082_112(w_082_112, w_038_526, w_004_094);
  and2 I082_115(w_082_115, w_045_168, w_058_022);
  or2  I082_122(w_082_122, w_061_227, w_065_214);
  nand2 I082_123(w_082_123, w_062_088, w_028_117);
  nand2 I082_128(w_082_128, w_008_475, w_063_178);
  not1 I082_130(w_082_130, w_006_188);
  or2  I082_135(w_082_135, w_014_016, w_050_274);
  nand2 I082_139(w_082_139, w_058_597, w_057_058);
  or2  I082_140(w_082_140, w_029_101, w_034_003);
  or2  I082_141(w_082_141, w_040_373, w_030_367);
  not1 I082_142(w_082_142, w_081_000);
  nand2 I082_148(w_082_148, w_034_063, w_010_522);
  nand2 I082_150(w_082_150, w_002_055, w_076_421);
  and2 I082_154(w_082_154, w_033_462, w_031_124);
  and2 I082_160(w_082_160, w_059_479, w_060_030);
  or2  I082_162(w_082_162, w_027_104, w_053_009);
  not1 I082_166(w_082_166, w_013_301);
  not1 I082_167(w_082_167, w_075_018);
  nand2 I082_175(w_082_175, w_036_231, w_050_412);
  and2 I082_191(w_082_191, w_060_053, w_033_660);
  or2  I082_193(w_082_193, w_000_441, w_012_234);
  not1 I082_196(w_082_196, w_076_104);
  and2 I082_199(w_082_199, w_034_027, w_003_054);
  not1 I082_213(w_082_213, w_013_578);
  not1 I082_214(w_082_214, w_041_339);
  and2 I082_215(w_082_215, w_010_228, w_014_205);
  or2  I082_218(w_082_218, w_034_068, w_069_067);
  not1 I082_228(w_082_228, w_000_440);
  nand2 I082_235(w_082_235, w_009_096, w_065_107);
  nand2 I082_240(w_082_240, w_054_394, w_030_136);
  nand2 I082_244(w_082_244, w_021_251, w_018_026);
  nand2 I082_247(w_082_247, w_030_212, w_028_254);
  and2 I082_270(w_082_270, w_076_052, w_057_135);
  or2  I082_291(w_082_291, w_051_256, w_074_030);
  nand2 I082_299(w_082_299, w_037_231, w_069_022);
  or2  I082_303(w_082_303, w_030_020, w_009_523);
  nand2 I082_309(w_082_309, w_037_333, w_028_128);
  or2  I082_314(w_082_314, w_066_416, w_010_359);
  not1 I082_323(w_082_323, w_057_307);
  nand2 I082_336(w_082_336, w_068_346, w_013_078);
  and2 I082_338(w_082_338, w_081_019, w_012_009);
  not1 I082_383(w_082_383, w_002_048);
  or2  I082_389(w_082_389, w_059_533, w_011_253);
  nand2 I082_393(w_082_393, w_064_059, w_033_022);
  nand2 I082_409(w_082_409, w_061_256, w_010_522);
  and2 I082_423(w_082_423, w_065_407, w_014_271);
  and2 I082_425(w_082_425, w_027_140, w_041_088);
  or2  I082_431(w_082_431, w_080_085, w_011_333);
  not1 I082_455(w_082_455, w_070_480);
  not1 I082_463(w_082_463, w_045_191);
  nand2 I082_486(w_082_486, w_060_268, w_044_072);
  nand2 I082_487(w_082_487, w_015_183, w_058_536);
  and2 I082_502(w_082_502, w_078_070, w_050_611);
  not1 I082_505(w_082_505, w_081_019);
  or2  I082_511(w_082_511, w_002_329, w_079_016);
  or2  I082_526(w_082_526, w_010_258, w_012_003);
  nand2 I082_531(w_082_531, w_022_365, w_030_315);
  nand2 I082_538(w_082_538, w_056_332, w_022_271);
  and2 I082_540(w_082_540, w_057_060, w_001_012);
  or2  I082_541(w_082_541, w_038_053, w_070_089);
  nand2 I082_546(w_082_546, w_063_212, w_067_316);
  or2  I082_551(w_082_551, w_022_364, w_069_232);
  not1 I082_576(w_082_576, w_016_002);
  nand2 I082_577(w_082_577, w_073_042, w_078_053);
  nand2 I083_007(w_083_007, w_028_060, w_031_595);
  and2 I083_008(w_083_008, w_058_111, w_058_274);
  or2  I083_009(w_083_009, w_012_260, w_015_376);
  or2  I083_011(w_083_011, w_014_100, w_046_477);
  nand2 I083_013(w_083_013, w_063_059, w_059_552);
  and2 I083_017(w_083_017, w_081_003, w_050_161);
  nand2 I083_018(w_083_018, w_065_558, w_002_285);
  and2 I083_019(w_083_019, w_060_037, w_000_014);
  not1 I083_021(w_083_021, w_027_053);
  nand2 I083_022(w_083_022, w_068_224, w_017_073);
  nand2 I083_023(w_083_023, w_065_117, w_020_139);
  and2 I083_033(w_083_033, w_038_203, w_075_077);
  or2  I083_036(w_083_036, w_014_254, w_000_025);
  or2  I083_040(w_083_040, w_016_008, w_082_154);
  or2  I083_043(w_083_043, w_021_227, w_072_171);
  not1 I083_044(w_083_044, w_035_057);
  nand2 I083_046(w_083_046, w_077_026, w_012_273);
  and2 I083_052(w_083_052, w_063_469, w_003_011);
  nand2 I083_057(w_083_057, w_078_004, w_040_146);
  or2  I083_061(w_083_061, w_054_323, w_048_014);
  nand2 I083_066(w_083_066, w_081_022, w_016_008);
  not1 I083_067(w_083_067, w_056_317);
  or2  I083_068(w_083_068, w_050_602, w_025_290);
  and2 I083_071(w_083_071, w_070_253, w_062_140);
  or2  I083_073(w_083_073, w_001_014, w_070_325);
  or2  I083_085(w_083_085, w_067_021, w_029_090);
  nand2 I083_088(w_083_088, w_020_568, w_040_067);
  nand2 I083_093(w_083_093, w_033_181, w_080_182);
  nand2 I083_098(w_083_098, w_038_423, w_068_070);
  and2 I083_103(w_083_103, w_081_000, w_032_121);
  not1 I083_110(w_083_110, w_071_206);
  nand2 I083_113(w_083_113, w_011_566, w_055_255);
  not1 I083_115(w_083_115, w_020_598);
  nand2 I083_116(w_083_116, w_005_042, w_009_181);
  and2 I083_118(w_083_118, w_000_725, w_045_375);
  or2  I083_123(w_083_123, w_060_354, w_074_337);
  nand2 I083_127(w_083_127, w_078_083, w_046_609);
  not1 I083_129(w_083_129, w_044_348);
  or2  I083_135(w_083_135, w_030_007, w_014_288);
  nand2 I083_138(w_083_138, w_080_476, w_010_533);
  not1 I083_140(w_083_140, w_017_337);
  or2  I083_144(w_083_144, w_021_105, w_001_028);
  or2  I083_147(w_083_147, w_066_627, w_052_042);
  not1 I083_149(w_083_149, w_056_046);
  and2 I083_151(w_083_151, w_049_190, w_020_024);
  not1 I083_153(w_083_153, w_019_009);
  and2 I083_154(w_083_154, w_029_081, w_034_009);
  and2 I083_155(w_083_155, w_036_393, w_026_382);
  not1 I083_156(w_083_156, w_052_026);
  not1 I083_158(w_083_158, w_067_104);
  or2  I083_163(w_083_163, w_020_169, w_009_132);
  and2 I083_165(w_083_165, w_060_058, w_060_126);
  not1 I083_166(w_083_166, w_034_054);
  not1 I083_168(w_083_168, w_039_263);
  nand2 I083_169(w_083_169, w_054_534, w_030_354);
  nand2 I083_170(w_083_170, w_006_062, w_054_410);
  and2 I083_175(w_083_175, w_040_102, w_070_232);
  not1 I083_181(w_083_181, w_060_323);
  not1 I083_182(w_083_182, w_017_380);
  or2  I083_183(w_083_183, w_070_191, w_003_057);
  or2  I083_187(w_083_187, w_073_499, w_020_010);
  or2  I083_189(w_083_189, w_042_111, w_030_035);
  or2  I083_190(w_083_190, w_008_205, w_075_014);
  nand2 I083_191(w_083_191, w_025_157, w_062_484);
  not1 I083_192(w_083_192, w_006_071);
  not1 I083_193(w_083_193, w_020_084);
  or2  I084_000(w_084_000, w_076_240, w_017_540);
  not1 I084_001(w_084_001, w_016_008);
  not1 I084_002(w_084_002, w_039_625);
  nand2 I084_003(w_084_003, w_073_071, w_043_005);
  or2  I084_004(w_084_004, w_006_054, w_052_008);
  not1 I084_005(w_084_005, w_020_001);
  nand2 I084_006(w_084_006, w_045_041, w_051_351);
  and2 I084_007(w_084_007, w_008_364, w_065_084);
  or2  I084_008(w_084_008, w_021_148, w_049_020);
  and2 I084_009(w_084_009, w_004_269, w_071_155);
  or2  I084_010(w_084_010, w_070_142, w_006_224);
  or2  I084_011(w_084_011, w_058_442, w_075_054);
  and2 I084_012(w_084_012, w_050_236, w_073_101);
  nand2 I084_013(w_084_013, w_062_745, w_031_471);
  or2  I084_014(w_084_014, w_064_080, w_011_026);
  and2 I084_015(w_084_015, w_076_098, w_037_051);
  and2 I084_016(w_084_016, w_054_230, w_003_056);
  not1 I084_017(w_084_017, w_037_295);
  or2  I084_018(w_084_018, w_028_058, w_041_399);
  or2  I084_020(w_084_020, w_048_018, w_060_336);
  nand2 I084_021(w_084_021, w_080_019, w_063_166);
  and2 I084_023(w_084_023, w_039_068, w_079_020);
  nand2 I084_024(w_084_024, w_032_123, w_048_005);
  or2  I084_025(w_084_025, w_005_204, w_043_019);
  and2 I084_026(w_084_026, w_033_016, w_002_405);
  and2 I084_028(w_084_028, w_014_243, w_040_415);
  not1 I084_029(w_084_029, w_076_295);
  nand2 I084_030(w_084_030, w_027_161, w_014_279);
  nand2 I084_032(w_084_032, w_023_137, w_078_078);
  or2  I084_033(w_084_033, w_027_083, w_016_000);
  not1 I084_034(w_084_034, w_026_311);
  nand2 I084_036(w_084_036, w_043_021, w_007_226);
  and2 I084_037(w_084_037, w_034_045, w_038_002);
  nand2 I084_038(w_084_038, w_016_006, w_046_171);
  and2 I084_039(w_084_039, w_040_054, w_058_376);
  and2 I084_040(w_084_040, w_074_296, w_026_668);
  not1 I084_042(w_084_042, w_042_298);
  nand2 I084_043(w_084_043, w_005_076, w_068_361);
  or2  I084_044(w_084_044, w_022_316, w_068_307);
  or2  I084_045(w_084_045, w_030_051, w_002_022);
  and2 I084_046(w_084_046, w_060_310, w_013_194);
  nand2 I084_047(w_084_047, w_039_646, w_071_055);
  or2  I084_048(w_084_048, w_014_180, w_047_129);
  not1 I085_001(w_085_001, w_071_031);
  or2  I085_011(w_085_011, w_034_006, w_071_250);
  nand2 I085_015(w_085_015, w_042_339, w_061_314);
  and2 I085_016(w_085_016, w_010_570, w_065_606);
  and2 I085_017(w_085_017, w_004_177, w_061_365);
  nand2 I085_022(w_085_022, w_079_043, w_003_031);
  or2  I085_024(w_085_024, w_036_400, w_056_500);
  or2  I085_026(w_085_026, w_079_003, w_084_006);
  and2 I085_027(w_085_027, w_043_036, w_051_136);
  nand2 I085_028(w_085_028, w_054_203, w_035_117);
  or2  I085_029(w_085_029, w_041_380, w_044_306);
  not1 I085_030(w_085_030, w_000_094);
  and2 I085_034(w_085_034, w_072_135, w_060_036);
  or2  I085_037(w_085_037, w_080_186, w_070_478);
  or2  I085_038(w_085_038, w_005_002, w_044_670);
  or2  I085_040(w_085_040, w_083_181, w_032_540);
  nand2 I085_042(w_085_042, w_065_311, w_084_004);
  and2 I085_045(w_085_045, w_068_012, w_079_059);
  and2 I085_048(w_085_048, w_049_172, w_034_062);
  or2  I085_051(w_085_051, w_054_133, w_030_340);
  nand2 I085_056(w_085_056, w_016_001, w_071_277);
  not1 I085_059(w_085_059, w_024_032);
  or2  I085_068(w_085_068, w_030_048, w_025_192);
  not1 I085_070(w_085_070, w_031_392);
  or2  I085_074(w_085_074, w_030_325, w_061_205);
  and2 I085_080(w_085_080, w_083_022, w_050_440);
  and2 I085_084(w_085_084, w_072_215, w_021_261);
  and2 I085_085(w_085_085, w_037_177, w_054_003);
  not1 I085_087(w_085_087, w_024_300);
  or2  I085_088(w_085_088, w_049_074, w_000_138);
  or2  I085_092(w_085_092, w_010_089, w_055_039);
  nand2 I085_096(w_085_096, w_036_368, w_021_266);
  nand2 I085_116(w_085_116, w_001_032, w_069_191);
  or2  I085_125(w_085_125, w_065_066, w_040_441);
  nand2 I085_129(w_085_129, w_049_130, w_027_093);
  or2  I085_139(w_085_139, w_023_197, w_009_228);
  or2  I085_141(w_085_141, w_030_220, w_043_011);
  nand2 I085_146(w_085_146, w_077_032, w_062_138);
  or2  I085_150(w_085_150, w_010_102, w_026_502);
  or2  I085_152(w_085_152, w_028_142, w_048_018);
  not1 I085_158(w_085_158, w_084_005);
  not1 I085_161(w_085_161, w_053_024);
  not1 I085_162(w_085_162, w_023_053);
  nand2 I085_164(w_085_164, w_058_182, w_011_024);
  or2  I085_167(w_085_167, w_007_088, w_072_120);
  or2  I085_173(w_085_173, w_072_184, w_075_001);
  or2  I085_176(w_085_176, w_072_060, w_002_206);
  or2  I085_190(w_085_190, w_037_251, w_057_029);
  or2  I085_199(w_085_199, w_018_017, w_060_284);
  not1 I085_201(w_085_201, w_064_328);
  or2  I085_202(w_085_202, w_002_072, w_008_193);
  nand2 I085_203(w_085_203, w_016_006, w_065_015);
  and2 I085_205(w_085_205, w_080_079, w_013_201);
  nand2 I085_219(w_085_219, w_081_016, w_045_067);
  and2 I085_220(w_085_220, w_020_105, w_001_020);
  nand2 I085_226(w_085_226, w_010_497, w_006_100);
  and2 I085_230(w_085_230, w_022_305, w_041_627);
  or2  I085_244(w_085_244, w_011_260, w_045_014);
  not1 I085_246(w_085_246, w_017_496);
  nand2 I085_255(w_085_255, w_045_204, w_027_178);
  and2 I085_257(w_085_257, w_038_120, w_043_026);
  not1 I085_265(w_085_265, w_035_031);
  nand2 I085_272(w_085_272, w_000_514, w_014_072);
  or2  I085_277(w_085_277, w_009_160, w_050_205);
  and2 I085_294(w_085_294, w_030_229, w_014_219);
  or2  I085_295(w_085_295, w_048_003, w_016_000);
  nand2 I085_298(w_085_298, w_049_324, w_063_326);
  and2 I085_299(w_085_299, w_044_723, w_076_130);
  and2 I085_305(w_085_305, w_058_550, w_064_029);
  or2  I085_306(w_085_306, w_055_257, w_015_047);
  or2  I085_309(w_085_309, w_043_029, w_081_018);
  nand2 I085_320(w_085_320, w_039_104, w_015_382);
  or2  I085_327(w_085_327, w_065_253, w_066_084);
  and2 I085_329(w_085_329, w_003_069, w_010_576);
  nand2 I085_338(w_085_338, w_013_093, w_030_274);
  not1 I085_340(w_085_340, w_074_250);
  nand2 I085_349(w_085_349, w_040_617, w_048_007);
  nand2 I085_350(w_085_350, w_024_391, w_073_026);
  not1 I085_353(w_085_353, w_036_267);
  and2 I085_354(w_085_356, w_085_355, w_003_080);
  nand2 I085_355(w_085_357, w_085_356, w_068_200);
  not1 I085_356(w_085_358, w_085_357);
  nand2 I085_357(w_085_359, w_012_176, w_085_358);
  nand2 I085_358(w_085_360, w_085_359, w_006_008);
  or2  I085_359(w_085_361, w_085_360, w_005_292);
  and2 I085_360(w_085_362, w_001_001, w_085_361);
  not1 I085_361(w_085_355, w_085_362);
  nand2 I086_003(w_086_003, w_076_145, w_055_045);
  and2 I086_007(w_086_007, w_026_480, w_047_246);
  not1 I086_009(w_086_009, w_020_149);
  and2 I086_010(w_086_010, w_066_224, w_078_043);
  or2  I086_022(w_086_022, w_028_190, w_003_034);
  not1 I086_024(w_086_024, w_061_084);
  nand2 I086_028(w_086_028, w_018_020, w_021_006);
  nand2 I086_029(w_086_029, w_041_197, w_025_135);
  and2 I086_032(w_086_032, w_056_665, w_060_259);
  and2 I086_033(w_086_033, w_036_211, w_054_081);
  not1 I086_034(w_086_034, w_080_255);
  and2 I086_043(w_086_043, w_006_096, w_049_164);
  nand2 I086_046(w_086_046, w_006_095, w_021_223);
  not1 I086_049(w_086_049, w_050_110);
  not1 I086_051(w_086_051, w_027_056);
  or2  I086_055(w_086_055, w_013_150, w_070_404);
  nand2 I086_059(w_086_059, w_075_145, w_037_097);
  and2 I086_062(w_086_062, w_015_431, w_071_099);
  nand2 I086_064(w_086_064, w_000_405, w_032_596);
  or2  I086_065(w_086_065, w_031_160, w_026_354);
  nand2 I086_067(w_086_067, w_024_178, w_034_022);
  not1 I086_073(w_086_073, w_033_727);
  nand2 I086_078(w_086_078, w_066_343, w_011_319);
  not1 I086_081(w_086_081, w_007_263);
  not1 I086_083(w_086_083, w_044_454);
  nand2 I086_089(w_086_089, w_000_144, w_045_043);
  and2 I086_091(w_086_091, w_014_015, w_036_245);
  and2 I086_093(w_086_093, w_081_016, w_049_249);
  and2 I086_095(w_086_095, w_082_336, w_000_291);
  and2 I086_097(w_086_097, w_039_221, w_026_009);
  not1 I086_098(w_086_098, w_037_207);
  and2 I086_101(w_086_101, w_079_036, w_054_085);
  and2 I086_119(w_086_119, w_035_115, w_036_294);
  or2  I086_122(w_086_122, w_047_050, w_070_010);
  and2 I086_124(w_086_124, w_016_008, w_039_425);
  or2  I086_133(w_086_133, w_032_445, w_053_119);
  nand2 I086_134(w_086_134, w_064_289, w_032_297);
  not1 I086_144(w_086_144, w_065_658);
  not1 I086_151(w_086_151, w_008_206);
  and2 I086_158(w_086_158, w_085_320, w_006_000);
  not1 I086_160(w_086_160, w_080_185);
  nand2 I086_161(w_086_161, w_019_001, w_057_052);
  or2  I086_164(w_086_164, w_053_071, w_076_418);
  nand2 I086_173(w_086_173, w_034_068, w_011_341);
  and2 I086_175(w_086_175, w_015_288, w_016_005);
  nand2 I086_179(w_086_179, w_033_148, w_005_023);
  not1 I086_181(w_086_181, w_010_122);
  not1 I086_182(w_086_182, w_026_217);
  nand2 I086_185(w_086_185, w_014_254, w_072_201);
  and2 I086_187(w_086_187, w_012_008, w_068_334);
  not1 I086_189(w_086_189, w_028_079);
  and2 I086_190(w_086_190, w_027_102, w_080_011);
  and2 I086_192(w_086_192, w_047_413, w_062_546);
  or2  I086_195(w_086_195, w_066_512, w_013_230);
  and2 I086_197(w_086_197, w_006_155, w_000_308);
  or2  I086_201(w_086_201, w_049_204, w_068_153);
  or2  I086_208(w_086_208, w_002_359, w_081_007);
  or2  I086_232(w_086_232, w_053_010, w_048_007);
  nand2 I086_236(w_086_236, w_077_242, w_027_139);
  and2 I086_237(w_086_237, w_048_003, w_022_188);
  or2  I086_253(w_086_253, w_047_465, w_067_206);
  or2  I086_264(w_086_264, w_011_162, w_001_003);
  nand2 I086_265(w_086_265, w_047_209, w_067_119);
  or2  I086_270(w_086_270, w_051_140, w_078_101);
  nand2 I086_275(w_086_275, w_012_297, w_041_346);
  not1 I086_277(w_086_277, w_073_150);
  not1 I086_307(w_086_307, w_078_016);
  nand2 I086_312(w_086_312, w_007_439, w_048_014);
  and2 I086_313(w_086_313, w_065_228, w_068_124);
  and2 I086_320(w_086_320, w_085_203, w_082_423);
  or2  I086_321(w_086_321, w_068_113, w_081_011);
  or2  I086_332(w_086_332, w_084_045, w_052_001);
  not1 I086_336(w_086_336, w_079_028);
  or2  I086_343(w_086_343, w_050_007, w_010_709);
  and2 I086_344(w_085_364, w_030_041, w_085_355);
  nand2 I087_013(w_087_013, w_072_167, w_043_022);
  or2  I087_015(w_087_015, w_079_053, w_035_108);
  not1 I087_018(w_087_018, w_052_038);
  not1 I087_025(w_087_025, w_026_457);
  nand2 I087_028(w_087_028, w_044_690, w_054_149);
  or2  I087_037(w_087_037, w_064_009, w_005_102);
  not1 I087_040(w_087_040, w_017_305);
  and2 I087_043(w_087_043, w_004_228, w_023_027);
  nand2 I087_048(w_087_048, w_082_140, w_037_208);
  nand2 I087_051(w_087_051, w_015_534, w_026_513);
  not1 I087_054(w_087_054, w_082_538);
  or2  I087_058(w_087_058, w_006_116, w_021_200);
  not1 I087_065(w_087_065, w_051_286);
  or2  I087_069(w_087_069, w_022_000, w_065_063);
  and2 I087_071(w_087_071, w_061_241, w_075_105);
  and2 I087_086(w_087_086, w_081_018, w_032_194);
  or2  I087_088(w_087_088, w_025_094, w_063_297);
  not1 I087_098(w_087_098, w_020_266);
  and2 I087_100(w_087_100, w_060_148, w_063_456);
  or2  I087_102(w_087_102, w_009_540, w_041_489);
  or2  I087_106(w_087_106, w_035_018, w_012_191);
  not1 I087_117(w_087_117, w_000_176);
  and2 I087_118(w_087_118, w_068_174, w_001_033);
  and2 I087_120(w_087_120, w_027_105, w_024_119);
  not1 I087_125(w_087_125, w_059_150);
  or2  I087_127(w_087_127, w_032_149, w_011_071);
  nand2 I087_134(w_087_134, w_055_324, w_060_190);
  not1 I087_137(w_087_137, w_009_359);
  or2  I087_149(w_087_149, w_037_267, w_021_093);
  or2  I087_154(w_087_154, w_010_131, w_075_083);
  and2 I087_156(w_087_156, w_007_296, w_068_098);
  and2 I087_160(w_087_160, w_011_132, w_039_536);
  or2  I087_162(w_087_162, w_076_476, w_038_386);
  or2  I087_165(w_087_165, w_083_187, w_061_443);
  and2 I087_168(w_087_168, w_032_464, w_008_181);
  not1 I087_182(w_087_182, w_061_300);
  and2 I087_186(w_087_186, w_054_058, w_073_037);
  or2  I087_189(w_087_189, w_045_013, w_079_057);
  and2 I087_190(w_087_190, w_030_172, w_073_016);
  nand2 I087_195(w_087_195, w_056_620, w_075_140);
  and2 I087_204(w_087_204, w_051_074, w_017_128);
  not1 I087_205(w_087_205, w_049_231);
  or2  I087_207(w_087_207, w_084_034, w_021_009);
  or2  I087_215(w_087_215, w_045_039, w_075_155);
  and2 I087_216(w_087_216, w_041_524, w_058_699);
  and2 I087_219(w_087_219, w_045_151, w_066_089);
  or2  I087_227(w_087_227, w_031_570, w_028_064);
  not1 I087_228(w_087_228, w_085_364);
  or2  I087_230(w_087_230, w_035_126, w_078_188);
  nand2 I087_235(w_087_235, w_036_053, w_001_005);
  nand2 I087_243(w_087_243, w_058_088, w_081_018);
  not1 I087_247(w_087_247, w_052_025);
  not1 I087_249(w_087_249, w_064_327);
  or2  I087_253(w_087_253, w_038_472, w_039_650);
  not1 I087_255(w_087_255, w_031_218);
  nand2 I087_258(w_087_258, w_004_212, w_075_010);
  and2 I087_273(w_087_273, w_083_135, w_047_221);
  or2  I087_286(w_087_286, w_062_785, w_015_069);
  or2  I087_292(w_087_292, w_084_014, w_046_272);
  and2 I087_293(w_087_293, w_065_557, w_083_013);
  and2 I087_298(w_087_298, w_033_162, w_017_555);
  not1 I087_310(w_087_310, w_069_048);
  or2  I087_311(w_087_311, w_074_344, w_048_008);
  not1 I087_323(w_087_323, w_018_021);
  not1 I087_326(w_087_326, w_030_315);
  and2 I087_333(w_087_333, w_068_062, w_020_378);
  and2 I087_335(w_087_335, w_038_337, w_002_443);
  nand2 I087_343(w_087_343, w_044_219, w_068_322);
  and2 I087_357(w_087_357, w_085_129, w_033_191);
  nand2 I087_358(w_087_358, w_018_036, w_019_004);
  and2 I087_366(w_087_366, w_059_730, w_046_341);
  not1 I087_372(w_087_372, w_074_111);
  and2 I087_379(w_087_379, w_007_130, w_004_453);
  not1 I087_381(w_087_381, w_022_347);
  and2 I087_387(w_087_387, w_023_023, w_024_056);
  nand2 I087_407(w_087_407, w_062_220, w_021_150);
  or2  I087_408(w_087_408, w_025_102, w_037_133);
  or2  I087_425(w_087_425, w_064_027, w_005_300);
  or2  I087_431(w_087_431, w_035_025, w_020_078);
  or2  I088_002(w_088_002, w_006_011, w_069_068);
  not1 I088_003(w_088_003, w_030_106);
  or2  I088_005(w_088_005, w_059_084, w_070_386);
  and2 I088_011(w_088_011, w_038_521, w_013_106);
  or2  I088_012(w_088_012, w_084_040, w_055_154);
  and2 I088_013(w_088_013, w_010_042, w_066_035);
  or2  I088_015(w_088_015, w_037_323, w_049_342);
  or2  I088_016(w_088_016, w_030_101, w_073_735);
  nand2 I088_018(w_088_018, w_007_221, w_049_107);
  and2 I088_019(w_088_019, w_080_159, w_024_339);
  not1 I088_020(w_088_020, w_066_559);
  or2  I088_021(w_088_021, w_052_031, w_066_385);
  nand2 I088_022(w_088_022, w_015_256, w_028_029);
  not1 I088_023(w_088_023, w_059_131);
  nand2 I088_024(w_088_024, w_026_381, w_045_286);
  or2  I088_025(w_088_025, w_053_151, w_034_028);
  nand2 I088_028(w_088_028, w_025_005, w_085_088);
  not1 I088_029(w_088_029, w_077_251);
  or2  I088_031(w_088_031, w_077_440, w_055_035);
  not1 I088_032(w_088_032, w_063_388);
  nand2 I088_033(w_088_033, w_038_070, w_035_001);
  not1 I088_036(w_088_036, w_076_347);
  and2 I088_041(w_088_041, w_014_145, w_053_023);
  or2  I088_043(w_088_043, w_036_157, w_062_313);
  and2 I088_044(w_088_044, w_049_140, w_077_372);
  not1 I088_045(w_088_045, w_056_229);
  and2 I088_046(w_088_046, w_062_653, w_052_008);
  nand2 I088_048(w_088_048, w_023_054, w_018_025);
  nand2 I088_050(w_088_050, w_007_014, w_050_280);
  not1 I088_051(w_088_051, w_011_421);
  nand2 I088_052(w_088_052, w_015_423, w_019_003);
  and2 I088_053(w_088_053, w_081_020, w_024_145);
  and2 I088_055(w_088_055, w_025_179, w_078_056);
  nand2 I088_060(w_088_060, w_050_130, w_079_031);
  nand2 I088_061(w_088_061, w_080_440, w_059_201);
  not1 I088_062(w_088_062, w_050_257);
  not1 I088_063(w_088_063, w_011_508);
  not1 I088_065(w_088_065, w_056_491);
  or2  I088_066(w_088_066, w_000_344, w_040_286);
  not1 I088_067(w_088_067, w_017_349);
  or2  I088_069(w_088_069, w_068_357, w_022_240);
  nand2 I088_070(w_088_070, w_032_022, w_002_564);
  not1 I088_076(w_088_076, w_011_172);
  and2 I088_079(w_088_079, w_009_294, w_046_314);
  or2  I088_080(w_088_080, w_024_193, w_046_092);
  not1 I088_089(w_088_089, w_050_334);
  not1 I088_090(w_088_090, w_004_098);
  nand2 I088_093(w_088_093, w_024_039, w_033_086);
  nand2 I088_094(w_088_094, w_007_045, w_085_017);
  not1 I088_102(w_088_102, w_060_198);
  and2 I088_106(w_088_106, w_001_028, w_049_174);
  not1 I088_117(w_088_117, w_058_658);
  not1 I088_119(w_088_119, w_031_234);
  not1 I088_121(w_088_121, w_068_268);
  not1 I088_125(w_088_125, w_085_190);
  or2  I088_126(w_088_126, w_069_055, w_005_159);
  not1 I088_129(w_088_129, w_018_035);
  or2  I088_130(w_088_130, w_004_135, w_040_174);
  not1 I088_131(w_088_131, w_028_523);
  or2  I088_132(w_088_132, w_002_681, w_019_008);
  and2 I088_135(w_088_135, w_069_009, w_016_004);
  not1 I088_136(w_088_136, w_048_008);
  or2  I088_143(w_088_143, w_000_432, w_002_516);
  not1 I089_006(w_089_006, w_006_078);
  or2  I089_009(w_089_009, w_059_029, w_056_622);
  nand2 I089_012(w_089_012, w_083_140, w_047_049);
  not1 I089_013(w_089_013, w_086_083);
  and2 I089_017(w_089_017, w_020_010, w_030_101);
  nand2 I089_025(w_089_025, w_003_027, w_050_475);
  nand2 I089_026(w_089_026, w_044_036, w_082_044);
  and2 I089_028(w_089_028, w_078_588, w_079_004);
  not1 I089_033(w_089_033, w_044_686);
  nand2 I089_042(w_089_042, w_048_016, w_071_031);
  nand2 I089_045(w_089_045, w_008_698, w_032_053);
  and2 I089_051(w_089_051, w_007_289, w_080_394);
  and2 I089_053(w_089_053, w_017_298, w_062_162);
  or2  I089_055(w_089_055, w_056_412, w_065_333);
  and2 I089_057(w_089_057, w_003_035, w_011_089);
  and2 I089_060(w_089_060, w_077_313, w_014_292);
  not1 I089_061(w_089_061, w_008_577);
  nand2 I089_068(w_089_068, w_061_088, w_079_012);
  nand2 I089_070(w_089_070, w_005_157, w_001_026);
  not1 I089_071(w_089_071, w_022_381);
  or2  I089_072(w_089_072, w_060_326, w_000_225);
  or2  I089_075(w_089_075, w_029_075, w_040_395);
  or2  I089_078(w_089_078, w_003_031, w_055_034);
  or2  I089_085(w_089_085, w_021_175, w_064_103);
  nand2 I089_086(w_089_086, w_051_200, w_022_155);
  not1 I089_089(w_089_089, w_026_216);
  nand2 I089_094(w_089_094, w_018_027, w_029_058);
  and2 I089_096(w_089_096, w_018_022, w_035_025);
  or2  I089_098(w_089_098, w_017_502, w_025_012);
  and2 I089_100(w_089_100, w_025_135, w_004_197);
  or2  I089_106(w_089_106, w_070_390, w_052_001);
  not1 I089_107(w_089_107, w_079_045);
  not1 I089_111(w_089_111, w_084_015);
  and2 I089_118(w_089_118, w_080_231, w_056_184);
  and2 I089_126(w_089_126, w_024_092, w_051_011);
  or2  I089_128(w_089_128, w_062_435, w_004_411);
  or2  I089_129(w_089_129, w_004_134, w_082_122);
  and2 I089_132(w_089_132, w_075_001, w_076_458);
  not1 I089_134(w_089_134, w_033_392);
  or2  I089_135(w_089_135, w_060_355, w_081_004);
  or2  I089_136(w_089_136, w_074_218, w_032_399);
  nand2 I089_138(w_089_138, w_024_079, w_033_224);
  not1 I089_140(w_089_140, w_086_009);
  or2  I089_142(w_089_142, w_042_199, w_072_103);
  not1 I089_144(w_089_144, w_057_235);
  not1 I089_149(w_089_149, w_078_428);
  nand2 I089_150(w_089_150, w_027_072, w_017_026);
  and2 I089_151(w_089_151, w_008_261, w_066_327);
  nand2 I089_155(w_089_155, w_058_050, w_037_024);
  or2  I089_156(w_089_156, w_026_348, w_012_045);
  or2  I089_160(w_089_160, w_067_297, w_056_020);
  not1 I089_164(w_089_164, w_044_500);
  or2  I089_166(w_089_166, w_069_105, w_027_016);
  nand2 I089_167(w_089_167, w_005_071, w_053_111);
  not1 I089_178(w_089_178, w_048_001);
  nand2 I089_185(w_089_185, w_014_274, w_074_144);
  not1 I089_190(w_089_190, w_006_034);
  or2  I089_191(w_089_191, w_076_015, w_079_017);
  not1 I089_197(w_089_197, w_020_100);
  not1 I089_198(w_089_198, w_070_473);
  nand2 I089_199(w_089_199, w_034_072, w_088_021);
  nand2 I089_206(w_089_206, w_054_033, w_073_085);
  and2 I089_210(w_089_210, w_069_168, w_048_004);
  nand2 I089_211(w_089_211, w_007_168, w_017_479);
  not1 I089_213(w_089_213, w_063_025);
  or2  I089_215(w_089_215, w_049_120, w_013_118);
  not1 I089_217(w_089_217, w_087_431);
  not1 I089_219(w_089_219, w_034_075);
  not1 I089_221(w_089_221, w_003_074);
  or2  I089_230(w_089_230, w_083_115, w_059_500);
  not1 I089_232(w_089_232, w_017_017);
  nand2 I089_258(w_089_258, w_036_272, w_001_016);
  and2 I089_259(w_089_259, w_009_570, w_068_298);
  nand2 I089_266(w_089_266, w_004_187, w_000_134);
  and2 I089_269(w_089_269, w_013_573, w_026_564);
  not1 I089_282(w_089_282, w_023_172);
  or2  I089_289(w_089_289, w_059_698, w_077_152);
  nand2 I089_291(w_089_291, w_070_499, w_016_006);
  and2 I089_300(w_089_300, w_086_182, w_053_119);
  nand2 I090_001(w_090_001, w_009_421, w_070_008);
  nand2 I090_011(w_090_011, w_008_725, w_063_003);
  nand2 I090_016(w_090_016, w_035_057, w_064_020);
  and2 I090_035(w_090_035, w_017_536, w_045_264);
  or2  I090_036(w_090_036, w_070_190, w_087_018);
  not1 I090_042(w_090_042, w_034_015);
  or2  I090_047(w_090_047, w_045_016, w_005_117);
  and2 I090_048(w_090_048, w_039_085, w_051_291);
  nand2 I090_052(w_090_052, w_036_256, w_017_495);
  or2  I090_061(w_090_061, w_029_089, w_053_066);
  or2  I090_063(w_090_063, w_075_050, w_056_487);
  not1 I090_066(w_090_066, w_059_159);
  not1 I090_067(w_090_067, w_084_005);
  nand2 I090_068(w_090_068, w_075_097, w_081_019);
  nand2 I090_072(w_090_072, w_034_037, w_051_084);
  not1 I090_080(w_090_080, w_034_005);
  or2  I090_086(w_090_086, w_018_035, w_074_111);
  nand2 I090_088(w_090_088, w_000_286, w_063_036);
  nand2 I090_117(w_090_117, w_055_345, w_048_013);
  or2  I090_122(w_090_122, w_045_044, w_036_221);
  nand2 I090_126(w_090_126, w_014_205, w_069_146);
  and2 I090_131(w_090_131, w_028_110, w_059_553);
  or2  I090_151(w_090_151, w_065_218, w_080_397);
  nand2 I090_168(w_090_168, w_067_382, w_029_066);
  nand2 I090_171(w_090_171, w_021_128, w_065_181);
  or2  I090_191(w_090_191, w_049_312, w_002_532);
  and2 I090_195(w_090_195, w_061_050, w_081_006);
  and2 I090_203(w_090_203, w_043_003, w_062_017);
  or2  I090_206(w_090_206, w_060_277, w_054_035);
  nand2 I090_218(w_090_218, w_088_045, w_079_055);
  not1 I090_221(w_090_221, w_030_235);
  not1 I090_222(w_090_222, w_030_269);
  or2  I090_223(w_090_223, w_018_024, w_019_003);
  nand2 I090_224(w_090_224, w_006_070, w_043_003);
  nand2 I090_232(w_090_232, w_010_183, w_074_175);
  and2 I090_242(w_090_242, w_035_040, w_058_332);
  nand2 I090_266(w_090_266, w_010_739, w_040_501);
  not1 I090_272(w_090_272, w_030_174);
  not1 I090_275(w_090_275, w_018_022);
  not1 I090_295(w_090_295, w_062_355);
  and2 I090_306(w_090_306, w_070_327, w_035_016);
  and2 I090_310(w_090_310, w_053_000, w_074_321);
  and2 I090_358(w_090_358, w_020_319, w_060_313);
  nand2 I090_362(w_090_362, w_037_152, w_061_057);
  not1 I090_370(w_090_370, w_060_071);
  and2 I090_380(w_090_380, w_063_233, w_005_055);
  or2  I090_384(w_090_384, w_028_198, w_018_023);
  nand2 I090_392(w_090_392, w_036_170, w_083_103);
  and2 I090_405(w_090_405, w_020_114, w_054_365);
  or2  I090_415(w_090_415, w_084_002, w_032_197);
  nand2 I090_420(w_090_420, w_037_235, w_080_225);
  or2  I090_442(w_090_442, w_059_147, w_022_343);
  and2 I090_451(w_090_451, w_027_161, w_025_201);
  and2 I090_464(w_090_464, w_086_179, w_034_017);
  not1 I090_469(w_090_469, w_004_149);
  not1 I090_472(w_090_472, w_067_347);
  nand2 I090_478(w_090_478, w_079_035, w_053_143);
  or2  I090_487(w_090_487, w_059_512, w_028_254);
  and2 I090_489(w_090_489, w_064_327, w_081_012);
  or2  I090_505(w_090_505, w_073_041, w_050_062);
  not1 I090_510(w_090_510, w_029_011);
  and2 I090_523(w_090_523, w_040_430, w_017_133);
  not1 I090_528(w_090_528, w_064_020);
  not1 I090_531(w_090_531, w_047_210);
  and2 I090_532(w_090_532, w_056_030, w_069_053);
  not1 I090_535(w_090_535, w_020_024);
  nand2 I090_536(w_090_536, w_075_144, w_076_099);
  and2 I090_542(w_090_542, w_009_354, w_009_097);
  not1 I090_543(w_090_543, w_085_164);
  not1 I090_564(w_090_564, w_027_155);
  not1 I091_000(w_091_000, w_035_069);
  and2 I091_008(w_091_008, w_056_017, w_061_012);
  and2 I091_012(w_091_012, w_042_258, w_089_033);
  and2 I091_014(w_091_014, w_089_282, w_059_348);
  or2  I091_020(w_091_020, w_001_014, w_066_516);
  and2 I091_024(w_091_024, w_048_014, w_070_104);
  nand2 I091_028(w_091_028, w_042_217, w_046_478);
  or2  I091_030(w_091_030, w_046_580, w_066_099);
  or2  I091_032(w_091_032, w_062_342, w_033_689);
  nand2 I091_033(w_091_033, w_011_325, w_076_296);
  not1 I091_034(w_091_034, w_032_102);
  and2 I091_036(w_091_036, w_017_042, w_019_014);
  not1 I091_037(w_091_037, w_085_265);
  and2 I091_039(w_091_039, w_078_170, w_088_053);
  or2  I091_040(w_091_040, w_063_019, w_034_006);
  not1 I091_041(w_091_041, w_067_062);
  not1 I091_042(w_091_042, w_018_032);
  or2  I091_043(w_091_043, w_007_089, w_019_011);
  nand2 I091_044(w_091_044, w_046_561, w_022_038);
  nand2 I091_046(w_091_046, w_013_471, w_073_499);
  not1 I091_056(w_091_056, w_024_347);
  or2  I091_059(w_091_059, w_047_404, w_033_278);
  nand2 I091_063(w_091_063, w_084_030, w_001_008);
  and2 I091_067(w_091_067, w_019_009, w_075_009);
  or2  I091_073(w_091_073, w_063_238, w_050_405);
  not1 I091_074(w_091_074, w_030_257);
  and2 I091_075(w_091_075, w_063_545, w_073_052);
  nand2 I091_077(w_091_077, w_079_017, w_062_696);
  and2 I091_078(w_091_078, w_024_070, w_035_126);
  and2 I091_080(w_091_080, w_020_479, w_018_025);
  or2  I091_081(w_091_081, w_042_222, w_010_050);
  not1 I091_085(w_091_085, w_051_231);
  or2  I091_088(w_091_088, w_007_271, w_022_201);
  nand2 I091_091(w_091_091, w_008_463, w_054_049);
  and2 I091_094(w_091_094, w_056_200, w_022_077);
  nand2 I091_095(w_091_095, w_008_278, w_080_417);
  not1 I091_105(w_091_105, w_027_134);
  nand2 I091_109(w_091_109, w_089_053, w_060_017);
  nand2 I091_111(w_091_111, w_089_210, w_021_035);
  and2 I091_112(w_091_112, w_048_011, w_038_193);
  not1 I091_117(w_091_117, w_044_743);
  nand2 I091_119(w_091_119, w_046_238, w_034_018);
  not1 I091_122(w_091_122, w_081_012);
  and2 I091_123(w_091_123, w_072_061, w_012_030);
  not1 I091_125(w_091_125, w_044_599);
  nand2 I091_127(w_091_127, w_015_614, w_052_006);
  and2 I091_129(w_091_129, w_087_048, w_054_073);
  and2 I091_133(w_091_133, w_087_216, w_021_209);
  and2 I091_134(w_091_134, w_011_474, w_062_591);
  or2  I091_135(w_091_135, w_031_494, w_080_192);
  nand2 I091_137(w_091_137, w_018_012, w_081_012);
  or2  I091_143(w_091_143, w_065_046, w_044_657);
  or2  I091_144(w_091_144, w_025_235, w_052_020);
  nand2 I091_151(w_091_151, w_087_088, w_021_114);
  nand2 I091_152(w_091_152, w_043_022, w_079_053);
  and2 I091_153(w_091_153, w_015_432, w_027_075);
  or2  I091_154(w_091_154, w_000_695, w_011_286);
  or2  I091_157(w_091_157, w_075_025, w_087_387);
  or2  I091_160(w_091_160, w_019_016, w_018_012);
  nand2 I091_161(w_091_161, w_005_276, w_027_121);
  not1 I091_162(w_091_162, w_007_215);
  nand2 I091_163(w_091_163, w_077_223, w_060_123);
  nand2 I091_164(w_091_164, w_056_466, w_031_101);
  not1 I091_166(w_091_166, w_032_409);
  and2 I091_169(w_091_169, w_004_171, w_005_171);
  and2 I091_170(w_091_170, w_045_338, w_047_119);
  or2  I091_176(w_091_176, w_045_292, w_050_295);
  and2 I092_001(w_092_001, w_040_449, w_035_044);
  or2  I092_009(w_092_009, w_042_233, w_046_338);
  and2 I092_011(w_092_011, w_037_162, w_047_270);
  and2 I092_027(w_092_027, w_052_008, w_031_558);
  and2 I092_029(w_092_029, w_018_008, w_054_155);
  or2  I092_032(w_092_032, w_043_031, w_043_029);
  nand2 I092_043(w_092_043, w_007_451, w_055_236);
  or2  I092_045(w_092_045, w_050_264, w_090_067);
  or2  I092_046(w_092_046, w_082_487, w_074_375);
  or2  I092_049(w_092_049, w_009_333, w_069_091);
  nand2 I092_050(w_092_050, w_020_102, w_011_150);
  and2 I092_059(w_092_059, w_001_008, w_002_183);
  not1 I092_062(w_092_062, w_069_068);
  and2 I092_068(w_092_068, w_088_089, w_077_107);
  nand2 I092_070(w_092_070, w_040_328, w_004_330);
  or2  I092_073(w_092_073, w_050_460, w_033_506);
  and2 I092_080(w_092_080, w_035_099, w_029_080);
  nand2 I092_088(w_092_088, w_049_222, w_075_011);
  not1 I092_089(w_092_089, w_037_172);
  or2  I092_107(w_092_107, w_013_065, w_054_131);
  and2 I092_112(w_092_112, w_058_540, w_054_013);
  not1 I092_131(w_092_131, w_084_007);
  and2 I092_151(w_092_151, w_014_194, w_085_327);
  nand2 I092_154(w_092_154, w_088_033, w_032_086);
  and2 I092_159(w_092_159, w_001_012, w_020_516);
  not1 I092_162(w_092_162, w_061_123);
  and2 I092_189(w_092_189, w_086_046, w_062_513);
  not1 I092_190(w_092_190, w_009_619);
  and2 I092_191(w_092_191, w_083_123, w_084_021);
  or2  I092_200(w_092_200, w_018_017, w_082_003);
  nand2 I092_203(w_092_203, w_047_238, w_083_193);
  nand2 I092_209(w_092_209, w_048_011, w_091_163);
  or2  I092_220(w_092_220, w_089_068, w_049_233);
  not1 I092_225(w_092_225, w_011_368);
  not1 I092_229(w_092_229, w_048_016);
  not1 I092_242(w_092_242, w_054_199);
  nand2 I092_264(w_092_264, w_084_033, w_041_023);
  nand2 I092_272(w_092_272, w_032_225, w_013_242);
  nand2 I092_277(w_092_277, w_071_091, w_049_239);
  and2 I092_287(w_092_287, w_062_253, w_015_497);
  not1 I092_292(w_092_292, w_088_069);
  and2 I092_307(w_092_307, w_068_204, w_014_084);
  and2 I092_324(w_092_324, w_066_558, w_035_055);
  and2 I092_331(w_092_331, w_016_002, w_015_604);
  and2 I092_360(w_092_360, w_032_569, w_025_162);
  not1 I092_377(w_092_377, w_056_242);
  and2 I092_391(w_092_391, w_013_322, w_009_010);
  not1 I092_412(w_092_412, w_046_702);
  or2  I092_429(w_092_429, w_050_085, w_035_037);
  not1 I092_439(w_092_439, w_058_060);
  or2  I092_447(w_092_447, w_041_128, w_005_147);
  nand2 I092_458(w_092_458, w_051_170, w_015_272);
  not1 I092_471(w_092_471, w_080_477);
  or2  I092_478(w_092_478, w_033_129, w_049_130);
  and2 I092_480(w_092_480, w_067_122, w_075_144);
  and2 I092_481(w_092_481, w_063_228, w_078_445);
  and2 I092_484(w_092_484, w_054_001, w_005_057);
  and2 I092_489(w_092_489, w_088_130, w_051_041);
  or2  I092_492(w_092_492, w_056_540, w_037_333);
  or2  I092_494(w_092_494, w_006_213, w_044_459);
  and2 I092_504(w_092_504, w_058_095, w_084_020);
  and2 I092_516(w_092_516, w_088_046, w_018_024);
  nand2 I092_530(w_092_530, w_035_045, w_015_529);
  and2 I092_548(w_092_548, w_043_013, w_037_051);
  nand2 I092_551(w_092_551, w_063_062, w_086_097);
  not1 I092_560(w_092_560, w_052_021);
  and2 I092_562(w_092_562, w_047_113, w_087_227);
  nand2 I092_563(w_092_563, w_082_425, w_041_359);
  and2 I092_572(w_092_572, w_015_129, w_037_158);
  not1 I092_580(w_092_580, w_072_034);
  or2  I092_588(w_092_588, w_027_134, w_085_199);
  not1 I092_595(w_092_595, w_058_171);
  not1 I092_609(w_092_609, w_017_029);
  and2 I092_610(w_092_610, w_017_567, w_081_000);
  not1 I092_628(w_092_628, w_064_207);
  nand2 I092_636(w_092_636, w_004_028, w_060_344);
  not1 I092_650(w_092_650, w_082_160);
  nand2 I092_673(w_092_673, w_002_540, w_044_055);
  and2 I092_690(w_092_690, w_035_122, w_011_232);
  nand2 I092_715(w_092_715, w_012_123, w_005_010);
  nand2 I092_723(w_092_725, w_092_738, w_092_724);
  and2 I092_724(w_092_726, w_062_177, w_092_725);
  or2  I092_725(w_092_724, w_092_726, w_051_167);
  and2 I092_726(w_092_731, w_038_591, w_092_730);
  or2  I092_727(w_092_732, w_019_012, w_092_731);
  and2 I092_728(w_092_733, w_092_732, w_057_070);
  or2  I092_729(w_092_734, w_092_733, w_003_042);
  or2  I092_730(w_092_735, w_010_498, w_092_734);
  and2 I092_731(w_092_736, w_092_735, w_034_031);
  not1 I092_732(w_092_730, w_092_725);
  and2 I092_733(w_092_738, w_018_007, w_092_736);
  not1 I093_006(w_093_006, w_078_464);
  not1 I093_016(w_093_016, w_053_088);
  and2 I093_028(w_093_028, w_017_508, w_022_177);
  or2  I093_032(w_093_032, w_070_530, w_015_113);
  and2 I093_035(w_093_035, w_062_666, w_021_056);
  not1 I093_041(w_093_041, w_077_127);
  not1 I093_043(w_093_043, w_052_009);
  nand2 I093_050(w_093_050, w_034_002, w_012_046);
  nand2 I093_054(w_093_054, w_001_002, w_069_104);
  nand2 I093_055(w_093_055, w_018_025, w_043_018);
  nand2 I093_057(w_093_057, w_043_002, w_024_026);
  or2  I093_059(w_093_059, w_075_077, w_068_075);
  not1 I093_060(w_093_060, w_083_057);
  not1 I093_067(w_093_067, w_085_306);
  and2 I093_073(w_093_073, w_069_014, w_029_061);
  or2  I093_077(w_093_077, w_010_733, w_085_085);
  not1 I093_080(w_093_080, w_090_531);
  not1 I093_081(w_093_081, w_045_088);
  not1 I093_084(w_093_084, w_057_013);
  and2 I093_086(w_093_086, w_081_010, w_065_304);
  not1 I093_088(w_093_088, w_092_636);
  nand2 I093_089(w_093_089, w_028_215, w_009_220);
  and2 I093_091(w_093_091, w_005_103, w_042_265);
  not1 I093_097(w_093_097, w_046_250);
  or2  I093_101(w_093_101, w_003_009, w_085_349);
  nand2 I093_105(w_093_105, w_077_321, w_064_328);
  and2 I093_119(w_093_119, w_001_009, w_080_032);
  and2 I093_123(w_093_123, w_077_123, w_057_140);
  not1 I093_128(w_093_128, w_041_623);
  not1 I093_132(w_093_132, w_037_077);
  not1 I093_133(w_093_133, w_066_594);
  or2  I093_143(w_093_143, w_017_648, w_020_115);
  not1 I093_151(w_093_151, w_005_150);
  and2 I093_162(w_093_162, w_038_106, w_049_303);
  not1 I093_177(w_093_177, w_028_470);
  not1 I093_178(w_093_178, w_081_017);
  not1 I093_180(w_093_180, w_057_081);
  and2 I093_186(w_093_186, w_036_076, w_022_290);
  not1 I093_200(w_093_200, w_037_186);
  not1 I093_208(w_093_208, w_084_037);
  or2  I093_217(w_093_217, w_054_231, w_061_106);
  nand2 I093_224(w_093_224, w_050_322, w_007_403);
  or2  I093_225(w_093_225, w_041_668, w_046_339);
  and2 I093_239(w_093_239, w_061_073, w_074_186);
  or2  I093_245(w_093_245, w_027_140, w_008_755);
  or2  I093_252(w_093_252, w_041_594, w_038_100);
  nand2 I093_256(w_093_256, w_092_027, w_083_067);
  not1 I093_270(w_093_270, w_076_321);
  and2 I093_321(w_093_321, w_071_034, w_046_062);
  or2  I093_332(w_093_332, w_061_051, w_028_135);
  not1 I093_339(w_093_339, w_073_068);
  or2  I093_354(w_093_354, w_004_141, w_084_039);
  and2 I093_360(w_093_360, w_062_057, w_049_017);
  or2  I093_362(w_093_362, w_041_010, w_058_208);
  nand2 I093_371(w_093_371, w_048_009, w_020_565);
  and2 I093_389(w_093_389, w_060_126, w_091_161);
  or2  I093_390(w_093_390, w_091_012, w_068_360);
  or2  I093_391(w_093_391, w_015_431, w_049_209);
  or2  I093_393(w_093_393, w_070_216, w_071_289);
  nand2 I093_395(w_093_395, w_005_013, w_084_048);
  nand2 I093_409(w_093_409, w_082_130, w_046_264);
  or2  I093_413(w_093_413, w_082_104, w_017_591);
  not1 I093_417(w_093_417, w_041_432);
  not1 I093_420(w_093_420, w_072_175);
  or2  I093_421(w_093_421, w_088_022, w_074_044);
  not1 I093_430(w_093_430, w_058_660);
  and2 I093_442(w_093_442, w_063_111, w_053_049);
  or2  I093_448(w_093_448, w_028_528, w_045_000);
  or2  I093_458(w_093_458, w_050_099, w_034_043);
  not1 I093_497(w_093_497, w_016_006);
  and2 I093_504(w_093_504, w_018_040, w_071_303);
  nand2 I093_559(w_093_561, w_056_371, w_093_560);
  and2 I093_560(w_093_562, w_089_045, w_093_561);
  and2 I093_561(w_093_563, w_010_331, w_093_562);
  and2 I093_562(w_093_560, w_009_250, w_093_563);
  and2 I093_563(w_092_728, w_093_362, w_092_724);
  nand2 I094_006(w_094_006, w_089_149, w_081_016);
  and2 I094_009(w_094_009, w_012_010, w_039_242);
  and2 I094_021(w_094_021, w_024_060, w_086_312);
  not1 I094_027(w_094_027, w_039_127);
  not1 I094_038(w_094_038, w_057_061);
  and2 I094_043(w_094_043, w_080_289, w_041_131);
  nand2 I094_044(w_094_044, w_056_048, w_091_123);
  or2  I094_051(w_094_051, w_072_064, w_071_143);
  and2 I094_052(w_094_052, w_065_296, w_057_229);
  not1 I094_056(w_094_056, w_018_019);
  nand2 I094_057(w_094_057, w_003_045, w_062_245);
  not1 I094_064(w_094_064, w_018_032);
  and2 I094_079(w_094_079, w_067_343, w_038_499);
  or2  I094_083(w_094_083, w_012_330, w_068_265);
  and2 I094_095(w_094_095, w_062_206, w_000_153);
  not1 I094_101(w_094_101, w_081_007);
  nand2 I094_110(w_094_110, w_064_125, w_047_090);
  and2 I094_114(w_094_114, w_085_202, w_055_254);
  and2 I094_116(w_094_116, w_060_305, w_015_302);
  not1 I094_120(w_094_120, w_070_293);
  not1 I094_138(w_094_138, w_003_017);
  not1 I094_150(w_094_150, w_002_190);
  nand2 I094_159(w_094_159, w_091_040, w_093_371);
  or2  I094_162(w_094_162, w_022_164, w_082_090);
  or2  I094_167(w_094_167, w_026_298, w_035_088);
  not1 I094_173(w_094_173, w_033_275);
  and2 I094_182(w_094_182, w_072_161, w_015_081);
  or2  I094_193(w_094_193, w_023_003, w_041_583);
  and2 I094_195(w_094_195, w_059_162, w_003_007);
  not1 I094_222(w_094_222, w_010_585);
  nand2 I094_234(w_094_234, w_072_208, w_011_410);
  and2 I094_246(w_094_246, w_026_655, w_008_353);
  or2  I094_267(w_094_267, w_011_517, w_000_556);
  nand2 I094_271(w_094_271, w_038_304, w_046_422);
  not1 I094_286(w_094_286, w_089_089);
  not1 I094_288(w_094_288, w_002_513);
  not1 I094_296(w_094_296, w_003_063);
  or2  I094_299(w_094_299, w_036_141, w_016_006);
  nand2 I094_317(w_094_317, w_058_256, w_050_093);
  nand2 I094_336(w_094_336, w_006_187, w_037_157);
  and2 I094_344(w_094_344, w_068_209, w_054_467);
  or2  I094_363(w_094_363, w_058_092, w_055_097);
  not1 I094_370(w_094_370, w_003_073);
  nand2 I094_373(w_094_373, w_066_578, w_040_032);
  or2  I094_376(w_094_376, w_093_057, w_089_258);
  nand2 I094_380(w_094_380, w_085_338, w_010_123);
  not1 I094_381(w_094_381, w_066_489);
  nand2 I094_386(w_094_386, w_045_287, w_054_319);
  nand2 I094_387(w_094_387, w_090_442, w_059_170);
  and2 I094_399(w_094_399, w_075_034, w_058_596);
  nand2 I094_419(w_094_419, w_068_224, w_035_080);
  nand2 I094_421(w_094_421, w_000_213, w_029_091);
  or2  I094_432(w_094_432, w_072_102, w_014_116);
  not1 I094_434(w_094_434, w_025_161);
  not1 I094_440(w_094_440, w_074_232);
  nand2 I094_444(w_094_444, w_032_045, w_051_148);
  or2  I094_449(w_094_449, w_001_024, w_026_028);
  or2  I094_462(w_094_462, w_030_244, w_077_412);
  not1 I094_469(w_094_469, w_010_149);
  not1 I094_475(w_094_475, w_061_356);
  and2 I094_514(w_094_514, w_074_000, w_008_150);
  not1 I094_522(w_094_522, w_014_022);
  nand2 I094_527(w_094_527, w_092_728, w_049_024);
  or2  I094_534(w_094_534, w_066_045, w_051_333);
  nand2 I094_542(w_094_542, w_085_299, w_029_073);
  or2  I094_544(w_094_544, w_012_045, w_048_017);
  nand2 I094_545(w_094_545, w_047_077, w_061_283);
  not1 I094_546(w_094_546, w_032_313);
  not1 I094_564(w_094_564, w_064_327);
  not1 I094_574(w_094_574, w_042_180);
  nand2 I094_587(w_094_587, w_016_004, w_043_025);
  not1 I094_599(w_094_599, w_079_041);
  nand2 I094_600(w_094_600, w_011_273, w_020_387);
  or2  I094_607(w_094_607, w_034_033, w_086_089);
  or2  I094_609(w_094_609, w_012_311, w_092_045);
  nand2 I094_610(w_094_610, w_062_508, w_040_327);
  and2 I094_624(w_094_624, w_042_035, w_000_525);
  nand2 I094_662(w_094_664, w_094_663, w_084_047);
  nand2 I094_663(w_094_665, w_094_664, w_017_292);
  not1 I094_664(w_094_666, w_094_665);
  and2 I094_665(w_094_667, w_094_666, w_040_228);
  or2  I094_666(w_094_663, w_094_667, w_019_012);
  and2 I094_667(w_093_565, w_052_024, w_093_560);
  or2  I095_000(w_095_000, w_092_429, w_018_042);
  not1 I095_001(w_095_001, w_001_033);
  or2  I095_002(w_095_002, w_042_331, w_074_360);
  not1 I095_003(w_095_003, w_070_071);
  or2  I095_004(w_095_004, w_082_148, w_012_036);
  not1 I095_005(w_095_005, w_013_346);
  and2 I095_006(w_095_006, w_006_165, w_075_062);
  and2 I095_008(w_095_008, w_028_029, w_052_042);
  and2 I095_010(w_095_010, w_025_187, w_052_008);
  or2  I095_012(w_095_012, w_022_352, w_065_372);
  or2  I095_014(w_095_014, w_026_187, w_085_017);
  and2 I095_018(w_095_018, w_091_152, w_089_061);
  nand2 I095_019(w_095_019, w_068_231, w_084_024);
  not1 I095_021(w_095_021, w_022_252);
  and2 I095_022(w_095_022, w_074_288, w_015_524);
  not1 I095_023(w_095_023, w_047_294);
  nand2 I095_026(w_095_026, w_089_140, w_031_346);
  nand2 I095_027(w_095_027, w_017_263, w_073_402);
  or2  I095_029(w_095_029, w_059_405, w_024_206);
  nand2 I095_030(w_095_030, w_067_239, w_081_012);
  not1 I095_031(w_095_031, w_015_043);
  or2  I095_033(w_095_033, w_030_274, w_068_334);
  and2 I095_034(w_095_034, w_082_511, w_053_097);
  or2  I095_036(w_095_036, w_042_041, w_000_319);
  and2 I095_038(w_095_038, w_074_340, w_056_090);
  and2 I095_039(w_095_039, w_094_440, w_054_234);
  or2  I095_040(w_095_040, w_035_092, w_077_151);
  nand2 I095_041(w_095_041, w_017_536, w_079_030);
  and2 I095_042(w_095_042, w_058_271, w_059_165);
  not1 I095_043(w_095_043, w_036_059);
  not1 I095_046(w_095_046, w_086_122);
  nand2 I095_047(w_095_047, w_023_122, w_033_488);
  or2  I095_049(w_095_049, w_070_294, w_080_245);
  and2 I095_051(w_095_051, w_060_343, w_020_521);
  and2 I095_052(w_095_052, w_093_565, w_017_055);
  not1 I095_053(w_095_053, w_065_563);
  and2 I095_054(w_095_054, w_004_093, w_068_001);
  and2 I095_055(w_095_055, w_080_472, w_051_263);
  not1 I095_056(w_095_056, w_036_060);
  not1 I095_057(w_095_057, w_054_126);
  and2 I095_059(w_094_669, w_072_129, w_094_663);
  or2  I096_000(w_096_000, w_009_199, w_090_195);
  not1 I096_001(w_096_001, w_028_541);
  or2  I096_002(w_096_002, w_045_230, w_044_000);
  nand2 I096_003(w_096_003, w_094_669, w_064_087);
  and2 I096_004(w_096_004, w_094_381, w_037_085);
  nand2 I096_005(w_096_005, w_082_576, w_012_051);
  nand2 I097_002(w_097_002, w_072_152, w_086_032);
  not1 I097_004(w_097_004, w_022_001);
  not1 I097_007(w_097_007, w_079_023);
  not1 I097_009(w_097_009, w_055_097);
  or2  I097_012(w_097_012, w_091_094, w_088_002);
  not1 I097_016(w_097_016, w_052_046);
  or2  I097_033(w_097_033, w_011_235, w_027_026);
  or2  I097_035(w_097_035, w_017_094, w_015_439);
  and2 I097_038(w_097_038, w_027_125, w_079_030);
  not1 I097_039(w_097_039, w_047_134);
  nand2 I097_042(w_097_042, w_008_366, w_040_468);
  and2 I097_048(w_097_048, w_024_208, w_033_555);
  not1 I097_049(w_097_049, w_007_093);
  or2  I097_056(w_097_056, w_067_255, w_065_248);
  nand2 I097_061(w_097_061, w_031_413, w_067_046);
  not1 I097_063(w_097_063, w_028_129);
  not1 I097_070(w_097_070, w_060_016);
  or2  I097_077(w_097_077, w_040_348, w_019_018);
  nand2 I097_082(w_097_082, w_063_175, w_090_310);
  or2  I097_085(w_097_085, w_062_390, w_001_009);
  or2  I097_088(w_097_088, w_077_592, w_040_646);
  nand2 I097_090(w_097_090, w_060_381, w_083_021);
  not1 I097_102(w_097_102, w_075_025);
  or2  I097_105(w_097_105, w_084_026, w_036_071);
  or2  I097_108(w_097_108, w_087_098, w_007_103);
  not1 I097_118(w_097_118, w_028_098);
  or2  I097_121(w_097_121, w_001_030, w_030_138);
  or2  I097_122(w_097_122, w_061_148, w_060_109);
  and2 I097_125(w_097_125, w_004_110, w_049_135);
  nand2 I097_130(w_097_130, w_000_403, w_081_020);
  not1 I097_131(w_097_131, w_037_173);
  or2  I097_135(w_097_135, w_025_174, w_025_191);
  or2  I097_139(w_097_139, w_019_005, w_005_231);
  nand2 I097_142(w_097_142, w_034_007, w_015_612);
  or2  I097_144(w_097_144, w_034_074, w_066_029);
  or2  I097_153(w_097_153, w_061_307, w_092_439);
  nand2 I097_166(w_097_166, w_088_070, w_086_119);
  not1 I097_175(w_097_175, w_072_003);
  and2 I097_179(w_097_179, w_087_310, w_026_702);
  not1 I097_180(w_097_180, w_057_053);
  and2 I097_189(w_097_189, w_033_656, w_084_008);
  nand2 I097_195(w_097_195, w_095_056, w_026_331);
  or2  I097_201(w_097_201, w_004_068, w_026_182);
  nand2 I097_205(w_097_205, w_046_429, w_072_059);
  or2  I097_207(w_097_207, w_000_102, w_021_032);
  nand2 I097_212(w_097_212, w_036_237, w_073_088);
  and2 I097_224(w_097_224, w_038_359, w_087_189);
  nand2 I097_225(w_097_225, w_082_199, w_076_405);
  and2 I097_252(w_097_252, w_049_192, w_029_102);
  not1 I097_303(w_097_303, w_054_106);
  nand2 I097_331(w_097_331, w_054_173, w_079_018);
  nand2 I097_335(w_097_335, w_001_020, w_077_232);
  and2 I097_360(w_097_360, w_013_470, w_065_512);
  nand2 I097_366(w_097_366, w_091_000, w_079_053);
  or2  I097_373(w_097_373, w_010_700, w_007_123);
  and2 I097_374(w_097_374, w_073_507, w_033_619);
  not1 I097_393(w_097_393, w_007_285);
  and2 I097_430(w_097_430, w_038_011, w_013_130);
  nand2 I097_471(w_097_471, w_010_127, w_005_066);
  not1 I097_480(w_097_480, w_070_083);
  or2  I097_492(w_097_492, w_028_000, w_046_209);
  and2 I097_502(w_097_502, w_046_659, w_044_721);
  or2  I097_504(w_097_504, w_044_510, w_087_190);
  not1 I097_507(w_097_507, w_090_218);
  not1 I097_514(w_097_514, w_025_243);
  nand2 I097_521(w_097_521, w_089_300, w_094_110);
  nand2 I097_526(w_097_526, w_083_190, w_079_000);
  and2 I097_548(w_097_548, w_076_461, w_003_050);
  or2  I097_553(w_097_553, w_029_107, w_093_105);
  or2  I097_566(w_097_566, w_069_065, w_024_447);
  not1 I097_570(w_097_570, w_088_080);
  or2  I098_000(w_098_000, w_017_228, w_089_070);
  or2  I098_001(w_098_001, w_057_057, w_083_040);
  and2 I098_003(w_098_003, w_007_124, w_097_548);
  nand2 I098_004(w_098_004, w_016_007, w_075_037);
  not1 I098_005(w_098_005, w_024_088);
  or2  I098_008(w_098_008, w_010_353, w_052_031);
  nand2 I098_009(w_098_009, w_014_144, w_031_088);
  or2  I098_010(w_098_010, w_085_092, w_082_383);
  or2  I098_011(w_098_011, w_059_734, w_053_004);
  nand2 I098_012(w_098_012, w_052_027, w_062_329);
  nand2 I098_013(w_098_013, w_023_156, w_077_444);
  not1 I098_014(w_098_014, w_047_276);
  nand2 I098_015(w_098_015, w_055_094, w_028_088);
  nand2 I098_016(w_098_016, w_059_125, w_010_388);
  nand2 I098_017(w_098_017, w_092_049, w_078_016);
  not1 I098_018(w_098_018, w_087_102);
  or2  I098_019(w_098_019, w_041_630, w_070_069);
  or2  I098_020(w_098_020, w_093_225, w_089_217);
  and2 I098_022(w_098_022, w_052_042, w_045_225);
  not1 I098_024(w_098_024, w_061_300);
  and2 I098_025(w_098_025, w_006_133, w_068_041);
  not1 I098_027(w_098_027, w_011_467);
  or2  I098_028(w_098_028, w_005_016, w_043_012);
  or2  I098_031(w_098_031, w_011_361, w_007_253);
  nand2 I098_032(w_098_032, w_075_062, w_046_024);
  and2 I098_033(w_098_033, w_066_052, w_058_005);
  and2 I098_034(w_098_034, w_078_142, w_010_010);
  not1 I098_035(w_098_035, w_067_171);
  not1 I098_036(w_098_036, w_081_005);
  and2 I098_038(w_098_038, w_019_004, w_097_189);
  not1 I098_040(w_098_040, w_058_479);
  and2 I098_041(w_098_041, w_077_110, w_063_149);
  not1 I098_042(w_098_042, w_057_182);
  or2  I098_043(w_098_043, w_061_467, w_032_121);
  and2 I098_044(w_098_044, w_040_705, w_041_011);
  or2  I098_045(w_098_045, w_048_019, w_040_553);
  or2  I098_046(w_098_046, w_033_183, w_030_208);
  or2  I098_047(w_098_047, w_088_020, w_071_316);
  and2 I098_048(w_098_048, w_090_011, w_070_381);
  not1 I098_050(w_098_050, w_038_077);
  and2 I098_052(w_098_052, w_062_151, w_097_002);
  not1 I098_053(w_098_053, w_029_071);
  and2 I098_055(w_098_055, w_052_017, w_008_011);
  or2  I098_057(w_098_057, w_053_035, w_085_230);
  not1 I098_058(w_098_058, w_023_018);
  not1 I098_059(w_098_059, w_009_372);
  and2 I098_061(w_098_061, w_010_413, w_080_171);
  or2  I098_062(w_098_062, w_079_047, w_027_058);
  not1 I098_063(w_098_063, w_040_481);
  or2  I098_065(w_098_065, w_011_033, w_020_508);
  not1 I098_068(w_098_068, w_008_076);
  and2 I098_069(w_098_069, w_015_105, w_004_463);
  or2  I098_071(w_098_071, w_064_049, w_057_001);
  nand2 I098_074(w_098_074, w_018_015, w_011_027);
  not1 I099_001(w_099_001, w_076_168);
  and2 I099_002(w_099_002, w_009_051, w_064_134);
  or2  I099_003(w_099_003, w_025_111, w_095_014);
  or2  I099_011(w_099_011, w_098_008, w_096_002);
  and2 I099_015(w_099_015, w_084_042, w_046_356);
  nand2 I099_019(w_099_019, w_028_205, w_000_221);
  or2  I099_025(w_099_025, w_030_121, w_028_123);
  and2 I099_036(w_099_036, w_025_061, w_089_075);
  and2 I099_037(w_099_037, w_049_363, w_022_267);
  not1 I099_044(w_099_044, w_066_281);
  or2  I099_047(w_099_047, w_014_026, w_036_206);
  nand2 I099_051(w_099_051, w_015_259, w_005_299);
  nand2 I099_053(w_099_053, w_015_132, w_001_007);
  nand2 I099_054(w_099_054, w_037_017, w_002_494);
  and2 I099_055(w_099_055, w_018_025, w_071_284);
  nand2 I099_057(w_099_057, w_038_021, w_080_303);
  nand2 I099_058(w_099_058, w_096_001, w_029_082);
  not1 I099_059(w_099_059, w_047_283);
  not1 I099_062(w_099_062, w_002_078);
  or2  I099_068(w_099_068, w_083_044, w_016_006);
  or2  I099_070(w_099_070, w_091_111, w_041_504);
  or2  I099_071(w_099_071, w_070_080, w_045_224);
  not1 I099_075(w_099_075, w_062_549);
  nand2 I099_077(w_099_077, w_041_576, w_031_386);
  and2 I099_078(w_099_078, w_077_610, w_054_173);
  not1 I099_081(w_099_081, w_063_251);
  and2 I099_087(w_099_087, w_018_019, w_029_023);
  and2 I099_088(w_099_088, w_090_392, w_002_706);
  and2 I099_091(w_099_091, w_078_475, w_045_024);
  or2  I099_093(w_099_093, w_075_044, w_098_009);
  nand2 I099_101(w_099_101, w_067_232, w_031_555);
  not1 I099_107(w_099_107, w_056_520);
  and2 I099_111(w_099_111, w_017_078, w_077_385);
  nand2 I099_113(w_099_113, w_034_025, w_075_063);
  not1 I099_114(w_099_114, w_023_017);
  not1 I099_123(w_099_123, w_060_296);
  not1 I099_131(w_099_131, w_023_071);
  nand2 I099_133(w_099_133, w_031_469, w_001_029);
  or2  I099_135(w_099_135, w_094_138, w_036_158);
  nand2 I099_136(w_099_136, w_042_092, w_093_054);
  not1 I099_141(w_099_141, w_059_639);
  or2  I099_148(w_099_148, w_046_104, w_027_142);
  not1 I099_150(w_099_150, w_074_045);
  or2  I099_159(w_099_159, w_017_080, w_071_105);
  or2  I099_163(w_099_163, w_076_033, w_070_573);
  not1 I099_169(w_099_169, w_057_296);
  or2  I099_172(w_099_172, w_028_021, w_007_144);
  and2 I099_173(w_099_173, w_032_300, w_080_290);
  nand2 I099_174(w_099_174, w_075_009, w_077_479);
  not1 I099_178(w_099_178, w_051_067);
  and2 I099_180(w_099_180, w_016_003, w_054_239);
  nand2 I099_188(w_099_188, w_070_396, w_055_022);
  or2  I099_192(w_099_192, w_091_033, w_017_234);
  nand2 I099_205(w_099_205, w_048_014, w_023_108);
  and2 I099_213(w_099_213, w_015_296, w_074_345);
  and2 I099_222(w_099_222, w_074_254, w_020_165);
  nand2 I099_223(w_099_223, w_073_512, w_008_183);
  and2 I099_229(w_099_229, w_030_293, w_096_002);
  or2  I099_240(w_099_240, w_049_305, w_002_188);
  not1 I099_248(w_099_248, w_079_018);
  or2  I099_256(w_099_256, w_061_437, w_016_008);
  and2 I099_257(w_099_257, w_066_058, w_090_035);
  or2  I099_261(w_099_261, w_065_016, w_091_129);
  or2  I099_262(w_099_262, w_071_265, w_002_557);
  not1 I099_263(w_099_263, w_063_194);
  and2 I099_274(w_099_274, w_019_014, w_009_430);
  or2  I099_276(w_099_276, w_013_515, w_076_181);
  nand2 I099_278(w_099_278, w_074_300, w_001_004);
  and2 I099_291(w_099_291, w_044_128, w_066_013);
  nand2 I099_301(w_099_303, w_020_188, w_099_302);
  nand2 I099_302(w_099_304, w_099_303, w_051_199);
  nand2 I099_303(w_099_305, w_051_045, w_099_304);
  nand2 I099_304(w_099_306, w_099_305, w_031_177);
  and2 I099_305(w_099_307, w_086_313, w_099_306);
  or2  I099_306(w_099_308, w_073_691, w_099_307);
  nand2 I099_307(w_099_309, w_099_308, w_064_005);
  nand2 I099_308(w_099_310, w_099_309, w_046_593);
  not1 I099_309(w_099_311, w_099_310);
  nand2 I099_310(w_099_312, w_099_311, w_028_029);
  and2 I099_311(w_099_313, w_099_329, w_099_312);
  not1 I099_312(w_099_302, w_099_313);
  not1 I099_313(w_099_318, w_099_317);
  not1 I099_314(w_099_319, w_099_318);
  or2  I099_315(w_099_320, w_097_016, w_099_319);
  or2  I099_316(w_099_321, w_099_320, w_031_599);
  or2  I099_317(w_099_322, w_068_321, w_099_321);
  and2 I099_318(w_099_323, w_099_322, w_073_714);
  and2 I099_319(w_099_324, w_060_262, w_099_323);
  or2  I099_320(w_099_325, w_068_307, w_099_324);
  and2 I099_321(w_099_326, w_099_325, w_051_307);
  and2 I099_322(w_099_327, w_099_326, w_056_089);
  not1 I099_323(w_099_317, w_099_313);
  and2 I099_324(w_099_329, w_079_045, w_099_327);
  nand2 I100_002(w_100_002, w_030_192, w_065_348);
  nand2 I100_007(w_100_007, w_096_005, w_029_079);
  not1 I100_008(w_100_008, w_012_082);
  or2  I100_010(w_100_010, w_037_318, w_036_239);
  or2  I100_012(w_100_012, w_013_088, w_000_209);
  or2  I100_013(w_100_013, w_060_222, w_038_302);
  or2  I100_014(w_100_014, w_086_007, w_026_490);
  not1 I100_018(w_100_018, w_056_016);
  nand2 I100_019(w_100_019, w_045_009, w_060_331);
  or2  I100_021(w_100_021, w_076_050, w_096_001);
  and2 I100_022(w_100_022, w_086_189, w_011_018);
  and2 I100_024(w_100_024, w_034_036, w_091_042);
  nand2 I100_030(w_100_030, w_021_219, w_038_247);
  or2  I100_031(w_100_031, w_024_208, w_096_002);
  not1 I100_036(w_100_036, w_051_323);
  or2  I100_037(w_100_037, w_072_292, w_035_088);
  not1 I100_038(w_100_038, w_059_012);
  and2 I100_044(w_100_044, w_012_254, w_008_284);
  or2  I100_046(w_100_046, w_030_382, w_080_096);
  or2  I100_049(w_100_049, w_090_131, w_074_327);
  and2 I100_051(w_100_051, w_005_044, w_099_276);
  and2 I100_053(w_100_053, w_000_128, w_059_049);
  nand2 I100_055(w_100_055, w_047_206, w_025_155);
  and2 I100_056(w_100_056, w_049_263, w_043_006);
  not1 I100_057(w_100_057, w_088_003);
  or2  I100_058(w_100_058, w_039_280, w_092_088);
  not1 I100_060(w_100_060, w_065_152);
  or2  I100_061(w_100_061, w_015_400, w_034_025);
  or2  I100_063(w_100_063, w_098_055, w_083_011);
  or2  I100_065(w_100_065, w_081_015, w_077_361);
  not1 I100_066(w_100_066, w_017_315);
  nand2 I100_071(w_100_071, w_022_153, w_085_309);
  or2  I100_074(w_100_074, w_088_136, w_030_155);
  and2 I100_077(w_100_077, w_092_715, w_072_266);
  not1 I100_078(w_100_078, w_009_129);
  and2 I100_080(w_100_080, w_009_520, w_007_175);
  not1 I100_081(w_100_081, w_095_019);
  and2 I100_082(w_100_082, w_029_004, w_081_015);
  and2 I100_084(w_100_084, w_042_312, w_072_057);
  or2  I100_085(w_100_085, w_038_064, w_002_320);
  not1 I100_086(w_100_086, w_083_147);
  not1 I100_087(w_100_087, w_092_458);
  and2 I100_092(w_100_092, w_045_084, w_027_055);
  nand2 I100_093(w_100_093, w_010_403, w_093_354);
  not1 I100_094(w_100_094, w_082_162);
  not1 I100_095(w_100_095, w_019_001);
  nand2 I100_096(w_100_096, w_085_048, w_017_085);
  and2 I100_100(w_100_100, w_068_225, w_074_194);
  nand2 I100_106(w_100_106, w_095_053, w_035_023);
  and2 I100_109(w_100_109, w_091_028, w_098_034);
  or2  I100_113(w_100_113, w_068_081, w_056_692);
  or2  I100_115(w_100_115, w_065_517, w_070_083);
  and2 I100_116(w_100_116, w_053_108, w_027_126);
  or2  I100_120(w_100_120, w_025_054, w_097_331);
  or2  I100_121(w_100_121, w_015_596, w_014_143);
  and2 I100_125(w_100_125, w_094_267, w_049_204);
  nand2 I100_127(w_100_127, w_047_008, w_041_414);
  nand2 I100_130(w_100_130, w_099_091, w_093_097);
  and2 I101_003(w_101_003, w_079_004, w_089_135);
  nand2 I101_004(w_101_004, w_006_003, w_083_158);
  or2  I101_006(w_101_006, w_070_174, w_069_063);
  nand2 I101_008(w_101_008, w_091_074, w_029_004);
  nand2 I101_020(w_101_020, w_057_146, w_070_489);
  not1 I101_038(w_101_038, w_029_091);
  nand2 I101_049(w_101_049, w_084_009, w_066_103);
  or2  I101_050(w_101_050, w_019_010, w_058_140);
  and2 I101_056(w_101_056, w_071_096, w_000_362);
  or2  I101_063(w_101_063, w_000_545, w_003_054);
  and2 I101_066(w_101_066, w_080_007, w_039_697);
  not1 I101_070(w_101_070, w_060_098);
  or2  I101_077(w_101_077, w_060_125, w_018_041);
  and2 I101_083(w_101_083, w_024_020, w_008_582);
  or2  I101_085(w_101_085, w_081_022, w_044_199);
  not1 I101_089(w_101_089, w_064_155);
  and2 I101_090(w_101_090, w_075_000, w_059_101);
  nand2 I101_092(w_101_092, w_002_195, w_007_088);
  and2 I101_094(w_101_094, w_099_107, w_069_107);
  and2 I101_095(w_101_095, w_067_137, w_042_316);
  nand2 I101_098(w_101_098, w_096_001, w_022_220);
  or2  I101_104(w_101_104, w_093_091, w_035_002);
  and2 I101_107(w_101_107, w_052_033, w_100_116);
  not1 I101_121(w_101_121, w_046_222);
  and2 I101_122(w_101_122, w_062_249, w_073_017);
  or2  I101_124(w_101_124, w_007_110, w_086_195);
  or2  I101_130(w_101_130, w_066_482, w_043_030);
  or2  I101_135(w_101_135, w_097_212, w_095_021);
  and2 I101_139(w_101_139, w_062_177, w_095_049);
  or2  I101_143(w_101_143, w_051_063, w_033_182);
  nand2 I101_156(w_101_156, w_089_060, w_096_002);
  nand2 I101_158(w_101_158, w_095_051, w_004_138);
  or2  I101_166(w_101_166, w_045_405, w_012_345);
  nand2 I101_168(w_101_168, w_021_086, w_089_096);
  or2  I101_170(w_101_170, w_063_010, w_085_255);
  not1 I101_171(w_101_171, w_013_352);
  and2 I101_176(w_101_176, w_001_029, w_046_427);
  not1 I101_188(w_101_188, w_054_109);
  and2 I101_194(w_101_194, w_046_576, w_097_009);
  or2  I101_207(w_101_207, w_024_545, w_040_616);
  or2  I101_209(w_101_209, w_074_348, w_004_288);
  and2 I101_214(w_101_214, w_057_187, w_045_057);
  or2  I101_223(w_101_223, w_087_117, w_063_183);
  nand2 I101_238(w_101_238, w_043_030, w_094_624);
  or2  I101_243(w_101_243, w_014_229, w_050_446);
  nand2 I101_244(w_101_244, w_085_045, w_028_463);
  or2  I101_246(w_101_246, w_016_008, w_045_012);
  not1 I101_247(w_101_247, w_024_530);
  nand2 I101_253(w_101_253, w_006_113, w_024_549);
  and2 I101_258(w_101_258, w_036_269, w_078_130);
  nand2 I101_261(w_101_261, w_080_225, w_063_397);
  not1 I101_266(w_101_266, w_065_172);
  and2 I101_269(w_101_269, w_042_159, w_035_055);
  nand2 I101_272(w_101_272, w_057_185, w_047_054);
  or2  I101_280(w_101_280, w_002_270, w_031_497);
  or2  I101_283(w_101_283, w_065_547, w_007_096);
  nand2 I101_284(w_101_284, w_039_119, w_051_189);
  or2  I101_285(w_101_285, w_023_105, w_027_057);
  not1 I101_293(w_101_293, w_005_182);
  nand2 I101_294(w_101_294, w_006_016, w_064_285);
  or2  I101_303(w_101_303, w_067_328, w_003_073);
  nand2 I101_307(w_101_307, w_055_313, w_007_036);
  not1 I101_312(w_101_314, w_101_313);
  nand2 I101_313(w_101_315, w_098_015, w_101_314);
  or2  I101_314(w_101_316, w_052_027, w_101_315);
  and2 I101_315(w_101_317, w_058_030, w_101_316);
  or2  I101_316(w_101_313, w_101_317, w_101_325);
  nand2 I101_317(w_101_322, w_101_321, w_012_079);
  and2 I101_318(w_101_323, w_101_322, w_056_241);
  not1 I101_319(w_101_321, w_101_313);
  and2 I101_320(w_101_325, w_005_191, w_101_323);
  nand2 I102_014(w_102_014, w_067_049, w_081_010);
  not1 I102_022(w_102_022, w_037_047);
  not1 I102_025(w_102_025, w_038_397);
  not1 I102_028(w_102_028, w_014_054);
  nand2 I102_035(w_102_035, w_096_000, w_033_475);
  not1 I102_036(w_102_036, w_010_151);
  and2 I102_042(w_102_042, w_054_020, w_099_222);
  or2  I102_047(w_102_047, w_074_322, w_051_185);
  nand2 I102_050(w_102_050, w_025_078, w_072_163);
  or2  I102_060(w_102_060, w_040_067, w_038_434);
  nand2 I102_068(w_102_068, w_087_013, w_096_004);
  and2 I102_070(w_102_070, w_004_012, w_029_002);
  and2 I102_076(w_102_076, w_090_489, w_038_288);
  and2 I102_093(w_102_093, w_076_220, w_027_055);
  not1 I102_097(w_102_097, w_014_001);
  not1 I102_115(w_102_115, w_071_022);
  and2 I102_116(w_102_116, w_051_150, w_013_140);
  or2  I102_123(w_102_123, w_003_019, w_089_191);
  or2  I102_133(w_102_133, w_011_481, w_093_332);
  not1 I102_144(w_102_144, w_044_713);
  not1 I102_152(w_102_152, w_065_320);
  nand2 I102_181(w_102_181, w_004_090, w_004_270);
  and2 I102_183(w_102_183, w_011_050, w_061_264);
  not1 I102_188(w_102_188, w_098_050);
  nand2 I102_193(w_102_193, w_078_103, w_042_005);
  not1 I102_195(w_102_195, w_027_059);
  nand2 I102_199(w_102_199, w_047_116, w_093_430);
  not1 I102_204(w_102_204, w_001_015);
  or2  I102_226(w_102_226, w_049_277, w_013_088);
  and2 I102_229(w_102_229, w_087_253, w_090_080);
  or2  I102_246(w_102_246, w_017_385, w_085_298);
  and2 I102_248(w_102_248, w_060_289, w_069_226);
  nand2 I102_250(w_102_250, w_036_307, w_061_213);
  not1 I102_252(w_102_252, w_066_023);
  not1 I102_274(w_102_274, w_023_111);
  not1 I102_282(w_102_282, w_073_009);
  and2 I102_304(w_102_304, w_061_356, w_082_041);
  and2 I102_308(w_102_308, w_062_149, w_008_336);
  nand2 I102_316(w_102_316, w_088_028, w_030_016);
  not1 I102_329(w_102_329, w_056_037);
  and2 I102_333(w_102_333, w_001_025, w_072_149);
  nand2 I102_337(w_102_337, w_071_217, w_008_190);
  not1 I102_345(w_102_345, w_012_230);
  nand2 I102_364(w_102_364, w_090_016, w_005_047);
  or2  I102_368(w_102_368, w_046_009, w_035_021);
  nand2 I102_392(w_102_392, w_046_041, w_065_307);
  or2  I102_421(w_102_421, w_017_087, w_047_309);
  and2 I102_424(w_102_424, w_084_025, w_006_111);
  nand2 I102_436(w_102_436, w_061_205, w_009_071);
  not1 I102_442(w_102_442, w_097_061);
  or2  I102_445(w_102_445, w_053_026, w_048_014);
  not1 I102_451(w_102_451, w_046_082);
  nand2 I102_458(w_102_458, w_093_225, w_031_049);
  or2  I102_462(w_102_462, w_000_619, w_059_612);
  or2  I102_476(w_102_476, w_068_224, w_074_342);
  and2 I102_479(w_102_479, w_083_189, w_034_031);
  nand2 I102_491(w_102_491, w_090_510, w_008_453);
  or2  I102_505(w_102_505, w_041_378, w_054_061);
  not1 I102_523(w_102_523, w_060_278);
  or2  I102_526(w_102_526, w_034_055, w_022_112);
  not1 I102_529(w_102_529, w_005_142);
  nand2 I102_542(w_102_542, w_016_007, w_076_300);
  nand2 I102_546(w_102_546, w_063_304, w_013_090);
  not1 I102_550(w_102_550, w_100_013);
  or2  I102_553(w_102_553, w_083_066, w_080_230);
  or2  I102_555(w_102_555, w_031_134, w_001_001);
  not1 I102_561(w_102_561, w_032_045);
  or2  I102_563(w_102_563, w_027_118, w_063_224);
  and2 I102_575(w_102_575, w_007_342, w_019_006);
  nand2 I102_589(w_102_589, w_015_436, w_082_115);
  or2  I102_597(w_102_597, w_042_198, w_045_267);
  and2 I102_601(w_102_601, w_052_046, w_034_040);
  nand2 I102_609(w_102_609, w_004_333, w_021_138);
  not1 I102_618(w_102_618, w_098_040);
  nand2 I102_619(w_102_619, w_000_154, w_054_081);
  or2  I102_646(w_102_646, w_071_029, w_002_150);
  nand2 I102_647(w_102_649, w_102_648, w_061_464);
  or2  I102_648(w_102_650, w_054_545, w_102_649);
  and2 I102_649(w_102_651, w_102_650, w_092_307);
  not1 I102_650(w_102_652, w_102_651);
  or2  I102_651(w_102_653, w_102_652, w_074_184);
  and2 I102_652(w_102_654, w_102_653, w_102_665);
  and2 I102_653(w_102_655, w_102_654, w_056_369);
  or2  I102_654(w_102_648, w_102_655, w_085_146);
  nand2 I102_655(w_102_660, w_102_659, w_033_235);
  not1 I102_656(w_102_661, w_102_660);
  or2  I102_657(w_102_662, w_044_691, w_102_661);
  and2 I102_658(w_102_663, w_102_662, w_100_080);
  not1 I102_659(w_102_659, w_102_654);
  and2 I102_660(w_102_665, w_051_298, w_102_663);
  not1 I102_661(w_102_668, w_102_667);
  not1 I102_662(w_102_669, w_102_668);
  not1 I102_663(w_102_670, w_102_669);
  not1 I102_664(w_102_671, w_102_670);
  or2  I102_665(w_102_672, w_102_690, w_102_671);
  or2  I102_666(w_102_673, w_102_672, w_044_458);
  or2  I102_667(w_102_674, w_102_673, w_045_199);
  nand2 I102_668(w_102_675, w_102_674, w_063_547);
  and2 I102_669(w_102_676, w_102_675, w_065_136);
  nand2 I102_670(w_102_667, w_102_676, w_040_101);
  not1 I102_671(w_102_681, w_102_680);
  and2 I102_672(w_102_682, w_072_232, w_102_681);
  and2 I102_673(w_102_683, w_040_404, w_102_682);
  not1 I102_674(w_102_684, w_102_683);
  nand2 I102_675(w_102_685, w_102_684, w_086_043);
  nand2 I102_676(w_102_686, w_012_118, w_102_685);
  or2  I102_677(w_102_687, w_021_022, w_102_686);
  and2 I102_678(w_102_688, w_038_340, w_102_687);
  not1 I102_679(w_102_680, w_102_672);
  and2 I102_680(w_102_690, w_049_003, w_102_688);
  or2  I103_002(w_103_002, w_076_258, w_010_255);
  or2  I103_006(w_103_006, w_053_014, w_045_332);
  and2 I103_007(w_103_007, w_053_028, w_070_408);
  or2  I103_015(w_103_015, w_022_247, w_082_123);
  or2  I103_016(w_103_016, w_052_009, w_035_083);
  nand2 I103_023(w_103_023, w_025_290, w_047_023);
  or2  I103_026(w_103_026, w_005_085, w_042_272);
  and2 I103_045(w_103_045, w_016_000, w_050_152);
  nand2 I103_048(w_103_048, w_092_377, w_003_062);
  or2  I103_053(w_103_053, w_040_583, w_084_034);
  nand2 I103_054(w_103_054, w_080_295, w_061_178);
  and2 I103_056(w_103_056, w_053_046, w_043_021);
  not1 I103_059(w_103_059, w_064_078);
  and2 I103_063(w_103_063, w_099_087, w_085_257);
  or2  I103_064(w_103_064, w_006_098, w_057_289);
  and2 I103_067(w_103_067, w_092_548, w_018_021);
  and2 I103_068(w_103_068, w_066_126, w_045_105);
  and2 I103_072(w_103_072, w_028_574, w_045_276);
  not1 I103_075(w_103_075, w_037_041);
  or2  I103_076(w_103_076, w_038_515, w_026_410);
  or2  I103_083(w_103_083, w_095_023, w_011_175);
  and2 I103_084(w_103_084, w_035_092, w_072_106);
  not1 I103_092(w_103_092, w_067_395);
  nand2 I103_098(w_103_098, w_000_412, w_025_297);
  and2 I103_105(w_103_105, w_073_347, w_052_025);
  and2 I103_108(w_103_108, w_029_075, w_061_058);
  not1 I103_113(w_103_113, w_027_027);
  and2 I103_114(w_103_114, w_002_297, w_064_289);
  or2  I103_117(w_103_117, w_047_021, w_036_140);
  nand2 I103_121(w_103_121, w_056_633, w_066_421);
  and2 I103_123(w_103_123, w_024_144, w_092_029);
  nand2 I103_128(w_103_128, w_069_265, w_080_238);
  or2  I103_136(w_103_136, w_098_019, w_080_237);
  and2 I103_137(w_103_137, w_029_002, w_092_011);
  not1 I103_140(w_103_140, w_077_519);
  or2  I103_143(w_103_143, w_066_319, w_022_023);
  nand2 I103_145(w_103_145, w_099_078, w_032_524);
  nand2 I103_147(w_103_147, w_074_100, w_040_254);
  and2 I103_149(w_103_149, w_005_148, w_004_138);
  not1 I103_156(w_103_156, w_041_441);
  and2 I103_162(w_103_162, w_012_178, w_050_135);
  nand2 I103_168(w_103_168, w_030_249, w_056_323);
  or2  I103_185(w_103_185, w_010_360, w_073_224);
  and2 I103_191(w_103_191, w_082_577, w_047_132);
  or2  I103_195(w_103_195, w_049_386, w_039_370);
  nand2 I103_199(w_103_199, w_081_020, w_068_342);
  or2  I103_206(w_103_206, w_015_095, w_031_165);
  and2 I103_210(w_103_210, w_034_039, w_012_013);
  and2 I103_213(w_103_213, w_027_081, w_088_126);
  not1 I103_220(w_103_220, w_035_007);
  not1 I103_228(w_103_228, w_090_088);
  nand2 I103_230(w_103_230, w_039_148, w_026_661);
  nand2 I103_232(w_103_232, w_072_090, w_026_006);
  not1 I103_240(w_103_240, w_012_345);
  and2 I103_248(w_103_248, w_069_053, w_093_321);
  and2 I103_260(w_103_260, w_033_513, w_078_063);
  nand2 I103_264(w_103_264, w_086_277, w_031_590);
  not1 I103_287(w_103_287, w_046_517);
  nand2 I103_289(w_103_289, w_067_382, w_055_259);
  nand2 I103_292(w_103_292, w_070_287, w_092_242);
  or2  I103_301(w_103_301, w_040_317, w_051_313);
  or2  I103_313(w_103_313, w_098_018, w_083_156);
  or2  I104_000(w_104_000, w_012_136, w_073_613);
  or2  I104_004(w_104_004, w_029_003, w_038_498);
  nand2 I104_007(w_104_007, w_094_587, w_001_031);
  not1 I104_009(w_104_009, w_059_026);
  not1 I104_021(w_104_021, w_103_098);
  nand2 I104_025(w_104_025, w_099_070, w_007_281);
  or2  I104_029(w_104_029, w_042_113, w_053_115);
  nand2 I104_033(w_104_033, w_012_078, w_006_020);
  not1 I104_040(w_104_040, w_034_061);
  or2  I104_042(w_104_042, w_010_073, w_029_072);
  and2 I104_047(w_104_047, w_079_029, w_003_065);
  and2 I104_053(w_104_053, w_083_066, w_072_107);
  and2 I104_057(w_104_057, w_059_001, w_048_008);
  nand2 I104_062(w_104_062, w_027_071, w_080_053);
  or2  I104_063(w_104_063, w_053_093, w_036_277);
  or2  I104_067(w_104_067, w_059_057, w_079_035);
  not1 I104_068(w_104_068, w_027_189);
  or2  I104_073(w_104_073, w_069_157, w_086_336);
  not1 I104_080(w_104_080, w_031_054);
  nand2 I104_091(w_104_091, w_010_563, w_025_158);
  nand2 I104_100(w_104_100, w_061_294, w_045_292);
  and2 I104_109(w_104_109, w_040_614, w_056_579);
  and2 I104_112(w_104_112, w_004_468, w_075_134);
  not1 I104_131(w_104_131, w_101_063);
  and2 I104_137(w_104_137, w_019_004, w_024_301);
  nand2 I104_138(w_104_138, w_072_043, w_005_160);
  not1 I104_143(w_104_143, w_087_249);
  or2  I104_144(w_104_144, w_087_118, w_037_063);
  nand2 I104_152(w_104_152, w_035_101, w_074_032);
  not1 I104_157(w_104_157, w_019_011);
  and2 I104_158(w_104_158, w_012_325, w_079_039);
  or2  I104_162(w_104_162, w_095_010, w_027_079);
  and2 I104_168(w_104_168, w_049_178, w_027_071);
  not1 I104_178(w_104_178, w_043_039);
  or2  I104_179(w_104_179, w_073_474, w_063_115);
  or2  I104_188(w_104_188, w_047_208, w_029_027);
  not1 I104_193(w_104_193, w_064_271);
  or2  I104_197(w_104_197, w_001_004, w_008_484);
  nand2 I104_199(w_104_199, w_047_051, w_009_087);
  or2  I104_213(w_104_213, w_070_096, w_063_198);
  and2 I104_216(w_104_216, w_020_500, w_061_182);
  not1 I104_221(w_104_221, w_051_147);
  nand2 I104_228(w_104_228, w_090_266, w_018_021);
  or2  I104_233(w_104_233, w_064_311, w_041_499);
  not1 I104_256(w_104_256, w_066_476);
  nand2 I104_260(w_104_260, w_054_549, w_078_381);
  and2 I104_263(w_104_263, w_073_569, w_079_037);
  and2 I104_264(w_104_264, w_004_175, w_024_139);
  or2  I104_266(w_104_266, w_068_250, w_025_105);
  and2 I104_271(w_104_271, w_082_393, w_032_095);
  not1 I104_273(w_104_273, w_063_244);
  or2  I104_278(w_104_278, w_016_005, w_021_175);
  nand2 I104_280(w_104_280, w_093_089, w_080_003);
  not1 I104_284(w_104_284, w_036_121);
  or2  I104_290(w_104_290, w_046_171, w_052_002);
  not1 I104_291(w_104_291, w_012_304);
  or2  I104_298(w_104_298, w_095_010, w_098_005);
  nand2 I104_299(w_104_299, w_043_039, w_056_438);
  or2  I104_310(w_104_310, w_024_065, w_058_478);
  nand2 I104_311(w_104_311, w_043_019, w_049_175);
  not1 I104_321(w_104_321, w_098_052);
  or2  I104_323(w_104_323, w_094_162, w_034_020);
  nand2 I104_326(w_104_326, w_078_416, w_019_011);
  not1 I104_335(w_104_335, w_045_272);
  or2  I104_342(w_104_342, w_016_003, w_058_251);
  not1 I104_354(w_104_354, w_024_127);
  and2 I104_357(w_104_357, w_058_056, w_001_035);
  and2 I104_362(w_104_362, w_044_371, w_003_083);
  nand2 I104_366(w_104_366, w_026_227, w_024_049);
  and2 I104_370(w_104_370, w_024_419, w_073_605);
  not1 I105_001(w_105_001, w_036_175);
  nand2 I105_005(w_105_005, w_015_322, w_090_122);
  not1 I105_016(w_105_016, w_057_022);
  and2 I105_029(w_105_029, w_004_059, w_035_099);
  not1 I105_045(w_105_045, w_091_063);
  nand2 I105_052(w_105_052, w_008_358, w_050_401);
  or2  I105_079(w_105_079, w_094_095, w_094_574);
  nand2 I105_082(w_105_082, w_082_082, w_028_127);
  or2  I105_088(w_105_088, w_099_148, w_089_055);
  or2  I105_091(w_105_091, w_044_197, w_009_510);
  and2 I105_093(w_105_093, w_016_003, w_013_562);
  not1 I105_097(w_105_097, w_005_012);
  nand2 I105_102(w_105_102, w_040_077, w_027_102);
  and2 I105_120(w_105_120, w_044_033, w_026_059);
  or2  I105_123(w_105_123, w_013_507, w_089_258);
  nand2 I105_129(w_105_129, w_063_072, w_102_097);
  and2 I105_130(w_105_130, w_087_227, w_000_379);
  or2  I105_132(w_105_132, w_072_097, w_100_109);
  nand2 I105_134(w_105_134, w_059_258, w_042_422);
  or2  I105_144(w_105_144, w_080_284, w_003_056);
  nand2 I105_163(w_105_163, w_104_109, w_077_029);
  and2 I105_169(w_105_169, w_041_053, w_083_061);
  or2  I105_182(w_105_182, w_097_570, w_092_059);
  not1 I105_192(w_105_192, w_000_592);
  or2  I105_198(w_105_198, w_030_061, w_054_114);
  not1 I105_199(w_105_199, w_031_049);
  nand2 I105_200(w_105_200, w_051_398, w_088_061);
  and2 I105_202(w_105_202, w_086_320, w_074_344);
  nand2 I105_211(w_105_211, w_058_498, w_056_214);
  nand2 I105_213(w_105_213, w_010_290, w_060_019);
  and2 I105_216(w_105_216, w_068_094, w_058_119);
  or2  I105_218(w_105_218, w_044_459, w_038_468);
  or2  I105_220(w_105_220, w_034_046, w_021_144);
  or2  I105_226(w_105_226, w_062_465, w_030_279);
  or2  I105_229(w_105_229, w_102_036, w_064_032);
  and2 I105_235(w_105_235, w_005_156, w_075_005);
  or2  I105_241(w_105_241, w_078_145, w_068_275);
  not1 I105_248(w_105_248, w_004_133);
  nand2 I105_249(w_105_249, w_043_018, w_070_185);
  and2 I105_251(w_105_251, w_009_343, w_056_129);
  not1 I105_253(w_105_253, w_026_092);
  and2 I105_264(w_105_264, w_076_014, w_035_019);
  or2  I105_265(w_105_265, w_009_159, w_083_033);
  not1 I105_267(w_105_267, w_016_006);
  nand2 I105_268(w_105_268, w_072_082, w_048_016);
  and2 I105_274(w_105_274, w_021_205, w_091_160);
  nand2 I105_282(w_105_282, w_002_035, w_047_277);
  and2 I105_284(w_105_284, w_069_001, w_044_296);
  and2 I105_294(w_105_294, w_102_526, w_054_184);
  not1 I105_305(w_105_305, w_074_252);
  nand2 I105_325(w_105_325, w_073_198, w_029_080);
  and2 I105_327(w_105_327, w_070_009, w_062_134);
  or2  I105_331(w_105_331, w_064_056, w_043_029);
  not1 I105_336(w_105_336, w_011_558);
  or2  I105_339(w_105_339, w_087_357, w_097_492);
  or2  I105_346(w_105_346, w_025_258, w_035_027);
  or2  I105_351(w_105_351, w_054_024, w_009_405);
  or2  I105_364(w_105_364, w_034_011, w_002_608);
  or2  I105_372(w_105_372, w_045_362, w_079_029);
  nand2 I105_384(w_105_384, w_095_014, w_060_155);
  not1 I105_386(w_105_386, w_092_595);
  and2 I105_388(w_105_388, w_094_542, w_097_033);
  nand2 I106_000(w_106_000, w_069_023, w_036_034);
  or2  I106_006(w_106_006, w_045_361, w_069_107);
  and2 I106_012(w_106_012, w_082_069, w_078_015);
  or2  I106_021(w_106_021, w_078_230, w_029_082);
  and2 I106_023(w_106_023, w_073_715, w_035_021);
  not1 I106_025(w_106_025, w_069_223);
  or2  I106_027(w_106_027, w_007_277, w_013_083);
  nand2 I106_032(w_106_032, w_050_406, w_060_208);
  and2 I106_037(w_106_037, w_084_007, w_056_709);
  and2 I106_043(w_106_043, w_014_188, w_047_275);
  not1 I106_044(w_106_044, w_032_521);
  nand2 I106_050(w_106_050, w_068_249, w_058_070);
  not1 I106_051(w_106_051, w_016_006);
  or2  I106_052(w_106_052, w_024_027, w_046_127);
  or2  I106_054(w_106_054, w_088_052, w_066_376);
  and2 I106_058(w_106_058, w_042_038, w_101_223);
  nand2 I106_062(w_106_062, w_052_001, w_081_006);
  not1 I106_065(w_106_065, w_044_532);
  or2  I106_066(w_106_066, w_045_231, w_051_330);
  and2 I106_067(w_106_067, w_023_026, w_078_573);
  not1 I106_069(w_106_069, w_004_274);
  or2  I106_072(w_106_072, w_061_042, w_051_103);
  nand2 I106_075(w_106_075, w_014_104, w_049_164);
  not1 I106_076(w_106_076, w_078_366);
  nand2 I106_081(w_106_081, w_092_673, w_057_213);
  not1 I106_083(w_106_083, w_020_034);
  not1 I106_084(w_106_084, w_059_708);
  not1 I106_089(w_106_089, w_048_006);
  or2  I106_091(w_106_091, w_040_682, w_057_070);
  not1 I106_093(w_106_093, w_051_025);
  nand2 I106_096(w_106_096, w_018_043, w_052_003);
  and2 I106_098(w_106_098, w_053_037, w_012_057);
  not1 I106_101(w_106_101, w_105_294);
  nand2 I106_105(w_106_105, w_040_571, w_043_008);
  and2 I106_107(w_106_107, w_046_174, w_024_371);
  or2  I106_108(w_106_108, w_097_480, w_096_001);
  or2  I106_116(w_106_116, w_091_119, w_044_675);
  not1 I106_123(w_106_123, w_066_118);
  nand2 I106_124(w_106_124, w_015_290, w_005_085);
  not1 I106_127(w_106_127, w_017_368);
  or2  I106_129(w_106_129, w_042_169, w_105_253);
  not1 I106_138(w_106_138, w_001_008);
  or2  I106_139(w_106_139, w_015_048, w_000_648);
  or2  I106_140(w_106_140, w_037_105, w_022_221);
  nand2 I106_141(w_106_141, w_044_588, w_074_127);
  and2 I106_144(w_106_144, w_032_025, w_006_222);
  and2 I106_146(w_106_146, w_063_197, w_039_609);
  or2  I106_147(w_106_147, w_074_200, w_031_277);
  not1 I106_160(w_106_160, w_018_043);
  nand2 I106_162(w_106_162, w_086_151, w_030_259);
  and2 I106_165(w_106_165, w_092_050, w_006_175);
  and2 I106_170(w_106_170, w_065_075, w_044_119);
  nand2 I106_181(w_106_181, w_017_102, w_016_001);
  nand2 I106_183(w_106_183, w_027_149, w_064_010);
  not1 I106_199(w_106_199, w_042_090);
  not1 I106_204(w_106_204, w_059_392);
  and2 I106_206(w_106_206, w_099_188, w_062_159);
  and2 I107_003(w_107_003, w_059_587, w_100_095);
  not1 I107_005(w_107_005, w_001_003);
  and2 I107_021(w_107_021, w_093_055, w_046_288);
  or2  I107_047(w_107_047, w_043_047, w_084_017);
  or2  I107_054(w_107_054, w_009_420, w_047_087);
  not1 I107_056(w_107_056, w_054_021);
  or2  I107_068(w_107_068, w_078_225, w_097_142);
  not1 I107_080(w_107_080, w_043_009);
  nand2 I107_082(w_107_082, w_039_543, w_000_006);
  and2 I107_091(w_107_091, w_022_153, w_087_219);
  not1 I107_094(w_107_094, w_034_030);
  nand2 I107_096(w_107_096, w_073_200, w_025_138);
  not1 I107_097(w_107_097, w_056_383);
  not1 I107_100(w_107_100, w_040_088);
  not1 I107_103(w_107_103, w_091_127);
  or2  I107_109(w_107_109, w_088_106, w_031_540);
  and2 I107_115(w_107_115, w_088_070, w_100_121);
  nand2 I107_118(w_107_118, w_069_199, w_047_317);
  and2 I107_121(w_107_121, w_078_318, w_076_046);
  nand2 I107_125(w_107_125, w_000_376, w_039_588);
  nand2 I107_126(w_107_126, w_034_036, w_039_527);
  nand2 I107_130(w_107_130, w_074_117, w_065_074);
  and2 I107_150(w_107_150, w_036_323, w_015_280);
  or2  I107_151(w_107_151, w_028_565, w_096_004);
  or2  I107_157(w_107_157, w_071_113, w_026_068);
  or2  I107_159(w_107_159, w_080_222, w_052_026);
  not1 I107_161(w_107_161, w_069_014);
  nand2 I107_177(w_107_177, w_073_258, w_032_579);
  or2  I107_180(w_107_180, w_045_344, w_068_237);
  or2  I107_181(w_107_181, w_083_088, w_077_586);
  nand2 I107_183(w_107_183, w_020_438, w_098_031);
  not1 I107_186(w_107_186, w_018_033);
  not1 I107_211(w_107_211, w_065_499);
  or2  I107_219(w_107_219, w_070_158, w_002_041);
  not1 I107_220(w_107_220, w_065_590);
  not1 I107_221(w_107_221, w_045_060);
  not1 I107_238(w_107_238, w_048_000);
  or2  I107_252(w_107_252, w_100_012, w_095_010);
  or2  I107_256(w_107_256, w_013_108, w_022_373);
  or2  I107_258(w_107_258, w_043_016, w_097_374);
  and2 I107_259(w_107_259, w_085_030, w_048_013);
  nand2 I107_272(w_107_272, w_099_025, w_033_008);
  or2  I107_279(w_107_279, w_104_100, w_101_209);
  or2  I107_288(w_107_288, w_102_523, w_078_038);
  not1 I107_292(w_107_292, w_015_223);
  and2 I107_293(w_107_293, w_082_139, w_065_389);
  and2 I107_302(w_107_302, w_051_150, w_022_334);
  nand2 I107_304(w_107_304, w_014_096, w_033_377);
  and2 I107_310(w_107_310, w_040_353, w_106_051);
  and2 I107_313(w_107_313, w_064_018, w_026_536);
  and2 I107_318(w_107_318, w_060_039, w_068_106);
  nand2 I107_329(w_107_329, w_019_017, w_105_134);
  or2  I107_345(w_107_345, w_016_007, w_049_210);
  and2 I107_349(w_107_349, w_083_071, w_067_390);
  and2 I107_355(w_107_355, w_102_115, w_034_003);
  and2 I107_370(w_107_370, w_049_337, w_072_195);
  and2 I107_379(w_107_379, w_064_265, w_031_148);
  not1 I107_396(w_107_396, w_106_091);
  not1 I107_400(w_107_400, w_083_052);
  not1 I107_415(w_107_415, w_031_541);
  and2 I107_425(w_107_425, w_082_526, w_005_014);
  or2  I108_000(w_108_000, w_044_338, w_038_022);
  or2  I108_001(w_108_001, w_050_035, w_039_377);
  and2 I108_002(w_108_002, w_004_061, w_094_449);
  nand2 I108_003(w_108_003, w_042_406, w_069_023);
  nand2 I108_006(w_108_006, w_011_240, w_098_010);
  or2  I108_015(w_108_015, w_103_313, w_094_386);
  and2 I108_021(w_108_021, w_054_133, w_098_042);
  not1 I108_024(w_108_024, w_019_013);
  or2  I108_026(w_108_026, w_033_534, w_090_061);
  or2  I108_031(w_108_031, w_013_526, w_037_206);
  or2  I108_035(w_108_035, w_082_019, w_103_117);
  nand2 I108_040(w_108_040, w_048_001, w_036_029);
  not1 I108_053(w_108_053, w_101_077);
  and2 I108_057(w_108_057, w_099_101, w_013_560);
  or2  I108_065(w_108_065, w_080_245, w_015_162);
  nand2 I108_067(w_108_067, w_039_093, w_054_186);
  and2 I108_073(w_108_073, w_040_133, w_105_211);
  and2 I108_078(w_108_078, w_102_250, w_028_228);
  and2 I108_085(w_108_085, w_092_307, w_077_577);
  not1 I108_086(w_108_086, w_038_032);
  nand2 I108_087(w_108_087, w_104_144, w_002_300);
  and2 I108_090(w_108_090, w_039_699, w_016_008);
  and2 I108_095(w_108_095, w_030_171, w_066_123);
  nand2 I108_097(w_108_097, w_019_006, w_003_064);
  nand2 I108_103(w_108_103, w_101_188, w_002_604);
  not1 I108_115(w_108_115, w_075_053);
  or2  I108_119(w_108_119, w_023_144, w_044_377);
  nand2 I108_122(w_108_122, w_042_255, w_027_051);
  or2  I108_127(w_108_127, w_100_094, w_041_243);
  or2  I108_130(w_108_130, w_077_551, w_019_005);
  nand2 I108_132(w_108_132, w_054_144, w_030_365);
  and2 I108_143(w_108_143, w_056_703, w_074_363);
  or2  I108_145(w_108_145, w_082_041, w_010_587);
  and2 I108_150(w_108_150, w_107_115, w_076_218);
  not1 I108_159(w_108_159, w_086_065);
  not1 I108_161(w_108_161, w_106_183);
  nand2 I108_166(w_108_166, w_081_013, w_009_351);
  nand2 I108_174(w_108_174, w_034_020, w_083_118);
  not1 I108_182(w_108_182, w_096_000);
  or2  I108_183(w_108_183, w_079_025, w_096_003);
  or2  I108_188(w_108_188, w_086_062, w_048_006);
  not1 I108_190(w_108_190, w_000_349);
  and2 I108_197(w_108_197, w_073_262, w_100_046);
  and2 I108_200(w_108_200, w_072_000, w_016_006);
  not1 I108_201(w_108_201, w_085_034);
  not1 I108_203(w_108_203, w_016_005);
  and2 I108_205(w_108_205, w_085_244, w_022_056);
  not1 I108_207(w_108_207, w_083_165);
  not1 I109_002(w_109_002, w_081_011);
  and2 I109_003(w_109_003, w_005_311, w_047_174);
  or2  I109_005(w_109_005, w_070_468, w_101_293);
  and2 I109_009(w_109_009, w_107_425, w_093_077);
  and2 I109_011(w_109_011, w_086_064, w_050_610);
  nand2 I109_028(w_109_028, w_019_015, w_042_116);
  or2  I109_053(w_109_053, w_045_378, w_089_150);
  and2 I109_054(w_109_054, w_019_009, w_034_006);
  or2  I109_068(w_109_068, w_031_494, w_098_013);
  and2 I109_100(w_109_100, w_051_005, w_046_171);
  not1 I109_104(w_109_104, w_059_165);
  not1 I109_114(w_109_114, w_069_064);
  and2 I109_124(w_109_124, w_093_413, w_031_605);
  not1 I109_127(w_109_127, w_035_078);
  nand2 I109_131(w_109_131, w_004_409, w_030_067);
  not1 I109_152(w_109_152, w_088_079);
  nand2 I109_169(w_109_169, w_000_500, w_073_326);
  not1 I109_177(w_109_177, w_008_250);
  or2  I109_199(w_109_199, w_107_118, w_062_099);
  nand2 I109_204(w_109_204, w_036_084, w_083_116);
  not1 I109_209(w_109_209, w_009_035);
  not1 I109_213(w_109_213, w_064_182);
  not1 I109_217(w_109_217, w_107_177);
  and2 I109_219(w_109_219, w_088_051, w_041_504);
  not1 I109_229(w_109_229, w_046_394);
  or2  I109_233(w_109_233, w_063_222, w_108_040);
  or2  I109_238(w_109_238, w_003_051, w_020_550);
  and2 I109_240(w_109_240, w_048_009, w_095_036);
  or2  I109_251(w_109_251, w_081_006, w_089_057);
  nand2 I109_252(w_109_252, w_086_265, w_032_328);
  and2 I109_259(w_109_259, w_034_021, w_048_005);
  or2  I109_264(w_109_264, w_033_427, w_082_228);
  and2 I109_279(w_109_279, w_083_168, w_096_004);
  nand2 I109_280(w_109_280, w_021_131, w_098_028);
  and2 I109_282(w_109_282, w_000_232, w_042_172);
  nand2 I109_284(w_109_284, w_073_422, w_076_162);
  not1 I109_285(w_109_285, w_039_104);
  or2  I109_291(w_109_291, w_052_035, w_108_026);
  or2  I109_293(w_109_293, w_100_044, w_073_026);
  nand2 I109_327(w_109_327, w_008_699, w_049_177);
  nand2 I109_331(w_109_331, w_082_336, w_052_018);
  not1 I109_350(w_109_350, w_025_004);
  nand2 I109_352(w_109_352, w_030_037, w_082_531);
  not1 I109_358(w_109_358, w_087_286);
  nand2 I109_363(w_109_363, w_045_102, w_012_224);
  nand2 I109_374(w_109_374, w_063_450, w_087_025);
  or2  I109_383(w_109_383, w_023_060, w_013_279);
  nand2 I109_385(w_109_385, w_033_207, w_062_661);
  or2  I109_392(w_109_392, w_034_017, w_065_593);
  not1 I109_394(w_109_394, w_070_143);
  and2 I109_407(w_109_407, w_067_213, w_094_462);
  nand2 I109_457(w_109_457, w_058_327, w_101_130);
  or2  I109_473(w_109_473, w_000_277, w_023_046);
  and2 I109_474(w_109_474, w_090_295, w_090_047);
  not1 I109_486(w_109_486, w_065_576);
  or2  I110_004(w_110_004, w_097_480, w_023_161);
  not1 I110_017(w_110_017, w_005_049);
  or2  I110_022(w_110_022, w_027_138, w_013_006);
  or2  I110_026(w_110_026, w_099_114, w_048_007);
  not1 I110_032(w_110_032, w_062_661);
  not1 I110_039(w_110_039, w_005_084);
  nand2 I110_041(w_110_041, w_093_073, w_101_066);
  or2  I110_042(w_110_042, w_004_241, w_050_091);
  not1 I110_047(w_110_047, w_097_039);
  or2  I110_064(w_110_064, w_048_011, w_049_049);
  and2 I110_075(w_110_075, w_096_005, w_097_514);
  nand2 I110_087(w_110_087, w_090_523, w_100_130);
  and2 I110_090(w_110_090, w_042_367, w_039_616);
  nand2 I110_092(w_110_092, w_044_180, w_051_340);
  or2  I110_117(w_110_117, w_021_215, w_074_215);
  and2 I110_124(w_110_124, w_074_014, w_068_260);
  and2 I110_125(w_110_125, w_046_480, w_108_150);
  or2  I110_132(w_110_132, w_022_331, w_032_152);
  or2  I110_135(w_110_135, w_019_007, w_071_176);
  or2  I110_139(w_110_139, w_054_431, w_039_143);
  nand2 I110_147(w_110_147, w_045_274, w_009_123);
  and2 I110_148(w_110_148, w_008_354, w_034_058);
  and2 I110_154(w_110_154, w_037_062, w_058_341);
  not1 I110_171(w_110_171, w_099_055);
  not1 I110_175(w_110_175, w_038_108);
  nand2 I110_187(w_110_187, w_062_089, w_058_541);
  nand2 I110_196(w_110_196, w_037_073, w_025_015);
  or2  I110_197(w_110_197, w_013_092, w_076_237);
  and2 I110_210(w_110_210, w_032_363, w_069_049);
  nand2 I110_237(w_110_237, w_004_343, w_069_049);
  and2 I110_239(w_110_239, w_071_173, w_108_182);
  nand2 I110_242(w_110_242, w_091_046, w_100_002);
  and2 I110_246(w_110_246, w_093_421, w_061_046);
  not1 I110_250(w_110_250, w_085_265);
  not1 I110_260(w_110_260, w_003_024);
  not1 I110_262(w_110_262, w_006_116);
  not1 I110_273(w_110_273, w_090_532);
  and2 I110_275(w_110_275, w_095_031, w_109_169);
  or2  I110_277(w_110_277, w_096_000, w_088_011);
  nand2 I110_279(w_110_279, w_039_175, w_018_003);
  and2 I110_282(w_110_282, w_030_349, w_017_375);
  or2  I110_289(w_110_289, w_087_230, w_091_176);
  nand2 I110_290(w_110_290, w_103_213, w_096_005);
  not1 I110_294(w_110_294, w_074_374);
  or2  I110_295(w_110_295, w_008_663, w_046_373);
  nand2 I110_304(w_110_304, w_088_051, w_045_026);
  nand2 I110_318(w_110_318, w_095_057, w_082_026);
  or2  I110_327(w_110_327, w_014_124, w_088_126);
  and2 I110_335(w_110_335, w_050_570, w_043_005);
  nand2 I110_352(w_110_352, w_030_172, w_013_571);
  and2 I110_358(w_110_358, w_063_090, w_063_445);
  not1 I110_362(w_110_362, w_108_115);
  nand2 I110_363(w_110_363, w_054_394, w_065_687);
  not1 I110_364(w_110_364, w_063_297);
  or2  I110_376(w_110_376, w_069_182, w_041_305);
  not1 I110_386(w_110_386, w_053_134);
  or2  I110_401(w_110_401, w_109_100, w_095_026);
  and2 I110_405(w_110_405, w_073_492, w_048_017);
  not1 I110_410(w_110_410, w_044_722);
  or2  I110_425(w_110_425, w_075_023, w_067_254);
  or2  I110_459(w_110_459, w_073_139, w_006_150);
  not1 I110_461(w_110_463, w_110_462);
  or2  I110_462(w_110_464, w_110_463, w_016_007);
  or2  I110_463(w_110_465, w_110_477, w_110_464);
  and2 I110_464(w_110_466, w_003_080, w_110_465);
  and2 I110_465(w_110_462, w_110_466, w_091_166);
  or2  I110_466(w_110_471, w_110_470, w_099_257);
  nand2 I110_467(w_110_472, w_007_357, w_110_471);
  and2 I110_468(w_110_473, w_110_472, w_102_491);
  not1 I110_469(w_110_474, w_110_473);
  and2 I110_470(w_110_475, w_110_474, w_086_197);
  not1 I110_471(w_110_470, w_110_465);
  and2 I110_472(w_110_477, w_010_338, w_110_475);
  not1 I111_003(w_111_003, w_025_054);
  not1 I111_007(w_111_007, w_103_240);
  not1 I111_008(w_111_008, w_103_083);
  nand2 I111_010(w_111_010, w_000_096, w_087_366);
  not1 I111_011(w_111_011, w_030_352);
  not1 I111_012(w_111_012, w_016_001);
  not1 I111_018(w_111_018, w_010_721);
  and2 I111_019(w_111_019, w_078_122, w_082_244);
  and2 I111_020(w_111_020, w_049_335, w_056_554);
  nand2 I111_021(w_111_021, w_060_294, w_049_022);
  nand2 I111_023(w_111_023, w_034_027, w_087_333);
  not1 I111_027(w_111_027, w_039_082);
  or2  I111_034(w_111_034, w_067_326, w_068_181);
  and2 I111_039(w_111_039, w_063_047, w_090_370);
  nand2 I111_041(w_111_041, w_028_226, w_045_258);
  not1 I111_046(w_111_046, w_034_054);
  nand2 I111_047(w_111_047, w_071_171, w_078_168);
  nand2 I111_049(w_111_049, w_039_256, w_007_443);
  nand2 I111_054(w_111_054, w_033_149, w_073_044);
  or2  I111_059(w_111_059, w_088_067, w_081_013);
  and2 I111_061(w_111_061, w_023_063, w_054_109);
  nand2 I111_062(w_111_062, w_079_029, w_092_190);
  or2  I111_070(w_111_070, w_008_124, w_025_095);
  nand2 I111_078(w_111_078, w_025_288, w_078_152);
  not1 I111_081(w_111_081, w_000_102);
  nand2 I111_091(w_111_091, w_087_343, w_016_002);
  not1 I111_099(w_111_099, w_001_011);
  or2  I111_102(w_111_102, w_083_155, w_094_475);
  or2  I111_106(w_111_106, w_043_036, w_083_022);
  and2 I111_111(w_110_468, w_095_033, w_110_462);
  not1 I112_000(w_112_000, w_017_625);
  and2 I112_006(w_112_006, w_028_052, w_011_320);
  nand2 I112_008(w_112_008, w_042_260, w_051_027);
  or2  I112_010(w_112_010, w_104_335, w_041_485);
  nand2 I112_018(w_112_018, w_086_321, w_085_220);
  not1 I112_019(w_112_019, w_019_003);
  nand2 I112_021(w_112_021, w_013_340, w_075_071);
  not1 I112_022(w_112_022, w_042_257);
  or2  I112_025(w_112_025, w_052_028, w_006_228);
  or2  I112_035(w_112_035, w_004_411, w_035_035);
  not1 I112_039(w_112_039, w_069_063);
  and2 I112_046(w_112_046, w_064_036, w_097_335);
  or2  I112_054(w_112_054, w_030_146, w_017_662);
  not1 I112_056(w_112_056, w_077_289);
  or2  I112_063(w_112_063, w_033_019, w_098_048);
  and2 I112_065(w_112_065, w_092_562, w_025_067);
  and2 I112_068(w_112_068, w_110_468, w_008_686);
  not1 I112_077(w_112_077, w_083_191);
  and2 I112_078(w_112_078, w_049_372, w_095_004);
  not1 I112_079(w_112_079, w_061_002);
  or2  I112_084(w_112_084, w_053_158, w_003_015);
  nand2 I112_085(w_112_085, w_023_141, w_104_299);
  or2  I112_095(w_112_095, w_069_087, w_048_018);
  or2  I112_104(w_112_104, w_097_048, w_021_240);
  or2  I112_107(w_112_107, w_076_040, w_051_106);
  or2  I112_120(w_112_120, w_085_125, w_067_053);
  and2 I112_121(w_112_121, w_069_188, w_021_093);
  nand2 I112_127(w_112_127, w_016_001, w_067_053);
  not1 I112_130(w_112_130, w_028_123);
  nand2 I112_131(w_112_131, w_002_580, w_006_091);
  and2 I112_134(w_112_134, w_064_066, w_051_262);
  or2  I112_140(w_112_140, w_051_319, w_050_365);
  nand2 I112_143(w_112_143, w_009_517, w_091_134);
  nand2 I112_144(w_112_144, w_042_001, w_093_043);
  not1 I112_145(w_112_145, w_054_486);
  or2  I112_160(w_112_160, w_101_158, w_102_246);
  not1 I112_161(w_112_161, w_073_687);
  nand2 I112_165(w_112_165, w_045_050, w_108_201);
  nand2 I112_169(w_112_169, w_017_234, w_047_225);
  or2  I112_172(w_112_172, w_105_336, w_018_018);
  and2 I112_173(w_112_173, w_091_075, w_102_097);
  nand2 I112_174(w_112_174, w_041_670, w_002_050);
  or2  I112_180(w_112_180, w_059_508, w_076_292);
  nand2 I112_182(w_112_182, w_010_240, w_087_086);
  nand2 I112_187(w_112_187, w_099_044, w_058_368);
  or2  I112_189(w_112_189, w_078_084, w_056_084);
  and2 I112_197(w_112_197, w_019_001, w_109_252);
  and2 I113_008(w_113_008, w_090_384, w_046_073);
  nand2 I113_010(w_113_010, w_056_035, w_107_211);
  not1 I113_015(w_113_015, w_094_607);
  nand2 I113_019(w_113_019, w_013_346, w_010_147);
  or2  I113_025(w_113_025, w_109_124, w_072_020);
  nand2 I113_029(w_113_029, w_029_074, w_045_330);
  not1 I113_031(w_113_031, w_110_363);
  nand2 I113_032(w_113_032, w_061_198, w_042_359);
  not1 I113_033(w_113_033, w_093_252);
  nand2 I113_034(w_113_034, w_060_344, w_009_443);
  and2 I113_047(w_113_047, w_047_141, w_051_349);
  or2  I113_048(w_113_048, w_063_251, w_063_198);
  not1 I113_049(w_113_049, w_014_250);
  and2 I113_050(w_113_050, w_041_510, w_109_394);
  not1 I113_061(w_113_061, w_026_433);
  not1 I113_062(w_113_062, w_010_711);
  nand2 I113_081(w_113_081, w_043_046, w_025_036);
  nand2 I113_090(w_113_090, w_081_011, w_065_507);
  or2  I113_106(w_113_106, w_038_005, w_032_325);
  or2  I113_107(w_113_107, w_039_571, w_065_285);
  or2  I113_109(w_113_109, w_094_043, w_008_489);
  or2  I113_110(w_113_110, w_053_086, w_021_088);
  not1 I113_112(w_113_112, w_056_586);
  nand2 I113_114(w_113_114, w_017_103, w_070_496);
  or2  I113_120(w_113_120, w_094_079, w_005_027);
  and2 I113_125(w_113_125, w_078_169, w_106_147);
  or2  I113_132(w_113_132, w_101_214, w_074_351);
  not1 I113_136(w_113_136, w_020_500);
  not1 I113_146(w_113_146, w_010_002);
  and2 I113_154(w_113_154, w_051_309, w_044_569);
  or2  I113_158(w_113_158, w_079_012, w_063_085);
  nand2 I113_171(w_113_171, w_048_000, w_110_004);
  nand2 I113_172(w_113_172, w_096_000, w_062_273);
  not1 I113_174(w_113_174, w_058_570);
  or2  I113_181(w_113_181, w_107_186, w_096_003);
  or2  I113_185(w_113_185, w_043_045, w_067_329);
  and2 I113_187(w_113_187, w_021_237, w_050_007);
  not1 I113_188(w_113_188, w_025_010);
  or2  I113_198(w_113_198, w_040_524, w_105_388);
  or2  I113_209(w_113_209, w_036_146, w_032_019);
  nand2 I113_211(w_113_211, w_064_135, w_097_122);
  and2 I113_218(w_113_218, w_079_048, w_053_078);
  and2 I113_219(w_113_219, w_052_038, w_046_168);
  and2 I113_227(w_113_227, w_025_164, w_059_056);
  nand2 I113_231(w_113_231, w_061_196, w_069_167);
  not1 I113_234(w_113_234, w_034_064);
  or2  I113_237(w_113_237, w_012_103, w_010_205);
  nand2 I113_238(w_113_238, w_036_200, w_093_389);
  and2 I113_250(w_113_250, w_087_125, w_018_043);
  and2 I113_258(w_113_258, w_018_005, w_027_163);
  nand2 I113_262(w_113_262, w_054_274, w_038_169);
  and2 I113_267(w_113_267, w_026_250, w_057_025);
  or2  I113_269(w_113_269, w_091_094, w_094_421);
  not1 I113_273(w_113_273, w_067_005);
  not1 I113_276(w_113_276, w_048_002);
  or2  I113_289(w_113_289, w_034_033, w_052_025);
  and2 I113_291(w_113_291, w_104_298, w_057_032);
  or2  I113_300(w_113_300, w_109_005, w_023_124);
  not1 I113_309(w_113_309, w_100_038);
  not1 I113_316(w_113_316, w_076_364);
  not1 I113_318(w_113_318, w_058_104);
  or2  I113_323(w_113_323, w_006_168, w_030_241);
  and2 I113_341(w_113_341, w_033_091, w_061_192);
  or2  I113_347(w_113_347, w_064_166, w_049_373);
  nand2 I113_348(w_113_348, w_102_226, w_072_024);
  nand2 I114_003(w_114_003, w_020_547, w_033_132);
  or2  I114_007(w_114_007, w_029_041, w_055_164);
  nand2 I114_009(w_114_009, w_059_432, w_071_144);
  nand2 I114_015(w_114_015, w_023_027, w_081_000);
  and2 I114_018(w_114_018, w_006_142, w_032_025);
  or2  I114_020(w_114_020, w_113_112, w_099_223);
  nand2 I114_032(w_114_032, w_066_064, w_066_240);
  nand2 I114_036(w_114_036, w_044_589, w_011_093);
  nand2 I114_037(w_114_037, w_105_202, w_029_020);
  not1 I114_039(w_114_039, w_068_080);
  and2 I114_047(w_114_047, w_053_047, w_049_386);
  nand2 I114_056(w_114_056, w_065_144, w_053_058);
  not1 I114_058(w_114_058, w_062_229);
  not1 I114_065(w_114_065, w_038_076);
  or2  I114_067(w_114_067, w_031_467, w_037_132);
  nand2 I114_068(w_114_068, w_102_646, w_050_032);
  and2 I114_069(w_114_069, w_063_268, w_002_217);
  or2  I114_106(w_114_106, w_069_141, w_009_485);
  nand2 I114_112(w_114_112, w_017_592, w_076_137);
  and2 I114_114(w_114_114, w_001_035, w_044_710);
  or2  I114_116(w_114_116, w_047_115, w_018_004);
  nand2 I114_117(w_114_117, w_107_272, w_108_078);
  nand2 I114_118(w_114_118, w_066_135, w_044_080);
  nand2 I114_119(w_114_119, w_006_217, w_030_370);
  nand2 I114_120(w_114_120, w_104_143, w_103_195);
  not1 I114_131(w_114_131, w_092_209);
  nand2 I114_134(w_114_134, w_014_007, w_045_266);
  not1 I114_135(w_114_135, w_074_045);
  not1 I114_138(w_114_138, w_018_006);
  and2 I114_141(w_114_141, w_061_301, w_015_651);
  not1 I114_144(w_114_144, w_031_131);
  not1 I114_148(w_114_148, w_021_015);
  or2  I114_150(w_114_150, w_048_010, w_045_215);
  not1 I114_152(w_114_152, w_036_134);
  nand2 I114_167(w_114_167, w_074_331, w_009_351);
  and2 I114_170(w_114_170, w_009_406, w_019_000);
  or2  I114_176(w_114_176, w_053_075, w_107_370);
  or2  I114_181(w_114_181, w_066_293, w_102_282);
  nand2 I114_186(w_114_186, w_046_092, w_112_131);
  and2 I114_188(w_114_188, w_104_025, w_053_112);
  or2  I114_189(w_114_189, w_025_143, w_029_027);
  nand2 I114_194(w_114_194, w_069_039, w_029_088);
  or2  I114_195(w_114_195, w_019_009, w_070_505);
  and2 I114_197(w_114_197, w_103_084, w_005_268);
  or2  I114_198(w_114_198, w_066_349, w_087_310);
  not1 I114_209(w_114_209, w_112_144);
  nand2 I114_211(w_114_211, w_061_172, w_041_070);
  nand2 I114_217(w_114_217, w_020_179, w_102_553);
  or2  I114_220(w_114_220, w_092_478, w_106_043);
  and2 I114_226(w_114_226, w_101_085, w_014_047);
  or2  I115_000(w_115_000, w_071_322, w_023_191);
  not1 I115_004(w_115_004, w_031_425);
  nand2 I115_005(w_115_005, w_036_010, w_036_314);
  nand2 I115_008(w_115_008, w_106_162, w_023_208);
  nand2 I115_016(w_115_016, w_007_413, w_014_140);
  nand2 I115_018(w_115_018, w_113_291, w_015_278);
  nand2 I115_019(w_115_019, w_098_032, w_065_280);
  nand2 I115_021(w_115_021, w_018_044, w_028_165);
  not1 I115_033(w_115_033, w_080_249);
  or2  I115_036(w_115_036, w_002_004, w_053_056);
  not1 I115_037(w_115_037, w_045_290);
  or2  I115_039(w_115_039, w_003_052, w_071_100);
  not1 I115_040(w_115_040, w_036_224);
  and2 I115_055(w_115_055, w_033_053, w_024_020);
  not1 I115_061(w_115_061, w_018_024);
  not1 I115_065(w_115_065, w_034_059);
  and2 I115_066(w_115_066, w_013_556, w_113_110);
  nand2 I115_075(w_115_075, w_001_008, w_051_203);
  nand2 I115_084(w_115_084, w_060_088, w_001_001);
  and2 I115_089(w_115_089, w_015_343, w_036_182);
  or2  I115_101(w_115_101, w_052_037, w_029_017);
  not1 I115_122(w_115_122, w_009_090);
  or2  I115_125(w_115_125, w_114_217, w_099_291);
  not1 I115_126(w_115_126, w_089_213);
  or2  I115_131(w_115_131, w_047_126, w_028_209);
  not1 I115_134(w_115_134, w_103_045);
  or2  I115_135(w_115_135, w_004_106, w_032_133);
  or2  I115_136(w_115_136, w_010_458, w_111_019);
  not1 I115_151(w_115_151, w_041_342);
  and2 I115_152(w_115_152, w_030_036, w_105_005);
  and2 I115_162(w_115_162, w_044_229, w_067_343);
  nand2 I115_169(w_115_169, w_096_001, w_108_035);
  not1 I115_178(w_115_178, w_087_326);
  nand2 I115_179(w_115_179, w_113_185, w_082_551);
  not1 I115_190(w_115_190, w_106_027);
  or2  I115_191(w_115_191, w_025_189, w_102_152);
  nand2 I115_194(w_115_194, w_083_013, w_030_280);
  nand2 I115_209(w_115_209, w_070_027, w_112_046);
  and2 I115_215(w_115_215, w_029_013, w_070_161);
  not1 I115_219(w_115_219, w_033_109);
  not1 I115_228(w_115_228, w_063_072);
  or2  I115_240(w_115_240, w_110_187, w_007_343);
  not1 I115_241(w_115_241, w_032_514);
  nand2 I115_251(w_115_251, w_021_123, w_025_055);
  and2 I116_001(w_116_001, w_074_107, w_009_104);
  not1 I116_004(w_116_004, w_097_070);
  not1 I116_008(w_116_008, w_009_114);
  and2 I116_023(w_116_023, w_011_080, w_075_049);
  and2 I116_030(w_116_030, w_021_205, w_028_541);
  nand2 I116_042(w_116_042, w_055_298, w_021_079);
  not1 I116_061(w_116_061, w_058_425);
  nand2 I116_077(w_116_077, w_096_001, w_113_238);
  or2  I116_079(w_116_079, w_102_308, w_001_004);
  not1 I116_092(w_116_092, w_113_125);
  and2 I116_112(w_116_112, w_045_282, w_047_088);
  and2 I116_118(w_116_118, w_022_150, w_003_022);
  or2  I116_122(w_116_122, w_018_044, w_034_049);
  and2 I116_124(w_116_124, w_058_527, w_104_152);
  and2 I116_126(w_116_126, w_010_343, w_079_022);
  not1 I116_136(w_116_136, w_034_018);
  or2  I116_140(w_116_140, w_071_213, w_066_341);
  nand2 I116_142(w_116_142, w_115_005, w_043_037);
  not1 I116_150(w_116_150, w_047_148);
  and2 I116_153(w_116_153, w_013_419, w_051_200);
  nand2 I116_192(w_116_192, w_030_243, w_046_616);
  or2  I116_204(w_116_204, w_045_048, w_096_003);
  or2  I116_224(w_116_224, w_043_001, w_104_137);
  nand2 I116_231(w_116_231, w_085_088, w_012_032);
  not1 I116_238(w_116_238, w_092_068);
  and2 I116_260(w_116_260, w_064_069, w_009_501);
  not1 I116_261(w_116_261, w_096_000);
  and2 I116_287(w_116_287, w_011_260, w_079_002);
  nand2 I116_292(w_116_292, w_067_358, w_038_178);
  and2 I116_343(w_116_343, w_063_120, w_050_602);
  and2 I116_345(w_116_345, w_071_217, w_018_013);
  and2 I116_348(w_116_348, w_072_067, w_100_056);
  nand2 I116_365(w_116_365, w_073_722, w_084_033);
  nand2 I116_373(w_116_373, w_055_226, w_093_084);
  and2 I116_387(w_116_387, w_105_305, w_015_271);
  not1 I116_407(w_116_407, w_009_399);
  not1 I116_412(w_116_412, w_089_013);
  or2  I116_414(w_116_414, w_044_418, w_030_225);
  not1 I116_420(w_116_420, w_088_043);
  or2  I116_424(w_116_424, w_084_028, w_030_057);
  and2 I116_426(w_116_426, w_031_319, w_042_147);
  nand2 I116_428(w_116_428, w_034_072, w_110_290);
  not1 I116_495(w_116_495, w_071_124);
  or2  I116_497(w_116_497, w_086_208, w_055_033);
  and2 I116_500(w_116_500, w_046_336, w_047_142);
  and2 I116_510(w_116_510, w_088_094, w_031_009);
  and2 I116_513(w_116_513, w_012_109, w_003_061);
  not1 I116_530(w_116_530, w_030_167);
  not1 I116_532(w_116_532, w_069_025);
  nand2 I116_545(w_116_545, w_078_401, w_107_126);
  not1 I116_554(w_116_554, w_059_425);
  or2  I116_570(w_116_570, w_094_167, w_040_386);
  nand2 I116_576(w_116_576, w_070_175, w_104_063);
  or2  I116_601(w_116_601, w_010_045, w_064_174);
  and2 I116_628(w_116_628, w_078_396, w_034_039);
  or2  I116_636(w_116_636, w_075_061, w_061_240);
  not1 I116_638(w_116_640, w_116_639);
  or2  I116_639(w_116_641, w_089_026, w_116_640);
  and2 I116_640(w_116_642, w_015_005, w_116_641);
  or2  I116_641(w_116_643, w_116_642, w_105_129);
  nand2 I116_642(w_116_644, w_115_219, w_116_643);
  not1 I116_643(w_116_645, w_116_644);
  and2 I116_644(w_116_646, w_116_645, w_115_191);
  nand2 I116_645(w_116_647, w_116_646, w_042_008);
  and2 I116_646(w_116_648, w_066_315, w_116_647);
  and2 I116_647(w_116_649, w_116_648, w_057_141);
  and2 I116_648(w_116_639, w_007_327, w_116_649);
  or2  I117_000(w_117_000, w_058_195, w_025_174);
  or2  I117_004(w_117_004, w_032_264, w_013_055);
  and2 I117_005(w_117_005, w_103_105, w_115_004);
  nand2 I117_008(w_117_008, w_027_159, w_015_477);
  or2  I117_010(w_117_010, w_025_000, w_012_005);
  nand2 I117_011(w_117_011, w_095_036, w_069_128);
  nand2 I117_012(w_117_012, w_100_010, w_064_097);
  not1 I117_014(w_117_014, w_112_021);
  and2 I117_016(w_117_016, w_048_005, w_071_047);
  not1 I117_017(w_117_017, w_096_004);
  and2 I117_018(w_117_018, w_006_085, w_009_024);
  nand2 I117_020(w_117_020, w_060_209, w_078_037);
  and2 I117_022(w_117_022, w_085_199, w_040_509);
  or2  I117_024(w_117_024, w_028_267, w_096_000);
  or2  I117_026(w_117_026, w_061_064, w_035_000);
  nand2 I117_028(w_117_028, w_098_071, w_102_491);
  and2 I117_029(w_117_029, w_080_311, w_093_224);
  nand2 I117_033(w_117_033, w_089_026, w_113_090);
  nand2 I117_035(w_117_035, w_064_036, w_083_182);
  and2 I117_036(w_117_036, w_035_050, w_046_033);
  not1 I117_038(w_117_038, w_075_032);
  and2 I117_040(w_117_040, w_041_446, w_025_130);
  and2 I117_043(w_117_043, w_084_018, w_089_106);
  nand2 I117_045(w_117_045, w_108_006, w_083_018);
  not1 I117_046(w_117_046, w_084_034);
  or2  I117_048(w_117_048, w_067_292, w_064_338);
  nand2 I117_050(w_117_050, w_058_447, w_031_100);
  nand2 I117_051(w_117_051, w_096_001, w_042_206);
  nand2 I117_053(w_117_053, w_037_130, w_085_150);
  not1 I117_054(w_117_054, w_077_424);
  and2 I117_055(w_117_055, w_050_041, w_038_142);
  nand2 I117_056(w_117_056, w_005_134, w_059_522);
  nand2 I117_057(w_117_057, w_107_096, w_017_538);
  or2  I117_058(w_117_058, w_102_505, w_043_037);
  nand2 I117_059(w_117_059, w_055_330, w_085_350);
  and2 I117_060(w_117_060, w_053_054, w_050_112);
  not1 I117_062(w_117_062, w_053_031);
  not1 I117_063(w_117_063, w_113_106);
  or2  I117_064(w_117_064, w_092_628, w_039_708);
  or2  I117_066(w_117_066, w_002_196, w_039_528);
  not1 I117_072(w_117_072, w_053_126);
  and2 I117_074(w_117_074, w_102_458, w_028_122);
  nand2 I117_075(w_117_075, w_047_294, w_064_194);
  or2  I117_078(w_117_078, w_020_287, w_009_465);
  and2 I117_079(w_117_079, w_115_228, w_106_140);
  or2  I117_088(w_117_088, w_075_024, w_074_190);
  or2  I118_000(w_118_000, w_060_330, w_077_086);
  or2  I118_005(w_118_005, w_041_349, w_018_002);
  or2  I118_010(w_118_010, w_026_025, w_088_012);
  and2 I118_012(w_118_012, w_040_356, w_106_083);
  nand2 I118_017(w_118_017, w_063_035, w_021_152);
  and2 I118_018(w_118_018, w_084_047, w_064_070);
  nand2 I118_019(w_118_019, w_108_130, w_065_132);
  and2 I118_023(w_118_023, w_064_118, w_075_136);
  nand2 I118_029(w_118_029, w_096_001, w_008_122);
  and2 I118_030(w_118_030, w_076_241, w_005_095);
  nand2 I118_031(w_118_031, w_106_021, w_011_533);
  and2 I118_036(w_118_036, w_032_183, w_098_001);
  nand2 I118_040(w_118_040, w_117_033, w_054_190);
  or2  I118_041(w_118_041, w_104_007, w_056_645);
  and2 I118_043(w_118_043, w_015_547, w_116_428);
  nand2 I118_050(w_118_050, w_014_285, w_051_398);
  nand2 I118_054(w_118_054, w_094_419, w_020_550);
  not1 I118_060(w_118_060, w_116_287);
  not1 I118_061(w_118_061, w_023_171);
  or2  I118_062(w_118_062, w_015_418, w_040_281);
  not1 I118_067(w_118_067, w_008_018);
  not1 I118_070(w_118_070, w_038_255);
  and2 I118_071(w_118_071, w_048_000, w_070_488);
  or2  I118_079(w_118_079, w_035_045, w_005_102);
  nand2 I118_080(w_118_080, w_088_090, w_067_224);
  and2 I118_081(w_118_081, w_035_078, w_032_021);
  or2  I118_082(w_118_082, w_091_164, w_067_276);
  or2  I118_087(w_118_087, w_058_485, w_047_362);
  nand2 I118_090(w_118_090, w_067_292, w_076_351);
  not1 I118_093(w_118_093, w_022_170);
  and2 I118_094(w_118_094, w_080_171, w_009_556);
  not1 I118_099(w_118_099, w_093_101);
  not1 I118_101(w_118_101, w_076_233);
  not1 I118_104(w_118_104, w_031_021);
  nand2 I118_106(w_118_108, w_118_107, w_118_132);
  and2 I118_107(w_118_109, w_118_108, w_038_600);
  not1 I118_108(w_118_110, w_118_109);
  or2  I118_109(w_118_111, w_118_110, w_062_673);
  or2  I118_110(w_118_112, w_028_405, w_118_111);
  and2 I118_111(w_118_113, w_118_112, w_005_185);
  and2 I118_112(w_118_114, w_118_113, w_118_134);
  or2  I118_113(w_118_115, w_118_114, w_111_020);
  or2  I118_114(w_118_116, w_118_115, w_062_628);
  or2  I118_115(w_118_117, w_059_596, w_118_116);
  and2 I118_116(w_118_118, w_002_080, w_118_117);
  nand2 I118_117(w_118_107, w_104_228, w_118_118);
  nand2 I118_118(w_118_123, w_017_515, w_118_122);
  nand2 I118_119(w_118_124, w_103_185, w_118_123);
  and2 I118_120(w_118_125, w_118_124, w_114_167);
  or2  I118_121(w_118_126, w_114_068, w_118_125);
  not1 I118_122(w_118_127, w_118_126);
  and2 I118_123(w_118_128, w_118_127, w_016_004);
  or2  I118_124(w_118_129, w_118_128, w_099_077);
  and2 I118_125(w_118_130, w_118_129, w_049_019);
  not1 I118_126(w_118_122, w_118_108);
  and2 I118_127(w_118_132, w_067_199, w_118_130);
  not1 I118_128(w_118_134, w_016_004);
  and2 I119_001(w_119_001, w_077_133, w_029_063);
  and2 I119_003(w_119_003, w_105_169, w_116_204);
  nand2 I119_007(w_119_007, w_011_013, w_075_118);
  or2  I119_012(w_119_012, w_091_067, w_059_114);
  or2  I119_014(w_119_014, w_083_036, w_012_242);
  and2 I119_016(w_119_016, w_103_092, w_039_063);
  and2 I119_017(w_119_017, w_047_318, w_030_137);
  or2  I119_018(w_119_018, w_015_343, w_018_035);
  not1 I119_027(w_119_027, w_045_283);
  nand2 I119_029(w_119_029, w_012_337, w_013_100);
  not1 I119_040(w_119_040, w_096_002);
  nand2 I119_043(w_119_043, w_044_405, w_075_069);
  nand2 I119_050(w_119_050, w_006_199, w_086_232);
  or2  I119_053(w_119_053, w_106_105, w_035_030);
  not1 I119_063(w_119_063, w_040_021);
  nand2 I119_067(w_119_067, w_047_139, w_060_265);
  or2  I119_070(w_119_070, w_002_002, w_048_009);
  not1 I119_082(w_119_082, w_063_104);
  nand2 I119_083(w_119_083, w_032_152, w_118_029);
  not1 I119_085(w_119_085, w_089_051);
  not1 I119_086(w_119_086, w_113_219);
  not1 I119_087(w_119_087, w_081_009);
  and2 I119_099(w_119_099, w_045_186, w_000_648);
  nand2 I119_101(w_119_101, w_031_271, w_069_042);
  and2 I119_103(w_119_103, w_040_469, w_064_197);
  not1 I119_104(w_119_104, w_041_337);
  nand2 I119_106(w_119_106, w_091_091, w_117_056);
  not1 I119_109(w_119_109, w_085_305);
  and2 I119_117(w_119_117, w_082_193, w_083_019);
  not1 I119_119(w_119_119, w_000_085);
  or2  I119_123(w_119_123, w_108_090, w_046_023);
  and2 I119_125(w_119_125, w_083_068, w_064_077);
  not1 I119_135(w_119_135, w_043_006);
  or2  I119_139(w_119_139, w_062_058, w_100_049);
  or2  I119_142(w_119_142, w_118_040, w_114_118);
  and2 I119_143(w_119_143, w_092_504, w_059_220);
  and2 I119_146(w_119_146, w_080_134, w_107_259);
  not1 I119_149(w_119_149, w_046_270);
  or2  I119_156(w_119_156, w_082_049, w_062_511);
  or2  I119_157(w_119_157, w_039_553, w_071_315);
  or2  I119_162(w_119_162, w_006_184, w_101_269);
  and2 I119_164(w_119_164, w_074_157, w_089_178);
  or2  I119_165(w_119_165, w_042_112, w_016_000);
  not1 I119_171(w_119_171, w_014_056);
  nand2 I119_175(w_119_175, w_071_045, w_012_269);
  and2 I119_177(w_119_177, w_039_432, w_067_374);
  and2 I119_188(w_119_188, w_096_004, w_076_158);
  nand2 I119_189(w_119_189, w_006_102, w_011_016);
  and2 I120_008(w_120_008, w_021_167, w_112_161);
  or2  I120_029(w_120_029, w_099_111, w_028_064);
  nand2 I120_038(w_120_038, w_017_238, w_060_224);
  not1 I120_042(w_120_042, w_098_062);
  or2  I120_051(w_120_051, w_021_128, w_061_194);
  not1 I120_060(w_120_060, w_050_105);
  and2 I120_072(w_120_072, w_030_031, w_013_176);
  or2  I120_083(w_120_083, w_027_047, w_109_199);
  not1 I120_104(w_120_104, w_036_170);
  nand2 I120_126(w_120_126, w_109_282, w_113_048);
  not1 I120_135(w_120_135, w_102_076);
  and2 I120_140(w_120_140, w_019_004, w_104_004);
  nand2 I120_159(w_120_159, w_076_345, w_042_427);
  not1 I120_167(w_120_167, w_004_315);
  and2 I120_169(w_120_169, w_109_252, w_048_010);
  not1 I120_176(w_120_176, w_055_213);
  nand2 I120_177(w_120_177, w_005_204, w_071_038);
  not1 I120_215(w_120_215, w_080_399);
  and2 I120_222(w_120_222, w_059_196, w_112_018);
  not1 I120_223(w_120_223, w_094_288);
  and2 I120_241(w_120_241, w_004_084, w_105_029);
  not1 I120_244(w_120_244, w_091_117);
  or2  I120_262(w_120_262, w_006_150, w_113_188);
  not1 I120_269(w_120_269, w_090_224);
  not1 I120_289(w_120_289, w_102_575);
  and2 I120_305(w_120_305, w_098_025, w_018_002);
  and2 I120_311(w_120_311, w_074_009, w_012_012);
  and2 I120_332(w_120_332, w_108_053, w_093_391);
  or2  I120_343(w_120_343, w_115_075, w_014_185);
  or2  I120_345(w_120_345, w_042_219, w_073_457);
  nand2 I120_348(w_120_348, w_086_133, w_099_044);
  not1 I120_353(w_120_353, w_068_242);
  and2 I120_402(w_120_402, w_060_122, w_016_003);
  or2  I120_410(w_120_410, w_004_336, w_042_227);
  nand2 I120_430(w_120_430, w_112_022, w_081_018);
  nand2 I120_439(w_120_439, w_025_235, w_037_055);
  nand2 I120_454(w_120_454, w_011_312, w_113_154);
  nand2 I120_480(w_120_480, w_104_138, w_109_383);
  and2 I120_489(w_120_489, w_072_199, w_012_152);
  and2 I120_506(w_120_506, w_015_555, w_081_007);
  or2  I120_516(w_120_516, w_004_187, w_089_136);
  not1 I120_517(w_120_517, w_092_220);
  not1 I120_528(w_120_528, w_063_188);
  and2 I120_545(w_120_545, w_054_157, w_032_033);
  or2  I120_558(w_120_558, w_041_513, w_081_022);
  and2 I120_569(w_120_569, w_067_360, w_056_675);
  and2 I120_578(w_120_578, w_018_029, w_106_206);
  nand2 I120_594(w_120_594, w_092_032, w_064_339);
  nand2 I120_604(w_120_604, w_106_062, w_049_083);
  and2 I120_612(w_120_612, w_084_037, w_102_462);
  nand2 I120_626(w_120_626, w_088_135, w_082_409);
  not1 I120_633(w_120_633, w_025_216);
  nand2 I120_638(w_120_638, w_078_033, w_072_172);
  or2  I120_648(w_120_648, w_063_107, w_000_159);
  nand2 I120_666(w_120_666, w_102_392, w_012_045);
  nand2 I120_674(w_120_674, w_099_213, w_005_130);
  and2 I120_681(w_120_681, w_035_081, w_029_087);
  nand2 I120_684(w_120_684, w_012_226, w_064_237);
  or2  I120_689(w_120_689, w_103_147, w_106_006);
  not1 I120_693(w_120_693, w_030_091);
  nand2 I120_695(w_120_695, w_084_036, w_012_072);
  and2 I120_734(w_120_734, w_110_125, w_097_130);
  nand2 I121_004(w_121_004, w_044_293, w_105_327);
  or2  I121_009(w_121_009, w_105_339, w_003_026);
  nand2 I121_011(w_121_011, w_074_099, w_103_128);
  and2 I121_027(w_121_027, w_099_053, w_092_530);
  or2  I121_032(w_121_032, w_034_017, w_100_084);
  or2  I121_039(w_121_039, w_051_230, w_053_080);
  not1 I121_045(w_121_045, w_089_071);
  not1 I121_047(w_121_047, w_037_059);
  nand2 I121_048(w_121_048, w_103_228, w_044_027);
  or2  I121_050(w_121_050, w_074_152, w_081_001);
  or2  I121_051(w_121_051, w_059_455, w_050_363);
  nand2 I121_053(w_121_053, w_063_180, w_075_127);
  not1 I121_054(w_121_054, w_112_000);
  or2  I121_055(w_121_055, w_095_038, w_094_044);
  nand2 I121_057(w_121_057, w_045_206, w_036_262);
  and2 I121_058(w_121_058, w_076_107, w_014_101);
  or2  I121_082(w_121_082, w_013_546, w_098_000);
  and2 I121_084(w_121_084, w_082_090, w_107_221);
  and2 I121_086(w_121_086, w_017_071, w_054_096);
  not1 I121_088(w_121_088, w_107_150);
  nand2 I121_106(w_121_106, w_028_547, w_039_680);
  or2  I121_112(w_121_112, w_097_035, w_022_243);
  nand2 I121_115(w_121_115, w_060_372, w_013_292);
  or2  I121_117(w_121_117, w_016_007, w_118_054);
  or2  I121_120(w_121_120, w_041_488, w_043_047);
  not1 I121_121(w_121_121, w_000_081);
  and2 I121_125(w_121_125, w_075_128, w_081_017);
  not1 I121_126(w_121_126, w_055_344);
  nand2 I121_127(w_121_127, w_096_005, w_102_445);
  or2  I121_128(w_121_128, w_102_526, w_008_358);
  and2 I121_129(w_121_129, w_076_183, w_024_118);
  or2  I121_134(w_121_134, w_030_204, w_086_144);
  not1 I121_136(w_121_136, w_072_288);
  and2 I121_141(w_121_141, w_010_221, w_036_136);
  not1 I121_144(w_121_144, w_014_005);
  or2  I121_160(w_121_160, w_113_031, w_079_038);
  not1 I121_161(w_121_161, w_104_158);
  or2  I121_162(w_121_162, w_095_010, w_063_383);
  and2 I121_168(w_121_168, w_116_261, w_052_007);
  or2  I121_174(w_121_174, w_062_526, w_050_392);
  not1 I121_189(w_121_189, w_046_314);
  nand2 I121_190(w_121_190, w_074_343, w_119_188);
  and2 I121_192(w_121_192, w_101_171, w_073_204);
  or2  I121_194(w_121_194, w_063_089, w_065_646);
  and2 I121_199(w_121_199, w_046_294, w_000_360);
  nand2 I121_202(w_121_202, w_093_256, w_017_345);
  or2  I121_206(w_121_206, w_059_202, w_041_057);
  or2  I121_209(w_121_209, w_089_107, w_092_272);
  or2  I121_210(w_121_210, w_060_086, w_021_202);
  and2 I121_211(w_121_211, w_082_546, w_108_201);
  not1 I122_000(w_122_000, w_037_339);
  nand2 I122_001(w_122_001, w_029_008, w_053_038);
  not1 I122_005(w_122_005, w_024_088);
  nand2 I122_008(w_122_008, w_004_019, w_064_114);
  and2 I122_009(w_122_009, w_103_076, w_004_035);
  not1 I122_010(w_122_010, w_068_226);
  not1 I122_012(w_122_012, w_014_005);
  not1 I122_014(w_122_014, w_073_601);
  or2  I122_017(w_122_017, w_019_006, w_004_005);
  nand2 I122_020(w_122_020, w_116_126, w_070_018);
  and2 I122_021(w_122_021, w_024_121, w_089_211);
  and2 I122_022(w_122_022, w_090_068, w_050_054);
  and2 I122_026(w_122_026, w_053_137, w_005_307);
  nand2 I122_027(w_122_027, w_078_106, w_088_129);
  and2 I122_030(w_122_030, w_027_168, w_034_026);
  or2  I122_031(w_122_031, w_075_141, w_069_153);
  nand2 I122_032(w_122_032, w_053_054, w_054_494);
  and2 I122_034(w_122_034, w_094_114, w_078_089);
  or2  I122_035(w_122_035, w_012_003, w_080_403);
  not1 I122_040(w_122_040, w_082_323);
  not1 I122_041(w_122_041, w_100_031);
  or2  I122_049(w_122_049, w_009_305, w_092_650);
  or2  I122_055(w_122_055, w_119_067, w_054_029);
  not1 I122_056(w_122_056, w_066_125);
  and2 I122_058(w_122_058, w_103_068, w_095_008);
  nand2 I122_060(w_122_060, w_016_007, w_022_407);
  or2  I122_063(w_122_063, w_107_003, w_105_346);
  not1 I122_065(w_122_065, w_111_011);
  or2  I122_066(w_122_066, w_092_324, w_061_101);
  and2 I122_067(w_122_067, w_077_398, w_018_042);
  and2 I122_072(w_122_072, w_018_030, w_019_002);
  and2 I122_074(w_122_074, w_067_346, w_117_010);
  or2  I122_081(w_122_081, w_101_089, w_067_062);
  and2 I122_082(w_122_082, w_037_140, w_029_004);
  nand2 I122_083(w_122_083, w_035_097, w_097_566);
  not1 I122_084(w_122_084, w_077_483);
  nand2 I122_086(w_122_086, w_001_020, w_092_287);
  not1 I122_089(w_122_089, w_088_024);
  or2  I122_090(w_122_090, w_039_567, w_110_135);
  or2  I122_091(w_122_091, w_050_454, w_090_035);
  not1 I122_093(w_122_093, w_006_223);
  not1 I122_094(w_122_094, w_088_143);
  or2  I122_102(w_122_102, w_106_199, w_001_006);
  or2  I122_103(w_122_103, w_009_197, w_051_242);
  and2 I122_113(w_122_113, w_074_256, w_114_188);
  or2  I122_120(w_122_120, w_063_219, w_046_029);
  not1 I122_121(w_122_121, w_018_039);
  not1 I122_126(w_122_126, w_033_724);
  not1 I123_005(w_123_005, w_039_301);
  nand2 I123_013(w_123_013, w_025_084, w_097_042);
  nand2 I123_016(w_123_016, w_032_091, w_078_104);
  or2  I123_029(w_123_029, w_060_291, w_008_258);
  and2 I123_036(w_123_036, w_121_117, w_015_177);
  and2 I123_053(w_123_053, w_103_123, w_043_035);
  and2 I123_056(w_123_056, w_027_122, w_016_003);
  not1 I123_067(w_123_067, w_091_043);
  nand2 I123_087(w_123_087, w_021_026, w_036_313);
  or2  I123_096(w_123_096, w_007_263, w_085_045);
  and2 I123_097(w_123_097, w_004_469, w_018_018);
  nand2 I123_101(w_123_101, w_079_007, w_017_426);
  and2 I123_104(w_123_104, w_067_134, w_102_618);
  nand2 I123_112(w_123_112, w_107_302, w_084_039);
  or2  I123_122(w_123_122, w_047_436, w_099_135);
  or2  I123_139(w_123_139, w_095_008, w_038_095);
  or2  I123_149(w_123_149, w_090_505, w_003_048);
  nand2 I123_153(w_123_153, w_103_162, w_102_304);
  not1 I123_162(w_123_162, w_113_109);
  or2  I123_169(w_123_169, w_008_485, w_087_311);
  and2 I123_172(w_123_172, w_103_191, w_098_027);
  not1 I123_174(w_123_174, w_054_162);
  or2  I123_187(w_123_187, w_120_734, w_036_282);
  not1 I123_195(w_123_195, w_108_203);
  and2 I123_251(w_123_251, w_037_085, w_081_013);
  nand2 I123_255(w_123_255, w_007_179, w_085_038);
  or2  I123_297(w_123_297, w_111_012, w_078_112);
  or2  I123_302(w_123_302, w_117_018, w_079_016);
  not1 I123_304(w_123_304, w_104_271);
  not1 I123_364(w_123_364, w_073_018);
  not1 I123_367(w_123_367, w_061_230);
  or2  I123_369(w_123_369, w_010_677, w_061_380);
  and2 I123_379(w_123_379, w_006_093, w_098_044);
  or2  I123_388(w_123_388, w_069_049, w_106_054);
  not1 I123_459(w_123_459, w_057_155);
  not1 I123_471(w_123_471, w_098_065);
  not1 I123_481(w_123_481, w_097_195);
  not1 I123_503(w_123_503, w_020_183);
  and2 I123_505(w_123_505, w_029_069, w_064_059);
  nand2 I123_511(w_123_511, w_022_399, w_030_061);
  nand2 I123_532(w_123_532, w_122_008, w_019_016);
  and2 I123_538(w_123_538, w_007_155, w_082_455);
  or2  I123_584(w_123_584, w_067_250, w_025_157);
  nand2 I123_592(w_123_592, w_024_093, w_018_028);
  nand2 I124_001(w_124_001, w_112_130, w_014_030);
  or2  I124_025(w_124_025, w_052_021, w_011_025);
  or2  I124_027(w_124_027, w_008_696, w_018_042);
  or2  I124_035(w_124_035, w_075_152, w_085_329);
  not1 I124_046(w_124_046, w_070_412);
  nand2 I124_052(w_124_052, w_027_033, w_053_066);
  or2  I124_056(w_124_056, w_005_052, w_078_446);
  and2 I124_057(w_124_057, w_105_045, w_043_000);
  not1 I124_061(w_124_061, w_113_050);
  and2 I124_065(w_124_065, w_102_542, w_025_160);
  not1 I124_070(w_124_070, w_043_035);
  nand2 I124_078(w_124_078, w_105_265, w_116_079);
  nand2 I124_089(w_124_089, w_089_199, w_111_041);
  and2 I124_091(w_124_091, w_013_141, w_000_264);
  not1 I124_094(w_124_094, w_026_331);
  not1 I124_096(w_124_096, w_027_131);
  or2  I124_104(w_124_104, w_101_020, w_048_018);
  not1 I124_105(w_124_105, w_087_335);
  nand2 I124_108(w_124_108, w_058_075, w_099_036);
  and2 I124_109(w_124_109, w_074_243, w_040_521);
  or2  I124_112(w_124_112, w_101_083, w_082_235);
  or2  I124_114(w_124_114, w_115_065, w_112_006);
  not1 I124_116(w_124_116, w_002_163);
  and2 I124_122(w_124_122, w_032_204, w_006_120);
  not1 I124_134(w_124_134, w_037_305);
  not1 I124_143(w_124_143, w_063_181);
  nand2 I124_145(w_124_145, w_110_117, w_011_409);
  not1 I124_156(w_124_156, w_074_227);
  or2  I124_171(w_124_171, w_016_003, w_002_354);
  nand2 I124_217(w_124_217, w_068_280, w_011_189);
  nand2 I124_220(w_124_220, w_008_183, w_019_018);
  and2 I124_232(w_124_232, w_087_100, w_066_595);
  and2 I124_242(w_124_242, w_050_133, w_100_051);
  and2 I124_244(w_124_244, w_031_251, w_025_199);
  not1 I124_252(w_124_252, w_081_003);
  and2 I124_256(w_124_256, w_033_116, w_058_479);
  or2  I124_273(w_124_273, w_108_174, w_019_000);
  or2  I124_281(w_124_281, w_123_369, w_061_059);
  nand2 I124_286(w_124_286, w_043_004, w_006_029);
  or2  I124_287(w_124_287, w_088_025, w_045_227);
  and2 I124_291(w_124_291, w_090_223, w_072_235);
  not1 I124_295(w_124_295, w_116_513);
  nand2 I124_319(w_124_319, w_072_165, w_015_041);
  nand2 I124_328(w_124_328, w_111_034, w_008_027);
  not1 I124_330(w_124_330, w_020_482);
  or2  I125_003(w_125_003, w_094_380, w_074_221);
  or2  I125_025(w_125_025, w_066_503, w_074_287);
  not1 I125_030(w_125_030, w_034_066);
  or2  I125_031(w_125_031, w_084_005, w_015_603);
  or2  I125_036(w_125_036, w_036_148, w_048_013);
  or2  I125_057(w_125_057, w_027_164, w_061_005);
  and2 I125_059(w_125_059, w_042_261, w_070_018);
  nand2 I125_065(w_125_065, w_097_360, w_033_646);
  not1 I125_069(w_125_069, w_083_175);
  or2  I125_072(w_125_072, w_008_682, w_070_329);
  not1 I125_079(w_125_079, w_071_317);
  nand2 I125_081(w_125_081, w_045_166, w_048_010);
  or2  I125_084(w_125_084, w_104_042, w_065_565);
  not1 I125_118(w_125_118, w_024_523);
  not1 I125_124(w_125_124, w_107_109);
  or2  I125_128(w_125_128, w_001_007, w_103_075);
  or2  I125_129(w_125_129, w_066_110, w_021_010);
  nand2 I125_138(w_125_138, w_035_124, w_067_005);
  not1 I125_150(w_125_150, w_037_153);
  or2  I125_187(w_125_187, w_095_018, w_044_499);
  not1 I125_191(w_125_191, w_022_207);
  not1 I125_193(w_125_193, w_058_017);
  not1 I125_204(w_125_204, w_008_159);
  not1 I125_208(w_125_208, w_108_190);
  and2 I125_224(w_125_224, w_079_010, w_032_165);
  not1 I125_242(w_125_242, w_093_081);
  and2 I125_282(w_125_282, w_049_131, w_040_611);
  nand2 I125_297(w_125_297, w_012_300, w_063_193);
  not1 I125_308(w_125_308, w_118_079);
  or2  I125_318(w_125_318, w_016_000, w_122_027);
  or2  I125_332(w_125_332, w_058_477, w_041_113);
  and2 I125_347(w_125_347, w_077_176, w_073_503);
  not1 I125_354(w_125_354, w_107_238);
  or2  I125_386(w_125_386, w_117_012, w_109_054);
  and2 I125_397(w_125_397, w_052_024, w_009_528);
  nand2 I125_399(w_125_399, w_055_096, w_089_230);
  or2  I125_417(w_125_417, w_112_095, w_030_159);
  nand2 I125_439(w_125_439, w_080_233, w_038_043);
  or2  I125_446(w_125_446, w_055_181, w_044_398);
  or2  I125_466(w_125_466, w_007_395, w_120_480);
  not1 I125_497(w_125_497, w_103_067);
  nand2 I125_561(w_125_561, w_050_149, w_046_604);
  not1 I125_586(w_125_586, w_035_116);
  or2  I126_008(w_126_008, w_092_610, w_105_182);
  not1 I126_013(w_126_013, w_084_042);
  and2 I126_017(w_126_017, w_053_154, w_104_354);
  and2 I126_018(w_126_018, w_007_014, w_070_041);
  nand2 I126_024(w_126_024, w_113_171, w_025_251);
  or2  I126_027(w_126_027, w_120_454, w_020_502);
  or2  I126_028(w_126_028, w_044_122, w_000_448);
  not1 I126_034(w_126_034, w_020_452);
  nand2 I126_037(w_126_037, w_041_549, w_045_293);
  and2 I126_038(w_126_038, w_114_211, w_055_174);
  and2 I126_041(w_126_041, w_058_229, w_119_125);
  or2  I126_047(w_126_047, w_080_336, w_067_060);
  and2 I126_055(w_126_055, w_040_478, w_052_032);
  nand2 I126_056(w_126_056, w_032_031, w_096_000);
  nand2 I126_058(w_126_058, w_019_016, w_027_074);
  nand2 I126_061(w_126_061, w_050_597, w_075_091);
  not1 I126_063(w_126_063, w_101_303);
  or2  I126_064(w_126_064, w_051_157, w_008_584);
  nand2 I126_068(w_126_068, w_047_379, w_077_272);
  and2 I126_073(w_126_073, w_005_275, w_038_054);
  nand2 I126_078(w_126_078, w_113_120, w_034_059);
  nand2 I126_079(w_126_079, w_083_043, w_038_377);
  nand2 I126_082(w_126_082, w_063_301, w_033_217);
  nand2 I126_084(w_126_084, w_038_496, w_032_364);
  or2  I126_090(w_126_090, w_051_008, w_075_111);
  not1 I126_092(w_126_092, w_058_074);
  nand2 I126_095(w_126_095, w_111_003, w_044_562);
  nand2 I126_100(w_126_100, w_076_296, w_007_439);
  nand2 I126_104(w_126_104, w_004_148, w_120_269);
  nand2 I126_112(w_126_112, w_097_077, w_100_066);
  not1 I126_115(w_126_115, w_114_209);
  not1 I126_116(w_126_116, w_084_037);
  or2  I126_117(w_126_117, w_015_029, w_005_096);
  not1 I126_119(w_126_119, w_018_005);
  not1 I126_120(w_126_120, w_063_424);
  nand2 I126_127(w_126_127, w_024_157, w_012_264);
  nand2 I126_128(w_126_128, w_069_225, w_008_335);
  or2  I126_130(w_126_130, w_002_027, w_077_619);
  nand2 I126_133(w_126_133, w_075_033, w_015_501);
  or2  I126_135(w_126_135, w_043_021, w_103_136);
  not1 I126_139(w_126_139, w_085_092);
  nand2 I126_142(w_126_142, w_008_653, w_067_111);
  and2 I126_144(w_126_144, w_078_421, w_014_234);
  or2  I126_153(w_126_153, w_110_087, w_095_022);
  and2 I126_154(w_126_154, w_122_012, w_052_041);
  and2 I126_158(w_126_158, w_071_305, w_077_254);
  or2  I126_164(w_126_164, w_080_154, w_101_070);
  or2  I126_175(w_126_175, w_013_469, w_096_004);
  nand2 I126_187(w_126_187, w_028_473, w_023_199);
  nand2 I126_193(w_126_193, w_113_132, w_034_044);
  nand2 I127_000(w_127_000, w_043_041, w_071_281);
  and2 I127_003(w_127_003, w_040_050, w_096_002);
  and2 I127_004(w_127_004, w_016_008, w_014_176);
  or2  I127_007(w_127_007, w_032_066, w_108_000);
  not1 I127_008(w_127_008, w_022_368);
  not1 I127_011(w_127_011, w_022_045);
  and2 I127_015(w_127_015, w_095_029, w_070_482);
  not1 I127_017(w_127_017, w_072_084);
  and2 I127_018(w_127_018, w_046_450, w_018_037);
  nand2 I127_022(w_127_022, w_036_179, w_099_222);
  and2 I127_025(w_127_025, w_022_399, w_099_011);
  not1 I127_026(w_127_026, w_117_053);
  and2 I127_027(w_127_027, w_025_227, w_099_081);
  and2 I127_031(w_127_031, w_067_362, w_019_001);
  nand2 I127_034(w_127_034, w_089_138, w_105_248);
  or2  I127_035(w_127_035, w_096_000, w_102_204);
  and2 I127_038(w_127_038, w_049_187, w_012_314);
  or2  I127_041(w_127_041, w_009_503, w_036_068);
  nand2 I127_043(w_127_043, w_042_292, w_060_336);
  or2  I127_044(w_127_044, w_067_336, w_035_119);
  or2  I127_047(w_127_047, w_020_038, w_107_068);
  or2  I127_048(w_127_048, w_008_576, w_107_130);
  and2 I127_052(w_127_052, w_028_072, w_069_171);
  nand2 I127_053(w_127_053, w_082_214, w_024_051);
  and2 I127_054(w_127_054, w_036_023, w_077_382);
  not1 I127_057(w_127_057, w_057_145);
  or2  I127_061(w_127_061, w_035_018, w_021_139);
  not1 I127_065(w_127_065, w_073_382);
  and2 I127_067(w_127_067, w_118_101, w_034_019);
  and2 I127_069(w_127_069, w_063_227, w_035_070);
  nand2 I127_070(w_127_070, w_095_039, w_063_045);
  nand2 I127_071(w_127_071, w_123_101, w_028_277);
  not1 I127_073(w_127_073, w_109_291);
  or2  I127_074(w_127_074, w_016_001, w_053_077);
  or2  I128_000(w_128_000, w_032_137, w_066_134);
  and2 I128_010(w_128_010, w_048_011, w_091_020);
  not1 I128_021(w_128_021, w_057_053);
  nand2 I128_022(w_128_022, w_086_160, w_093_035);
  not1 I128_025(w_128_025, w_091_117);
  and2 I128_026(w_128_026, w_084_005, w_077_052);
  and2 I128_035(w_128_035, w_027_197, w_079_010);
  nand2 I128_048(w_128_048, w_087_204, w_013_099);
  or2  I128_051(w_128_051, w_029_031, w_019_001);
  not1 I128_055(w_128_055, w_040_488);
  or2  I128_067(w_128_067, w_072_134, w_110_064);
  not1 I128_070(w_128_070, w_092_131);
  and2 I128_073(w_128_073, w_006_115, w_077_057);
  nand2 I128_091(w_128_091, w_098_069, w_098_059);
  or2  I128_094(w_128_094, w_018_001, w_098_059);
  nand2 I128_103(w_128_103, w_105_218, w_048_016);
  and2 I128_111(w_128_111, w_060_038, w_049_081);
  and2 I128_115(w_128_115, w_021_041, w_124_217);
  or2  I128_122(w_128_122, w_019_010, w_083_067);
  nand2 I128_130(w_128_130, w_039_470, w_124_114);
  and2 I128_139(w_128_139, w_006_014, w_085_201);
  or2  I128_140(w_128_140, w_099_062, w_060_246);
  nand2 I128_152(w_128_152, w_014_280, w_120_517);
  nand2 I128_157(w_128_157, w_050_406, w_087_258);
  not1 I128_174(w_128_174, w_116_373);
  not1 I128_181(w_128_181, w_082_175);
  not1 I128_187(w_128_187, w_023_096);
  and2 I128_191(w_128_191, w_084_024, w_085_294);
  and2 I128_195(w_128_195, w_082_270, w_091_125);
  not1 I128_196(w_128_196, w_108_207);
  nand2 I128_233(w_128_233, w_003_039, w_047_237);
  and2 I128_234(w_128_234, w_104_168, w_028_013);
  or2  I128_268(w_128_268, w_065_348, w_108_122);
  not1 I128_291(w_128_291, w_124_001);
  or2  I128_295(w_128_295, w_078_013, w_102_555);
  and2 I128_297(w_128_297, w_051_265, w_090_171);
  not1 I128_306(w_128_306, w_040_080);
  and2 I128_318(w_128_318, w_017_636, w_110_318);
  not1 I128_327(w_128_327, w_018_038);
  or2  I128_329(w_128_329, w_075_058, w_127_003);
  and2 I128_345(w_128_345, w_029_083, w_105_192);
  and2 I128_353(w_128_353, w_073_627, w_055_219);
  or2  I128_380(w_128_380, w_032_138, w_069_042);
  nand2 I128_411(w_128_411, w_033_269, w_040_505);
  nand2 I128_414(w_128_414, w_050_271, w_052_042);
  or2  I128_417(w_128_417, w_092_191, w_082_389);
  nand2 I128_426(w_128_426, w_090_048, w_079_004);
  not1 I128_464(w_128_464, w_117_005);
  or2  I128_495(w_128_495, w_111_007, w_038_548);
  and2 I128_496(w_128_496, w_114_195, w_044_652);
  not1 I128_524(w_128_524, w_074_293);
  and2 I128_559(w_128_559, w_119_099, w_032_091);
  nand2 I128_571(w_128_571, w_000_582, w_039_170);
  and2 I128_580(w_128_580, w_027_111, w_114_141);
  and2 I128_608(w_128_608, w_047_248, w_090_451);
  nand2 I128_638(w_128_638, w_065_046, w_126_037);
  nand2 I128_640(w_128_640, w_068_079, w_099_150);
  not1 I129_005(w_129_005, w_092_046);
  not1 I129_017(w_129_017, w_045_172);
  nand2 I129_023(w_129_023, w_010_568, w_087_255);
  not1 I129_029(w_129_029, w_014_109);
  and2 I129_034(w_129_034, w_101_246, w_000_326);
  nand2 I129_041(w_129_041, w_027_124, w_031_466);
  or2  I129_044(w_129_044, w_024_434, w_047_390);
  not1 I129_048(w_129_048, w_012_323);
  and2 I129_065(w_129_065, w_116_636, w_017_206);
  and2 I129_067(w_129_067, w_046_118, w_046_097);
  nand2 I129_072(w_129_072, w_124_319, w_051_183);
  not1 I129_078(w_129_078, w_106_101);
  nand2 I129_082(w_129_082, w_018_027, w_087_195);
  nand2 I129_087(w_129_087, w_071_109, w_013_114);
  not1 I129_088(w_129_088, w_122_056);
  and2 I129_090(w_129_090, w_110_352, w_027_132);
  or2  I129_095(w_129_095, w_100_077, w_128_638);
  nand2 I129_100(w_129_100, w_118_030, w_073_489);
  not1 I129_106(w_129_106, w_067_156);
  not1 I129_108(w_129_108, w_074_309);
  nand2 I129_111(w_129_111, w_126_028, w_090_117);
  and2 I129_113(w_129_113, w_085_011, w_024_258);
  nand2 I129_117(w_129_117, w_001_001, w_126_084);
  not1 I129_120(w_129_120, w_071_082);
  not1 I129_133(w_129_133, w_119_014);
  not1 I129_135(w_129_135, w_119_171);
  nand2 I129_140(w_129_140, w_068_344, w_093_132);
  or2  I129_149(w_129_149, w_005_002, w_099_087);
  and2 I129_156(w_129_156, w_090_221, w_107_345);
  or2  I129_164(w_129_164, w_005_095, w_109_068);
  or2  I129_168(w_129_168, w_045_007, w_123_016);
  nand2 I129_170(w_129_170, w_119_053, w_065_028);
  nand2 I129_175(w_129_175, w_041_154, w_053_080);
  nand2 I129_180(w_129_180, w_066_276, w_121_115);
  nand2 I129_182(w_129_182, w_114_135, w_009_424);
  nand2 I129_186(w_129_186, w_006_004, w_119_103);
  or2  I129_198(w_129_198, w_002_702, w_068_024);
  nand2 I129_204(w_129_204, w_104_233, w_094_006);
  not1 I129_205(w_129_205, w_097_131);
  or2  I129_210(w_129_210, w_127_025, w_102_553);
  not1 I129_216(w_129_216, w_058_359);
  or2  I129_226(w_129_226, w_003_071, w_074_077);
  or2  I129_245(w_129_245, w_083_098, w_109_104);
  or2  I129_251(w_129_251, w_096_002, w_005_091);
  not1 I129_256(w_129_256, w_086_029);
  nand2 I129_275(w_129_275, w_002_074, w_070_213);
  nand2 I129_276(w_129_276, w_078_112, w_020_226);
  not1 I129_278(w_129_278, w_064_202);
  or2  I129_282(w_129_282, w_102_188, w_010_451);
  not1 I129_289(w_129_289, w_118_071);
  and2 I129_293(w_129_293, w_006_057, w_060_164);
  or2  I129_295(w_129_295, w_053_114, w_064_064);
  not1 I129_305(w_129_305, w_104_321);
  not1 I129_313(w_129_313, w_028_136);
  or2  I129_329(w_129_329, w_047_199, w_039_493);
  not1 I129_333(w_129_333, w_116_001);
  or2  I129_337(w_129_337, w_049_238, w_006_132);
  nand2 I129_342(w_129_342, w_122_020, w_005_125);
  or2  I129_348(w_129_348, w_019_010, w_054_310);
  or2  I129_349(w_129_349, w_052_035, w_052_004);
  and2 I129_351(w_129_351, w_002_529, w_048_008);
  not1 I129_353(w_129_353, w_120_689);
  nand2 I129_372(w_129_372, w_019_001, w_033_639);
  not1 I129_414(w_129_414, w_074_231);
  and2 I130_005(w_130_005, w_108_143, w_121_206);
  and2 I130_023(w_130_023, w_128_411, w_036_309);
  or2  I130_033(w_130_033, w_028_076, w_033_358);
  or2  I130_035(w_130_035, w_103_007, w_100_087);
  or2  I130_044(w_130_044, w_035_046, w_019_001);
  and2 I130_046(w_130_046, w_033_082, w_122_083);
  not1 I130_049(w_130_049, w_035_087);
  or2  I130_071(w_130_071, w_036_109, w_031_375);
  nand2 I130_075(w_130_075, w_045_092, w_059_660);
  nand2 I130_088(w_130_088, w_066_101, w_081_012);
  nand2 I130_089(w_130_089, w_004_507, w_071_104);
  not1 I130_122(w_130_122, w_075_055);
  not1 I130_134(w_130_134, w_108_097);
  and2 I130_171(w_130_171, w_023_135, w_052_000);
  and2 I130_184(w_130_184, w_079_024, w_124_089);
  not1 I130_191(w_130_191, w_088_060);
  not1 I130_194(w_130_194, w_120_029);
  nand2 I130_195(w_130_195, w_101_121, w_005_073);
  or2  I130_204(w_130_204, w_051_183, w_030_330);
  and2 I130_211(w_130_211, w_042_001, w_118_093);
  not1 I130_212(w_130_212, w_096_005);
  and2 I130_220(w_130_220, w_083_066, w_085_265);
  not1 I130_230(w_130_230, w_124_328);
  not1 I130_236(w_130_236, w_046_052);
  nand2 I130_239(w_130_239, w_022_103, w_127_044);
  or2  I130_252(w_130_252, w_009_223, w_066_544);
  not1 I130_254(w_130_254, w_020_022);
  not1 I130_260(w_130_260, w_126_139);
  or2  I130_264(w_130_264, w_096_001, w_045_157);
  or2  I130_278(w_130_278, w_123_511, w_074_070);
  not1 I130_280(w_130_280, w_058_292);
  or2  I130_283(w_130_283, w_099_054, w_071_260);
  nand2 I130_294(w_130_294, w_027_165, w_060_261);
  nand2 I130_295(w_130_295, w_028_437, w_034_012);
  not1 I130_321(w_130_321, w_030_292);
  nand2 I130_375(w_130_375, w_099_240, w_013_054);
  or2  I130_377(w_130_377, w_042_310, w_094_038);
  or2  I130_391(w_130_391, w_056_523, w_040_051);
  and2 I130_408(w_130_408, w_051_081, w_074_114);
  not1 I130_418(w_130_418, w_117_026);
  not1 I130_463(w_130_463, w_085_139);
  not1 I130_469(w_130_469, w_000_702);
  or2  I130_499(w_130_499, w_098_047, w_056_642);
  and2 I130_511(w_130_511, w_014_108, w_036_123);
  not1 I130_517(w_130_519, w_130_518);
  nand2 I130_518(w_130_520, w_030_191, w_130_519);
  or2  I130_519(w_130_521, w_130_520, w_029_018);
  nand2 I130_520(w_130_522, w_028_411, w_130_521);
  nand2 I130_521(w_130_523, w_088_023, w_130_522);
  and2 I130_522(w_130_524, w_130_523, w_130_538);
  nand2 I130_523(w_130_518, w_130_524, w_042_134);
  not1 I130_524(w_130_529, w_130_528);
  and2 I130_525(w_130_530, w_013_496, w_130_529);
  or2  I130_526(w_130_531, w_001_032, w_130_530);
  or2  I130_527(w_130_532, w_095_041, w_130_531);
  and2 I130_528(w_130_533, w_037_166, w_130_532);
  and2 I130_529(w_130_534, w_046_472, w_130_533);
  not1 I130_530(w_130_535, w_130_534);
  and2 I130_531(w_130_536, w_055_258, w_130_535);
  not1 I130_532(w_130_528, w_130_524);
  and2 I130_533(w_130_538, w_082_092, w_130_536);
  nand2 I131_000(w_131_000, w_089_266, w_056_249);
  nand2 I131_007(w_131_007, w_097_252, w_125_118);
  or2  I131_029(w_131_029, w_035_031, w_034_042);
  and2 I131_037(w_131_037, w_041_304, w_009_480);
  nand2 I131_040(w_131_040, w_012_051, w_011_521);
  nand2 I131_048(w_131_048, w_120_528, w_085_295);
  not1 I131_053(w_131_053, w_030_301);
  not1 I131_054(w_131_054, w_068_069);
  not1 I131_059(w_131_059, w_089_129);
  or2  I131_071(w_131_071, w_055_023, w_052_014);
  or2  I131_073(w_131_073, w_040_551, w_045_117);
  not1 I131_087(w_131_087, w_031_308);
  and2 I131_092(w_131_092, w_053_102, w_104_264);
  nand2 I131_101(w_131_101, w_121_032, w_037_303);
  or2  I131_109(w_131_109, w_021_060, w_055_185);
  nand2 I131_113(w_131_113, w_078_063, w_039_121);
  not1 I131_120(w_131_120, w_118_012);
  or2  I131_121(w_131_121, w_029_065, w_070_471);
  not1 I131_140(w_131_140, w_008_414);
  and2 I131_144(w_131_144, w_108_205, w_038_097);
  nand2 I131_147(w_131_147, w_009_120, w_027_015);
  and2 I131_149(w_131_149, w_106_083, w_087_071);
  nand2 I131_187(w_131_187, w_107_279, w_097_108);
  or2  I131_212(w_131_212, w_055_027, w_021_122);
  not1 I131_223(w_131_223, w_005_125);
  not1 I131_254(w_131_254, w_030_207);
  or2  I131_263(w_131_263, w_130_236, w_110_032);
  and2 I131_269(w_131_269, w_013_334, w_083_151);
  not1 I131_285(w_131_285, w_040_514);
  not1 I131_303(w_131_303, w_031_434);
  not1 I131_304(w_131_304, w_115_135);
  nand2 I131_308(w_131_308, w_077_165, w_043_002);
  or2  I131_318(w_131_318, w_093_186, w_050_011);
  and2 I131_345(w_131_345, w_110_090, w_069_096);
  not1 I131_430(w_131_430, w_104_260);
  or2  I131_431(w_131_431, w_053_149, w_071_107);
  not1 I131_432(w_131_432, w_130_005);
  and2 I131_450(w_131_450, w_032_180, w_114_170);
  and2 I131_472(w_131_472, w_060_155, w_098_028);
  or2  I131_480(w_131_480, w_090_362, w_098_036);
  and2 I131_483(w_131_483, w_026_005, w_122_090);
  not1 I131_486(w_131_486, w_096_002);
  not1 I131_511(w_131_511, w_126_008);
  nand2 I131_545(w_131_545, w_110_363, w_103_023);
  or2  I131_557(w_131_557, w_111_102, w_085_162);
  nand2 I131_566(w_131_566, w_077_060, w_080_052);
  not1 I132_012(w_132_012, w_024_219);
  not1 I132_026(w_132_026, w_052_037);
  nand2 I132_031(w_132_031, w_024_187, w_016_002);
  or2  I132_056(w_132_056, w_049_190, w_061_175);
  or2  I132_059(w_132_059, w_021_009, w_074_342);
  or2  I132_076(w_132_076, w_094_399, w_074_210);
  not1 I132_077(w_132_077, w_045_139);
  not1 I132_082(w_132_082, w_107_258);
  or2  I132_084(w_132_084, w_011_147, w_003_016);
  nand2 I132_087(w_132_087, w_086_098, w_016_003);
  or2  I132_089(w_132_089, w_063_319, w_061_266);
  nand2 I132_094(w_132_094, w_031_155, w_129_414);
  or2  I132_099(w_132_099, w_129_164, w_064_280);
  or2  I132_115(w_132_115, w_095_046, w_109_264);
  or2  I132_129(w_132_129, w_008_232, w_002_064);
  and2 I132_130(w_132_130, w_107_094, w_045_390);
  nand2 I132_152(w_132_152, w_029_096, w_113_061);
  nand2 I132_155(w_132_155, w_095_043, w_068_095);
  or2  I132_165(w_132_165, w_096_000, w_088_131);
  nand2 I132_179(w_132_179, w_116_420, w_104_178);
  nand2 I132_180(w_132_180, w_129_216, w_010_758);
  or2  I132_188(w_132_188, w_108_183, w_075_047);
  nand2 I132_196(w_132_196, w_022_161, w_047_154);
  or2  I132_202(w_132_202, w_059_588, w_085_068);
  not1 I132_204(w_132_204, w_063_213);
  or2  I132_206(w_132_206, w_053_023, w_051_333);
  or2  I132_217(w_132_217, w_113_227, w_106_144);
  not1 I132_219(w_132_219, w_127_057);
  nand2 I132_229(w_132_229, w_113_309, w_012_015);
  or2  I132_231(w_132_231, w_049_279, w_008_118);
  nand2 I132_249(w_132_249, w_051_342, w_004_284);
  nand2 I132_255(w_132_255, w_128_140, w_010_515);
  or2  I132_260(w_132_260, w_044_098, w_063_123);
  nand2 I132_262(w_132_262, w_085_277, w_059_521);
  and2 I132_281(w_132_281, w_102_068, w_010_187);
  nand2 I132_289(w_132_289, w_074_166, w_007_397);
  or2  I132_291(w_132_291, w_042_334, w_077_210);
  nand2 I132_305(w_132_305, w_086_237, w_001_006);
  nand2 I132_313(w_132_313, w_026_181, w_095_054);
  or2  I132_330(w_132_330, w_120_289, w_023_189);
  nand2 I132_331(w_132_331, w_100_074, w_101_066);
  not1 I132_333(w_132_333, w_002_692);
  and2 I132_384(w_132_384, w_064_165, w_131_318);
  not1 I132_386(w_132_386, w_077_019);
  nand2 I132_390(w_132_390, w_092_277, w_025_122);
  nand2 I132_393(w_132_393, w_123_388, w_076_074);
  nand2 I132_395(w_132_395, w_035_049, w_053_013);
  not1 I132_398(w_132_398, w_046_197);
  not1 I132_406(w_132_406, w_105_097);
  and2 I132_415(w_132_415, w_101_107, w_105_199);
  and2 I132_422(w_132_422, w_073_428, w_097_088);
  and2 I132_435(w_132_435, w_078_514, w_089_009);
  and2 I132_466(w_132_468, w_132_467, w_132_483);
  and2 I132_467(w_132_469, w_014_198, w_132_468);
  and2 I132_468(w_132_470, w_132_469, w_083_169);
  and2 I132_469(w_132_471, w_132_470, w_093_032);
  not1 I132_470(w_132_467, w_132_471);
  nand2 I132_471(w_132_476, w_101_307, w_132_475);
  or2  I132_472(w_132_477, w_127_065, w_132_476);
  and2 I132_473(w_132_478, w_132_477, w_033_321);
  and2 I132_474(w_132_479, w_132_478, w_120_545);
  nand2 I132_475(w_132_480, w_042_194, w_132_479);
  and2 I132_476(w_132_481, w_124_057, w_132_480);
  not1 I132_477(w_132_475, w_132_468);
  and2 I132_478(w_132_483, w_089_085, w_132_481);
  and2 I132_479(w_132_486, w_132_485, w_050_263);
  not1 I132_480(w_132_487, w_132_486);
  or2  I132_481(w_132_488, w_068_182, w_132_487);
  and2 I132_482(w_132_489, w_039_289, w_132_488);
  or2  I132_483(w_132_490, w_132_489, w_001_004);
  nand2 I132_484(w_132_491, w_132_490, w_039_264);
  and2 I132_485(w_132_492, w_072_057, w_132_491);
  and2 I132_486(w_132_493, w_132_492, w_066_011);
  or2  I132_487(w_132_494, w_132_493, w_105_284);
  nand2 I132_488(w_132_495, w_022_210, w_132_494);
  and2 I132_489(w_132_496, w_132_495, w_089_025);
  nand2 I132_490(w_132_485, w_132_496, w_095_005);
  nand2 I133_000(w_133_000, w_052_037, w_122_049);
  not1 I133_003(w_133_003, w_128_187);
  not1 I133_028(w_133_028, w_060_073);
  not1 I133_057(w_133_057, w_001_021);
  nand2 I133_061(w_133_061, w_085_042, w_001_004);
  not1 I133_066(w_133_066, w_099_261);
  nand2 I133_081(w_133_081, w_084_013, w_132_386);
  or2  I133_085(w_133_085, w_021_072, w_007_168);
  nand2 I133_095(w_133_095, w_085_056, w_129_108);
  not1 I133_097(w_133_097, w_022_232);
  or2  I133_099(w_133_099, w_010_616, w_115_151);
  or2  I133_117(w_133_117, w_051_036, w_119_086);
  nand2 I133_120(w_133_120, w_033_100, w_046_509);
  nand2 I133_134(w_133_134, w_102_601, w_077_282);
  or2  I133_143(w_133_143, w_016_001, w_063_400);
  nand2 I133_159(w_133_159, w_014_291, w_038_491);
  and2 I133_187(w_133_187, w_064_279, w_084_045);
  or2  I133_201(w_133_201, w_033_263, w_014_134);
  nand2 I133_223(w_133_223, w_052_031, w_095_014);
  and2 I133_235(w_133_235, w_044_019, w_029_033);
  and2 I133_244(w_133_244, w_041_494, w_090_001);
  and2 I133_249(w_133_249, w_059_181, w_015_353);
  or2  I133_290(w_133_290, w_105_229, w_068_101);
  not1 I133_313(w_133_313, w_069_245);
  nand2 I133_334(w_133_334, w_058_105, w_025_279);
  and2 I133_344(w_133_344, w_063_084, w_070_205);
  and2 I133_351(w_133_351, w_003_075, w_025_135);
  nand2 I133_362(w_133_362, w_098_001, w_060_285);
  not1 I133_368(w_133_368, w_006_005);
  or2  I133_373(w_133_373, w_037_036, w_009_625);
  or2  I133_374(w_133_374, w_105_386, w_087_040);
  or2  I133_376(w_133_376, w_058_208, w_019_011);
  or2  I133_378(w_133_378, w_001_011, w_059_242);
  not1 I134_001(w_134_001, w_114_197);
  or2  I134_002(w_134_002, w_086_081, w_069_038);
  and2 I134_017(w_134_017, w_114_194, w_128_496);
  not1 I134_018(w_134_018, w_073_219);
  or2  I134_066(w_134_066, w_009_314, w_024_178);
  not1 I134_071(w_134_071, w_129_048);
  nand2 I134_072(w_134_072, w_064_267, w_045_176);
  and2 I134_073(w_134_073, w_004_490, w_072_058);
  not1 I134_076(w_134_076, w_059_260);
  and2 I134_089(w_134_089, w_048_006, w_028_034);
  or2  I134_109(w_134_109, w_009_384, w_101_004);
  or2  I134_114(w_134_114, w_078_520, w_102_050);
  or2  I134_116(w_134_116, w_070_271, w_100_018);
  or2  I134_122(w_134_122, w_123_005, w_020_131);
  and2 I134_132(w_134_132, w_073_049, w_062_586);
  nand2 I134_135(w_134_135, w_081_021, w_090_543);
  not1 I134_138(w_134_138, w_019_007);
  nand2 I134_140(w_134_140, w_052_013, w_026_694);
  or2  I134_147(w_134_147, w_071_302, w_007_227);
  or2  I134_151(w_134_151, w_074_081, w_095_003);
  and2 I134_156(w_134_156, w_018_043, w_094_193);
  and2 I134_163(w_134_163, w_117_043, w_080_162);
  nand2 I134_169(w_134_169, w_099_053, w_126_187);
  not1 I134_173(w_134_173, w_081_008);
  not1 I134_185(w_134_185, w_052_014);
  and2 I134_200(w_134_200, w_098_041, w_041_359);
  nand2 I134_204(w_134_204, w_129_282, w_084_018);
  nand2 I134_218(w_134_218, w_094_344, w_020_067);
  or2  I134_230(w_134_230, w_082_166, w_115_194);
  or2  I134_251(w_134_251, w_104_109, w_086_028);
  not1 I134_256(w_134_256, w_074_012);
  nand2 I134_261(w_134_261, w_101_094, w_070_330);
  not1 I134_292(w_134_292, w_022_315);
  not1 I134_320(w_134_320, w_115_039);
  or2  I134_323(w_134_323, w_008_213, w_052_036);
  and2 I134_374(w_134_374, w_092_516, w_050_175);
  nand2 I134_375(w_134_375, w_012_121, w_121_126);
  not1 I134_396(w_134_396, w_093_208);
  nand2 I134_405(w_134_405, w_114_181, w_087_407);
  or2  I134_448(w_134_448, w_082_073, w_003_065);
  nand2 I134_451(w_134_451, w_002_471, w_037_032);
  or2  I134_474(w_134_474, w_062_264, w_077_500);
  or2  I134_488(w_134_490, w_134_489, w_125_242);
  or2  I134_489(w_134_491, w_134_490, w_097_526);
  and2 I134_490(w_134_492, w_134_491, w_133_099);
  nand2 I134_491(w_134_493, w_021_189, w_134_492);
  nand2 I134_492(w_134_494, w_134_493, w_047_225);
  nand2 I134_493(w_134_495, w_134_494, w_077_091);
  or2  I134_494(w_134_496, w_134_495, w_034_032);
  and2 I134_495(w_134_497, w_033_671, w_134_496);
  not1 I134_496(w_134_498, w_134_497);
  and2 I134_497(w_134_499, w_134_498, w_068_101);
  or2  I134_498(w_134_489, w_134_499, w_098_034);
  not1 I135_003(w_135_003, w_048_008);
  or2  I135_013(w_135_013, w_020_130, w_001_030);
  or2  I135_019(w_135_019, w_108_002, w_084_007);
  not1 I135_029(w_135_029, w_053_071);
  and2 I135_062(w_135_062, w_115_152, w_025_089);
  not1 I135_078(w_135_078, w_072_130);
  and2 I135_086(w_135_086, w_032_350, w_041_460);
  not1 I135_089(w_135_089, w_061_089);
  not1 I135_094(w_135_094, w_004_505);
  and2 I135_110(w_135_110, w_059_413, w_122_121);
  nand2 I135_111(w_135_111, w_071_075, w_057_131);
  and2 I135_119(w_135_119, w_118_061, w_131_223);
  nand2 I135_136(w_135_136, w_020_109, w_130_171);
  and2 I135_156(w_135_156, w_065_515, w_073_463);
  or2  I135_163(w_135_163, w_074_009, w_075_072);
  nand2 I135_164(w_135_164, w_077_043, w_027_165);
  nand2 I135_184(w_135_184, w_047_013, w_096_005);
  or2  I135_191(w_135_191, w_109_473, w_104_278);
  and2 I135_194(w_135_194, w_082_215, w_044_603);
  or2  I135_196(w_135_196, w_084_045, w_024_395);
  and2 I135_200(w_135_200, w_061_051, w_017_470);
  or2  I135_240(w_135_240, w_101_092, w_105_093);
  or2  I135_257(w_135_257, w_026_064, w_079_047);
  and2 I135_271(w_135_271, w_081_005, w_007_224);
  nand2 I135_286(w_135_286, w_012_333, w_036_440);
  or2  I135_348(w_135_348, w_005_135, w_086_190);
  or2  I135_354(w_135_354, w_036_028, w_037_086);
  nand2 I135_373(w_135_373, w_068_352, w_015_619);
  not1 I135_377(w_135_377, w_026_642);
  nand2 I135_398(w_135_398, w_090_469, w_067_196);
  or2  I135_429(w_135_429, w_044_705, w_073_634);
  or2  I135_438(w_135_438, w_127_069, w_026_598);
  or2  I135_457(w_135_457, w_027_127, w_086_181);
  and2 I135_487(w_135_487, w_032_346, w_047_197);
  not1 I135_488(w_135_488, w_040_340);
  not1 I135_528(w_135_528, w_112_068);
  nand2 I135_549(w_135_549, w_106_141, w_042_135);
  and2 I135_587(w_135_587, w_128_025, w_114_018);
  not1 I135_609(w_135_609, w_011_629);
  and2 I135_661(w_135_661, w_048_004, w_012_138);
  and2 I135_678(w_134_501, w_052_006, w_134_489);
  nand2 I136_002(w_136_002, w_003_015, w_021_100);
  or2  I136_004(w_136_004, w_096_005, w_112_174);
  nand2 I136_005(w_136_005, w_116_292, w_066_531);
  not1 I136_007(w_136_007, w_025_011);
  not1 I136_010(w_136_010, w_044_540);
  nand2 I136_011(w_136_011, w_012_028, w_104_357);
  and2 I136_013(w_136_013, w_001_011, w_072_047);
  and2 I136_014(w_136_014, w_105_268, w_064_058);
  and2 I136_017(w_136_017, w_109_293, w_088_018);
  not1 I136_020(w_136_020, w_035_021);
  or2  I136_024(w_136_024, w_014_054, w_030_044);
  and2 I136_025(w_136_025, w_023_053, w_008_307);
  and2 I136_030(w_136_030, w_132_330, w_041_581);
  nand2 I136_031(w_136_031, w_072_054, w_070_256);
  or2  I136_032(w_136_032, w_122_040, w_108_095);
  and2 I136_033(w_136_033, w_055_140, w_069_125);
  or2  I136_037(w_136_037, w_017_471, w_099_015);
  or2  I136_040(w_136_040, w_102_028, w_134_017);
  not1 I136_044(w_136_044, w_134_501);
  not1 I136_047(w_136_047, w_086_010);
  or2  I136_049(w_136_049, w_005_030, w_089_219);
  and2 I136_051(w_136_051, w_096_005, w_097_366);
  or2  I136_054(w_136_054, w_057_200, w_117_064);
  not1 I136_057(w_136_057, w_000_453);
  not1 I136_058(w_136_058, w_113_269);
  not1 I136_059(w_136_059, w_050_030);
  or2  I136_060(w_136_060, w_047_007, w_021_138);
  not1 I136_063(w_136_063, w_003_013);
  and2 I137_003(w_137_003, w_045_219, w_079_010);
  and2 I137_013(w_137_013, w_088_062, w_020_132);
  nand2 I137_017(w_137_017, w_035_048, w_050_359);
  nand2 I137_032(w_137_032, w_121_054, w_103_054);
  nand2 I137_034(w_137_034, w_098_004, w_030_328);
  nand2 I137_037(w_137_037, w_040_241, w_131_545);
  or2  I137_039(w_137_039, w_083_129, w_116_628);
  not1 I137_042(w_137_042, w_058_590);
  nand2 I137_045(w_137_045, w_015_049, w_105_268);
  not1 I137_061(w_137_061, w_103_113);
  or2  I137_075(w_137_075, w_058_660, w_044_286);
  and2 I137_076(w_137_076, w_064_233, w_031_017);
  nand2 I137_085(w_137_085, w_001_018, w_023_113);
  and2 I137_098(w_137_098, w_058_673, w_103_230);
  nand2 I137_099(w_137_099, w_054_256, w_055_207);
  nand2 I137_104(w_137_104, w_014_271, w_047_340);
  not1 I137_107(w_137_107, w_028_027);
  or2  I137_116(w_137_116, w_064_256, w_070_108);
  not1 I137_122(w_137_122, w_125_386);
  nand2 I137_123(w_137_123, w_035_061, w_089_232);
  or2  I137_146(w_137_146, w_118_062, w_010_488);
  not1 I137_162(w_137_162, w_136_025);
  and2 I137_164(w_137_164, w_052_028, w_026_693);
  or2  I137_176(w_137_176, w_074_193, w_080_138);
  or2  I137_183(w_137_183, w_096_005, w_127_061);
  nand2 I137_185(w_137_185, w_015_051, w_118_018);
  or2  I137_188(w_137_188, w_105_384, w_064_074);
  nand2 I137_190(w_137_190, w_075_067, w_048_000);
  nand2 I137_202(w_137_202, w_084_029, w_125_466);
  or2  I137_223(w_137_223, w_009_558, w_008_628);
  and2 I137_234(w_137_234, w_051_105, w_062_362);
  nand2 I137_235(w_137_235, w_017_124, w_047_014);
  or2  I137_255(w_137_255, w_105_235, w_114_003);
  and2 I137_266(w_137_266, w_062_027, w_081_017);
  nand2 I137_272(w_137_272, w_109_457, w_068_102);
  not1 I137_320(w_137_320, w_075_055);
  or2  I137_345(w_137_345, w_079_040, w_090_358);
  not1 I137_351(w_137_351, w_003_014);
  and2 I137_354(w_137_354, w_084_034, w_023_081);
  nand2 I137_356(w_137_356, w_004_162, w_065_031);
  or2  I137_443(w_137_443, w_069_260, w_001_008);
  not1 I137_464(w_137_464, w_071_312);
  and2 I137_469(w_137_469, w_084_018, w_099_123);
  or2  I137_473(w_137_473, w_071_093, w_013_359);
  not1 I138_023(w_138_023, w_015_584);
  or2  I138_024(w_138_024, w_132_082, w_128_025);
  not1 I138_037(w_138_037, w_132_130);
  and2 I138_047(w_138_047, w_102_060, w_096_002);
  nand2 I138_049(w_138_049, w_102_022, w_132_084);
  nand2 I138_051(w_138_051, w_088_050, w_061_285);
  not1 I138_056(w_138_056, w_095_012);
  or2  I138_058(w_138_058, w_119_007, w_035_037);
  or2  I138_060(w_138_060, w_118_010, w_119_040);
  or2  I138_061(w_138_061, w_114_009, w_113_158);
  nand2 I138_066(w_138_066, w_001_013, w_107_180);
  and2 I138_067(w_138_067, w_022_140, w_045_270);
  and2 I138_069(w_138_069, w_001_022, w_125_208);
  nand2 I138_073(w_138_073, w_080_076, w_031_205);
  and2 I138_078(w_138_078, w_029_027, w_022_249);
  not1 I138_083(w_138_083, w_059_213);
  and2 I138_093(w_138_093, w_120_135, w_076_221);
  or2  I138_094(w_138_094, w_002_392, w_010_373);
  not1 I138_096(w_138_096, w_003_002);
  not1 I138_100(w_138_100, w_006_120);
  nand2 I138_104(w_138_104, w_030_194, w_116_510);
  and2 I138_120(w_138_120, w_117_036, w_061_200);
  or2  I138_125(w_138_125, w_063_090, w_052_020);
  nand2 I138_134(w_138_134, w_137_234, w_135_164);
  nand2 I138_157(w_138_157, w_056_465, w_135_373);
  not1 I138_160(w_138_160, w_016_006);
  and2 I138_168(w_138_168, w_106_139, w_134_169);
  and2 I138_171(w_138_171, w_029_073, w_067_390);
  not1 I138_192(w_138_192, w_002_418);
  or2  I138_205(w_138_205, w_104_256, w_093_390);
  nand2 I138_206(w_138_206, w_112_035, w_053_109);
  nand2 I138_214(w_138_214, w_093_177, w_065_095);
  and2 I138_221(w_138_221, w_079_001, w_009_361);
  or2  I138_231(w_138_231, w_121_106, w_078_037);
  nand2 I138_238(w_138_238, w_074_141, w_085_015);
  nand2 I138_241(w_138_241, w_000_043, w_039_351);
  and2 I138_246(w_138_246, w_109_028, w_104_179);
  or2  I138_248(w_138_248, w_047_099, w_109_350);
  and2 I138_250(w_138_250, w_092_107, w_099_163);
  and2 I138_258(w_138_258, w_041_507, w_094_222);
  not1 I138_261(w_138_261, w_074_005);
  not1 I138_282(w_138_282, w_098_045);
  or2  I138_283(w_138_283, w_075_100, w_126_017);
  nand2 I138_304(w_138_304, w_113_276, w_084_047);
  and2 I138_308(w_138_308, w_129_210, w_039_055);
  nand2 I138_309(w_138_309, w_076_060, w_123_304);
  and2 I138_310(w_138_310, w_106_076, w_092_360);
  or2  I138_326(w_138_326, w_077_209, w_062_259);
  not1 I139_001(w_139_001, w_101_284);
  nand2 I139_002(w_139_002, w_044_694, w_061_217);
  not1 I139_004(w_139_004, w_138_282);
  not1 I139_005(w_139_005, w_062_330);
  nand2 I139_006(w_139_006, w_053_129, w_061_260);
  or2  I139_007(w_139_007, w_013_515, w_121_086);
  nand2 I139_009(w_139_009, w_126_127, w_087_120);
  or2  I139_010(w_139_010, w_074_313, w_080_269);
  nand2 I139_011(w_139_011, w_128_103, w_016_006);
  and2 I139_013(w_139_013, w_018_032, w_005_236);
  not1 I139_014(w_139_014, w_076_070);
  not1 I139_015(w_139_015, w_108_085);
  not1 I139_016(w_139_016, w_095_027);
  or2  I139_018(w_139_018, w_003_002, w_003_009);
  nand2 I139_019(w_139_019, w_104_131, w_057_066);
  nand2 I139_020(w_139_020, w_060_167, w_126_090);
  or2  I139_021(w_139_021, w_037_262, w_133_368);
  or2  I139_022(w_139_022, w_013_042, w_044_375);
  and2 I139_023(w_139_023, w_056_008, w_121_048);
  nand2 I139_024(w_139_024, w_135_094, w_125_124);
  or2  I139_025(w_139_025, w_101_122, w_005_282);
  and2 I139_026(w_139_026, w_114_065, w_046_620);
  not1 I139_027(w_139_027, w_013_155);
  and2 I140_001(w_140_001, w_138_049, w_031_446);
  or2  I140_009(w_140_009, w_116_554, w_138_241);
  or2  I140_010(w_140_010, w_054_533, w_139_022);
  and2 I140_015(w_140_015, w_094_444, w_058_593);
  and2 I140_020(w_140_020, w_128_091, w_027_124);
  not1 I140_021(w_140_021, w_023_032);
  not1 I140_024(w_140_024, w_099_159);
  and2 I140_027(w_140_027, w_053_132, w_137_098);
  nand2 I140_031(w_140_031, w_131_303, w_030_125);
  and2 I140_036(w_140_036, w_108_031, w_031_343);
  and2 I140_042(w_140_042, w_095_055, w_115_084);
  nand2 I140_052(w_140_052, w_028_117, w_017_538);
  or2  I140_062(w_140_062, w_116_008, w_098_071);
  or2  I140_068(w_140_068, w_048_015, w_054_456);
  and2 I140_071(w_140_071, w_037_315, w_130_089);
  and2 I140_073(w_140_073, w_032_172, w_093_217);
  and2 I140_074(w_140_074, w_031_128, w_129_034);
  nand2 I140_088(w_140_088, w_030_057, w_111_070);
  and2 I140_092(w_140_092, w_049_303, w_128_234);
  or2  I140_093(w_140_093, w_103_228, w_007_233);
  or2  I140_094(w_140_094, w_022_303, w_107_159);
  nand2 I140_096(w_140_096, w_121_106, w_031_058);
  not1 I140_137(w_140_137, w_079_029);
  and2 I140_155(w_140_155, w_022_341, w_127_038);
  nand2 I140_161(w_140_161, w_075_052, w_127_004);
  nand2 I140_165(w_140_165, w_053_072, w_028_151);
  not1 I140_176(w_140_176, w_132_305);
  nand2 I140_178(w_140_178, w_044_341, w_035_025);
  nand2 I140_180(w_140_180, w_040_423, w_082_299);
  and2 I140_184(w_140_184, w_018_012, w_081_001);
  nand2 I140_188(w_140_188, w_107_054, w_047_136);
  not1 I140_189(w_140_189, w_108_197);
  not1 I140_190(w_140_190, w_121_168);
  and2 I140_202(w_140_202, w_018_036, w_037_077);
  nand2 I140_216(w_140_216, w_046_059, w_032_295);
  and2 I140_230(w_140_230, w_132_255, w_071_247);
  not1 I140_233(w_140_233, w_047_045);
  and2 I140_234(w_140_234, w_046_526, w_128_329);
  and2 I140_241(w_140_243, w_140_242, w_062_125);
  nand2 I140_242(w_140_244, w_140_256, w_140_243);
  not1 I140_243(w_140_245, w_140_244);
  not1 I140_244(w_140_246, w_140_245);
  and2 I140_245(w_140_247, w_140_246, w_013_251);
  or2  I140_246(w_140_242, w_140_247, w_054_051);
  or2  I140_247(w_140_252, w_102_274, w_140_251);
  and2 I140_248(w_140_253, w_140_252, w_094_246);
  and2 I140_249(w_140_254, w_140_253, w_052_037);
  not1 I140_250(w_140_251, w_140_244);
  and2 I140_251(w_140_256, w_043_035, w_140_254);
  not1 I141_000(w_141_000, w_061_023);
  not1 I141_002(w_141_002, w_003_001);
  not1 I141_008(w_141_008, w_070_173);
  or2  I141_011(w_141_011, w_042_276, w_089_269);
  and2 I141_012(w_141_012, w_110_210, w_041_338);
  and2 I141_016(w_141_016, w_040_246, w_003_003);
  nand2 I141_018(w_141_018, w_015_095, w_068_139);
  nand2 I141_021(w_141_021, w_081_022, w_110_358);
  or2  I141_044(w_141_044, w_117_011, w_042_268);
  not1 I141_048(w_141_048, w_079_005);
  or2  I141_050(w_141_050, w_075_074, w_057_008);
  or2  I141_053(w_141_053, w_121_088, w_120_008);
  and2 I141_056(w_141_056, w_057_117, w_019_014);
  not1 I141_059(w_141_059, w_098_050);
  not1 I141_065(w_141_065, w_010_429);
  not1 I141_068(w_141_068, w_124_104);
  and2 I141_079(w_141_079, w_063_024, w_016_000);
  and2 I141_093(w_141_093, w_041_102, w_065_043);
  or2  I141_107(w_141_107, w_025_064, w_045_075);
  not1 I141_114(w_141_114, w_082_167);
  or2  I141_117(w_141_117, w_138_060, w_098_013);
  nand2 I141_128(w_141_128, w_042_109, w_121_047);
  nand2 I141_133(w_141_133, w_120_666, w_109_280);
  nand2 I141_139(w_141_139, w_084_023, w_050_367);
  not1 I141_143(w_141_143, w_129_289);
  and2 I141_149(w_141_149, w_009_268, w_063_376);
  nand2 I141_151(w_141_151, w_058_493, w_085_028);
  not1 I141_154(w_141_154, w_075_009);
  nand2 I141_168(w_141_168, w_062_060, w_014_226);
  not1 I141_171(w_141_171, w_057_117);
  or2  I141_175(w_141_175, w_094_522, w_125_187);
  nand2 I141_176(w_141_176, w_119_117, w_078_429);
  not1 I142_040(w_142_040, w_099_088);
  nand2 I142_076(w_142_076, w_095_055, w_127_071);
  or2  I142_095(w_142_095, w_072_295, w_035_064);
  not1 I142_101(w_142_101, w_016_003);
  and2 I142_129(w_142_129, w_141_065, w_040_539);
  nand2 I142_147(w_142_147, w_124_287, w_083_135);
  and2 I142_181(w_142_181, w_016_005, w_089_128);
  and2 I142_187(w_142_187, w_139_002, w_119_085);
  and2 I142_205(w_142_205, w_027_171, w_016_005);
  and2 I142_209(w_142_209, w_127_065, w_053_137);
  not1 I142_212(w_142_212, w_008_637);
  nand2 I142_258(w_142_258, w_010_570, w_116_530);
  not1 I142_276(w_142_276, w_021_024);
  nand2 I142_303(w_142_303, w_005_032, w_082_314);
  or2  I142_321(w_142_321, w_086_073, w_005_198);
  and2 I142_348(w_142_348, w_011_406, w_111_046);
  not1 I142_365(w_142_365, w_101_207);
  nand2 I142_421(w_142_421, w_075_011, w_012_253);
  or2  I142_442(w_142_442, w_130_075, w_069_060);
  and2 I142_494(w_142_494, w_011_328, w_077_048);
  not1 I142_499(w_142_499, w_007_004);
  or2  I142_503(w_142_503, w_075_138, w_090_487);
  or2  I142_517(w_142_517, w_102_193, w_072_058);
  and2 I142_559(w_142_559, w_028_105, w_011_127);
  or2  I142_587(w_142_587, w_128_464, w_132_331);
  nand2 I142_603(w_142_603, w_074_168, w_021_064);
  not1 I142_607(w_142_607, w_127_007);
  not1 I142_638(w_142_638, w_041_128);
  or2  I142_772(w_142_772, w_120_215, w_021_190);
  not1 I142_777(w_142_777, w_105_130);
  nand2 I142_792(w_142_792, w_064_056, w_004_227);
  and2 I143_000(w_143_000, w_089_156, w_049_252);
  not1 I143_004(w_143_004, w_100_036);
  not1 I143_014(w_143_014, w_112_160);
  not1 I143_018(w_143_018, w_063_066);
  not1 I143_019(w_143_019, w_045_255);
  not1 I143_044(w_143_044, w_086_161);
  and2 I143_061(w_143_061, w_125_030, w_140_180);
  or2  I143_066(w_143_066, w_078_080, w_043_027);
  not1 I143_068(w_143_068, w_115_016);
  or2  I143_076(w_143_076, w_012_272, w_120_674);
  and2 I143_081(w_143_081, w_112_077, w_037_031);
  or2  I143_082(w_143_082, w_068_042, w_110_148);
  nand2 I143_088(w_143_088, w_112_065, w_016_000);
  and2 I143_090(w_143_090, w_133_134, w_117_008);
  nand2 I143_106(w_143_106, w_009_449, w_014_131);
  and2 I143_107(w_143_107, w_130_375, w_120_410);
  not1 I143_111(w_143_111, w_036_215);
  and2 I143_116(w_143_116, w_060_073, w_124_091);
  or2  I143_209(w_143_209, w_000_218, w_045_400);
  nand2 I143_211(w_143_211, w_082_040, w_011_303);
  nand2 I143_243(w_143_243, w_091_030, w_120_140);
  not1 I143_257(w_143_257, w_000_245);
  nand2 I143_265(w_143_265, w_001_015, w_014_189);
  and2 I143_300(w_143_300, w_080_013, w_053_006);
  or2  I143_344(w_143_344, w_072_096, w_026_061);
  nand2 I143_353(w_143_353, w_087_293, w_067_275);
  nand2 I143_374(w_143_374, w_062_535, w_071_001);
  or2  I143_401(w_143_401, w_101_253, w_113_234);
  or2  I143_408(w_143_408, w_011_243, w_036_188);
  not1 I143_473(w_143_473, w_109_474);
  and2 I143_479(w_143_479, w_048_016, w_002_189);
  not1 I143_493(w_143_493, w_023_101);
  and2 I143_501(w_143_501, w_094_052, w_010_145);
  not1 I143_530(w_143_530, w_141_133);
  nand2 I143_535(w_143_535, w_133_066, w_052_009);
  not1 I143_554(w_143_554, w_049_093);
  and2 I143_568(w_143_568, w_014_192, w_083_183);
  nand2 I143_575(w_143_575, w_130_499, w_101_098);
  nand2 I143_581(w_143_581, w_075_013, w_116_150);
  and2 I143_598(w_143_598, w_131_269, w_041_434);
  nand2 I143_652(w_143_652, w_023_129, w_136_010);
  nand2 I144_006(w_144_006, w_041_491, w_050_027);
  or2  I144_010(w_144_010, w_006_054, w_084_000);
  not1 I144_032(w_144_032, w_104_263);
  not1 I144_035(w_144_035, w_120_674);
  not1 I144_043(w_144_043, w_023_184);
  or2  I144_044(w_144_044, w_013_439, w_054_332);
  or2  I144_045(w_144_045, w_032_177, w_076_197);
  not1 I144_061(w_144_061, w_086_101);
  not1 I144_062(w_144_062, w_071_026);
  or2  I144_077(w_144_077, w_130_418, w_111_054);
  not1 I144_079(w_144_079, w_128_021);
  not1 I144_105(w_144_105, w_049_184);
  nand2 I144_125(w_144_125, w_031_090, w_009_412);
  not1 I144_142(w_144_142, w_101_143);
  or2  I144_169(w_144_169, w_055_127, w_068_323);
  not1 I144_173(w_144_173, w_046_201);
  not1 I144_182(w_144_182, w_076_200);
  nand2 I144_185(w_144_185, w_117_062, w_107_091);
  nand2 I144_186(w_144_186, w_043_012, w_032_410);
  and2 I144_190(w_144_190, w_125_191, w_017_112);
  not1 I144_193(w_144_193, w_141_068);
  or2  I144_202(w_144_202, w_011_143, w_122_084);
  not1 I144_206(w_144_206, w_094_363);
  and2 I144_219(w_144_219, w_028_134, w_053_047);
  or2  I144_228(w_144_228, w_030_112, w_027_086);
  or2  I144_242(w_144_242, w_062_259, w_105_386);
  nand2 I144_302(w_144_302, w_133_095, w_055_225);
  nand2 I144_306(w_144_306, w_026_139, w_087_134);
  nand2 I144_309(w_144_309, w_142_503, w_030_191);
  nand2 I144_346(w_144_346, w_010_663, w_010_074);
  not1 I144_373(w_144_373, w_091_169);
  or2  I144_406(w_144_406, w_121_210, w_063_415);
  or2  I144_447(w_144_447, w_053_072, w_031_138);
  or2  I144_473(w_144_473, w_110_171, w_084_023);
  and2 I144_557(w_144_559, w_049_026, w_144_558);
  not1 I144_558(w_144_560, w_144_559);
  and2 I144_559(w_144_561, w_079_030, w_144_560);
  and2 I144_560(w_144_562, w_144_561, w_129_029);
  not1 I144_561(w_144_563, w_144_562);
  not1 I144_562(w_144_564, w_144_563);
  and2 I144_563(w_144_565, w_144_564, w_069_077);
  not1 I144_564(w_144_558, w_144_565);
  not1 I145_002(w_145_002, w_087_323);
  nand2 I145_005(w_145_005, w_068_295, w_072_017);
  and2 I145_011(w_145_011, w_006_060, w_089_190);
  nand2 I145_012(w_145_012, w_039_187, w_012_006);
  or2  I145_016(w_145_016, w_075_147, w_136_030);
  not1 I145_020(w_145_020, w_018_011);
  nand2 I145_022(w_145_022, w_073_717, w_036_271);
  not1 I145_027(w_145_027, w_013_501);
  nand2 I145_030(w_145_030, w_092_112, w_011_500);
  or2  I145_032(w_145_032, w_137_473, w_020_025);
  not1 I145_035(w_145_035, w_035_092);
  nand2 I145_037(w_145_037, w_108_003, w_080_080);
  nand2 I145_038(w_145_038, w_081_021, w_134_132);
  not1 I145_039(w_145_039, w_126_158);
  or2  I145_040(w_145_040, w_032_084, w_019_001);
  nand2 I145_046(w_145_046, w_005_092, w_012_076);
  nand2 I145_048(w_145_048, w_017_165, w_131_450);
  and2 I145_052(w_145_052, w_064_055, w_050_007);
  nand2 I145_066(w_145_066, w_127_031, w_069_067);
  or2  I145_068(w_145_068, w_069_202, w_045_353);
  or2  I145_070(w_145_070, w_092_225, w_046_677);
  or2  I145_075(w_145_075, w_143_473, w_128_073);
  or2  I145_077(w_145_077, w_029_086, w_059_173);
  and2 I145_079(w_145_079, w_081_003, w_033_486);
  or2  I146_001(w_146_001, w_018_022, w_018_037);
  nand2 I146_005(w_146_005, w_112_172, w_011_288);
  nand2 I146_008(w_146_008, w_029_050, w_005_191);
  not1 I146_036(w_146_036, w_075_058);
  and2 I146_042(w_146_042, w_002_190, w_058_258);
  nand2 I146_044(w_146_044, w_059_255, w_120_311);
  and2 I146_049(w_146_049, w_053_031, w_134_375);
  or2  I146_057(w_146_057, w_005_028, w_048_007);
  and2 I146_071(w_146_071, w_129_149, w_035_088);
  and2 I146_079(w_146_079, w_013_208, w_071_227);
  and2 I146_085(w_146_085, w_036_024, w_109_152);
  and2 I146_088(w_146_088, w_056_348, w_043_012);
  and2 I146_090(w_146_090, w_114_056, w_145_040);
  and2 I146_092(w_146_092, w_086_192, w_023_210);
  and2 I146_107(w_146_107, w_133_351, w_020_044);
  not1 I146_124(w_146_124, w_124_027);
  or2  I146_133(w_146_133, w_097_180, w_092_492);
  not1 I146_142(w_146_142, w_031_253);
  nand2 I146_168(w_146_168, w_100_007, w_121_082);
  nand2 I146_182(w_146_182, w_130_278, w_068_060);
  or2  I146_191(w_146_191, w_088_029, w_137_356);
  not1 I146_198(w_146_198, w_040_497);
  and2 I146_210(w_146_210, w_060_024, w_095_034);
  or2  I146_213(w_146_213, w_053_053, w_124_232);
  and2 I146_227(w_146_227, w_106_084, w_065_058);
  and2 I146_255(w_146_255, w_006_116, w_101_095);
  not1 I146_256(w_146_256, w_020_209);
  not1 I146_273(w_146_273, w_062_355);
  and2 I146_275(w_146_275, w_132_089, w_118_005);
  and2 I146_279(w_146_279, w_052_026, w_056_254);
  not1 I146_285(w_146_285, w_017_159);
  not1 I146_291(w_146_291, w_101_008);
  or2  I146_297(w_146_297, w_028_086, w_128_524);
  not1 I146_302(w_146_302, w_003_000);
  not1 I146_303(w_146_303, w_079_062);
  not1 I146_305(w_146_305, w_013_178);
  nand2 I146_309(w_146_309, w_038_176, w_137_037);
  not1 I146_311(w_146_311, w_038_600);
  and2 I146_320(w_146_320, w_028_170, w_089_164);
  not1 I146_321(w_146_321, w_012_215);
  and2 I146_323(w_146_323, w_054_276, w_048_017);
  not1 I146_324(w_146_324, w_050_131);
  nand2 I147_003(w_147_003, w_050_082, w_080_481);
  nand2 I147_007(w_147_007, w_116_414, w_070_004);
  or2  I147_020(w_147_020, w_046_575, w_091_037);
  or2  I147_022(w_147_022, w_071_102, w_143_575);
  or2  I147_027(w_147_027, w_091_105, w_104_193);
  nand2 I147_029(w_147_029, w_069_117, w_131_121);
  and2 I147_031(w_147_031, w_107_292, w_030_055);
  nand2 I147_032(w_147_032, w_069_185, w_010_669);
  and2 I147_037(w_147_037, w_032_173, w_124_220);
  or2  I147_040(w_147_040, w_008_562, w_018_009);
  nand2 I147_050(w_147_050, w_128_297, w_111_081);
  or2  I147_061(w_147_061, w_113_174, w_102_133);
  or2  I147_062(w_147_062, w_102_529, w_109_327);
  or2  I147_063(w_147_063, w_022_120, w_004_051);
  or2  I147_077(w_147_077, w_102_097, w_058_469);
  or2  I147_089(w_147_089, w_093_119, w_024_073);
  nand2 I147_097(w_147_097, w_091_014, w_050_534);
  nand2 I147_099(w_147_099, w_136_017, w_077_039);
  not1 I147_100(w_147_100, w_054_077);
  or2  I147_113(w_147_113, w_061_426, w_076_218);
  not1 I147_116(w_147_116, w_119_083);
  nand2 I147_118(w_147_118, w_040_367, w_083_166);
  and2 I147_146(w_147_146, w_094_064, w_058_402);
  not1 I147_147(w_147_147, w_128_139);
  not1 I147_160(w_147_160, w_048_005);
  and2 I147_162(w_147_162, w_127_035, w_102_589);
  and2 I147_165(w_147_165, w_019_017, w_075_148);
  nand2 I147_166(w_147_166, w_078_044, w_039_263);
  nand2 I147_168(w_147_168, w_047_287, w_063_267);
  not1 I147_173(w_147_173, w_123_162);
  or2  I147_175(w_147_175, w_111_023, w_097_063);
  nand2 I147_202(w_147_202, w_044_344, w_026_595);
  and2 I147_203(w_147_203, w_129_005, w_105_097);
  and2 I147_214(w_147_214, w_065_582, w_137_039);
  not1 I147_216(w_147_216, w_099_136);
  or2  I147_226(w_147_226, w_104_213, w_116_112);
  nand2 I148_004(w_148_004, w_022_204, w_059_695);
  nand2 I148_010(w_148_010, w_112_008, w_064_140);
  or2  I148_015(w_148_015, w_113_050, w_147_113);
  or2  I148_017(w_148_017, w_089_166, w_004_379);
  or2  I148_038(w_148_038, w_100_092, w_022_090);
  not1 I148_043(w_148_043, w_114_117);
  nand2 I148_060(w_148_060, w_147_147, w_120_353);
  nand2 I148_077(w_148_077, w_138_258, w_087_273);
  nand2 I148_085(w_148_085, w_135_348, w_082_487);
  and2 I148_087(w_148_087, w_110_196, w_012_098);
  not1 I148_106(w_148_106, w_012_262);
  and2 I148_123(w_148_123, w_111_008, w_111_047);
  not1 I148_164(w_148_164, w_046_551);
  or2  I148_209(w_148_209, w_129_182, w_133_061);
  nand2 I148_215(w_148_215, w_112_173, w_055_197);
  and2 I148_241(w_148_241, w_114_036, w_119_143);
  and2 I148_279(w_148_279, w_039_571, w_035_070);
  and2 I148_283(w_148_283, w_142_212, w_081_021);
  or2  I148_286(w_148_286, w_108_161, w_099_003);
  and2 I148_353(w_148_353, w_002_445, w_025_121);
  nand2 I148_371(w_148_371, w_054_194, w_009_059);
  nand2 I148_375(w_148_375, w_096_002, w_011_057);
  or2  I148_398(w_148_398, w_106_141, w_140_234);
  or2  I148_417(w_148_417, w_142_276, w_031_340);
  or2  I148_447(w_148_447, w_062_606, w_141_048);
  or2  I148_499(w_148_499, w_135_271, w_000_456);
  nand2 I148_528(w_148_528, w_093_458, w_037_002);
  nand2 I148_536(w_148_536, w_012_231, w_036_192);
  not1 I148_553(w_148_553, w_033_372);
  and2 I148_565(w_148_565, w_030_316, w_054_071);
  nand2 I148_574(w_148_574, w_096_000, w_087_207);
  and2 I148_576(w_148_576, w_071_063, w_089_025);
  or2  I148_581(w_148_581, w_036_294, w_108_015);
  and2 I148_595(w_148_595, w_053_054, w_046_255);
  or2  I148_609(w_148_609, w_071_257, w_034_046);
  not1 I148_611(w_148_611, w_061_287);
  not1 I148_650(w_148_650, w_122_017);
  not1 I148_670(w_148_670, w_003_058);
  not1 I148_684(w_148_684, w_093_128);
  not1 I148_688(w_148_690, w_148_689);
  and2 I148_689(w_148_691, w_079_004, w_148_690);
  nand2 I148_690(w_148_692, w_148_705, w_148_691);
  nand2 I148_691(w_148_693, w_148_692, w_139_007);
  and2 I148_692(w_148_694, w_148_693, w_050_344);
  or2  I148_693(w_148_689, w_148_694, w_040_361);
  not1 I148_694(w_148_699, w_148_698);
  not1 I148_695(w_148_700, w_148_699);
  nand2 I148_696(w_148_701, w_148_700, w_078_229);
  or2  I148_697(w_148_702, w_148_701, w_093_448);
  and2 I148_698(w_148_703, w_025_240, w_148_702);
  not1 I148_699(w_148_698, w_148_692);
  and2 I148_700(w_148_705, w_003_070, w_148_703);
  not1 I148_701(w_148_708, w_148_707);
  or2  I148_702(w_148_709, w_042_311, w_148_708);
  and2 I148_703(w_148_710, w_148_709, w_024_558);
  and2 I148_704(w_148_711, w_089_042, w_148_710);
  not1 I148_705(w_148_712, w_148_711);
  and2 I148_706(w_148_713, w_148_712, w_132_180);
  nand2 I148_707(w_148_707, w_148_721, w_148_713);
  or2  I148_708(w_148_718, w_135_354, w_148_717);
  and2 I148_709(w_148_719, w_106_050, w_148_718);
  not1 I148_710(w_148_717, w_148_707);
  and2 I148_711(w_148_721, w_092_189, w_148_719);
  not1 I149_004(w_149_004, w_007_291);
  or2  I149_015(w_149_015, w_142_076, w_126_082);
  and2 I149_018(w_149_018, w_015_235, w_106_183);
  nand2 I149_027(w_149_027, w_070_021, w_077_601);
  nand2 I149_032(w_149_032, w_137_107, w_143_243);
  or2  I149_041(w_149_041, w_000_733, w_096_005);
  not1 I149_056(w_149_056, w_089_025);
  and2 I149_060(w_149_060, w_071_099, w_002_366);
  or2  I149_063(w_149_063, w_065_386, w_128_187);
  not1 I149_075(w_149_075, w_041_439);
  nand2 I149_079(w_149_079, w_137_017, w_132_406);
  nand2 I149_080(w_149_080, w_093_143, w_064_143);
  and2 I149_081(w_149_081, w_015_343, w_064_086);
  nand2 I149_082(w_149_082, w_117_017, w_131_053);
  nand2 I149_126(w_149_126, w_067_290, w_004_075);
  or2  I149_138(w_149_138, w_094_173, w_044_740);
  and2 I149_159(w_149_159, w_041_618, w_103_145);
  and2 I149_179(w_149_179, w_101_266, w_039_383);
  not1 I149_207(w_149_207, w_067_270);
  not1 I149_261(w_149_261, w_102_476);
  and2 I149_302(w_149_302, w_130_295, w_019_002);
  and2 I149_314(w_149_314, w_081_003, w_090_206);
  not1 I149_364(w_149_364, w_014_058);
  or2  I149_367(w_149_367, w_110_246, w_068_084);
  not1 I149_368(w_149_368, w_096_003);
  or2  I149_430(w_149_430, w_146_279, w_094_546);
  or2  I149_438(w_149_438, w_009_184, w_001_029);
  or2  I149_450(w_149_450, w_062_013, w_058_335);
  nand2 I149_466(w_149_466, w_140_230, w_077_488);
  or2  I149_478(w_149_478, w_071_000, w_064_070);
  not1 I149_484(w_149_484, w_088_066);
  or2  I149_501(w_149_501, w_096_002, w_004_230);
  and2 I149_506(w_149_506, w_082_148, w_068_246);
  nand2 I149_517(w_149_517, w_045_043, w_092_412);
  or2  I149_590(w_149_590, w_095_053, w_128_640);
  and2 I149_600(w_149_600, w_043_029, w_078_024);
  or2  I149_612(w_149_612, w_101_283, w_029_002);
  not1 I149_619(w_149_619, w_008_638);
  or2  I149_631(w_149_631, w_140_036, w_110_250);
  or2  I149_636(w_149_636, w_059_636, w_049_338);
  or2  I150_000(w_150_000, w_038_265, w_013_208);
  and2 I150_003(w_150_003, w_085_016, w_140_176);
  and2 I150_008(w_150_008, w_003_044, w_016_001);
  nand2 I150_009(w_150_009, w_146_198, w_084_038);
  not1 I150_041(w_150_041, w_038_032);
  and2 I150_056(w_150_056, w_100_022, w_050_072);
  not1 I150_067(w_150_067, w_112_127);
  and2 I150_068(w_150_068, w_088_094, w_043_004);
  and2 I150_108(w_150_108, w_127_043, w_078_055);
  not1 I150_127(w_150_127, w_013_184);
  or2  I150_150(w_150_150, w_083_154, w_128_414);
  and2 I150_159(w_150_159, w_033_024, w_022_295);
  not1 I150_182(w_150_182, w_125_439);
  and2 I150_191(w_150_191, w_109_363, w_144_193);
  or2  I150_197(w_150_197, w_122_120, w_105_132);
  and2 I150_200(w_150_200, w_050_416, w_063_176);
  not1 I150_231(w_150_231, w_132_229);
  nand2 I150_239(w_150_239, w_042_117, w_115_136);
  or2  I150_241(w_150_241, w_067_007, w_031_543);
  or2  I150_253(w_150_253, w_114_119, w_012_275);
  nand2 I150_274(w_150_274, w_010_312, w_030_236);
  or2  I150_294(w_150_294, w_103_016, w_078_013);
  and2 I150_296(w_150_296, w_087_015, w_086_078);
  nand2 I150_300(w_150_300, w_082_338, w_040_667);
  and2 I150_318(w_150_318, w_058_310, w_061_465);
  not1 I150_324(w_150_324, w_012_316);
  or2  I150_333(w_150_333, w_040_555, w_036_273);
  not1 I150_334(w_150_334, w_097_303);
  and2 I150_345(w_150_345, w_009_470, w_149_368);
  or2  I150_361(w_150_361, w_004_069, w_032_085);
  not1 I150_363(w_150_363, w_075_025);
  and2 I150_378(w_150_378, w_008_550, w_121_112);
  not1 I150_393(w_150_393, w_119_040);
  not1 I150_394(w_150_394, w_023_191);
  not1 I150_449(w_150_449, w_134_320);
  nand2 I151_009(w_151_009, w_150_363, w_105_102);
  and2 I151_011(w_151_011, w_062_316, w_038_299);
  nand2 I151_013(w_151_013, w_056_039, w_025_094);
  and2 I151_034(w_151_034, w_103_168, w_047_126);
  and2 I151_048(w_151_048, w_043_011, w_026_692);
  not1 I151_057(w_151_057, w_030_069);
  nand2 I151_068(w_151_068, w_066_625, w_055_337);
  and2 I151_080(w_151_080, w_088_125, w_081_017);
  nand2 I151_086(w_151_086, w_071_267, w_011_565);
  not1 I151_088(w_151_088, w_097_125);
  and2 I151_099(w_151_099, w_043_023, w_077_185);
  or2  I151_108(w_151_108, w_020_001, w_122_074);
  and2 I151_116(w_151_116, w_021_182, w_078_441);
  nand2 I151_130(w_151_130, w_082_463, w_140_184);
  or2  I151_148(w_151_148, w_109_392, w_009_054);
  not1 I151_156(w_151_156, w_104_366);
  not1 I151_160(w_151_160, w_133_376);
  not1 I151_175(w_151_175, w_080_213);
  not1 I151_178(w_151_178, w_075_039);
  not1 I151_184(w_151_184, w_106_058);
  nand2 I151_200(w_151_200, w_067_165, w_007_062);
  and2 I151_203(w_151_203, w_144_309, w_076_136);
  nand2 I151_208(w_151_208, w_022_141, w_125_347);
  or2  I151_215(w_151_215, w_065_543, w_039_446);
  nand2 I151_222(w_151_222, w_129_305, w_024_571);
  and2 I151_247(w_151_247, w_136_037, w_088_005);
  not1 I151_259(w_151_259, w_073_675);
  or2  I151_262(w_151_262, w_041_336, w_149_517);
  not1 I151_264(w_151_264, w_091_112);
  and2 I151_268(w_151_268, w_084_040, w_000_703);
  or2  I151_276(w_151_276, w_025_168, w_033_695);
  and2 I151_284(w_151_284, w_033_617, w_133_097);
  nand2 I151_295(w_151_295, w_118_070, w_010_571);
  and2 I151_302(w_151_302, w_081_018, w_148_283);
  or2  I151_321(w_151_321, w_089_012, w_125_417);
  and2 I151_352(w_151_352, w_012_076, w_143_493);
  nand2 I151_366(w_151_366, w_077_401, w_009_058);
  nand2 I151_367(w_151_367, w_106_204, w_131_486);
  not1 I151_388(w_151_388, w_116_042);
  not1 I151_453(w_151_453, w_051_166);
  or2  I152_002(w_152_002, w_079_002, w_047_007);
  not1 I152_007(w_152_007, w_148_574);
  nand2 I152_008(w_152_008, w_042_123, w_108_065);
  and2 I152_045(w_152_045, w_127_048, w_084_015);
  not1 I152_073(w_152_073, w_103_006);
  and2 I152_089(w_152_089, w_107_415, w_096_002);
  and2 I152_108(w_152_108, w_106_165, w_080_118);
  and2 I152_118(w_152_118, w_126_073, w_058_513);
  or2  I152_153(w_152_153, w_034_024, w_001_009);
  not1 I152_161(w_152_161, w_099_093);
  not1 I152_167(w_152_167, w_062_768);
  nand2 I152_198(w_152_198, w_080_044, w_102_123);
  and2 I152_200(w_152_200, w_044_289, w_146_092);
  nand2 I152_221(w_152_221, w_050_226, w_080_251);
  not1 I152_234(w_152_234, w_014_130);
  and2 I152_236(w_152_236, w_114_131, w_116_545);
  not1 I152_337(w_152_337, w_095_038);
  nand2 I152_348(w_152_348, w_143_265, w_100_127);
  nand2 I152_387(w_152_387, w_084_046, w_124_112);
  not1 I152_428(w_152_428, w_010_770);
  nand2 I152_468(w_152_468, w_071_143, w_086_264);
  nand2 I152_511(w_152_511, w_076_351, w_086_033);
  and2 I152_513(w_152_513, w_094_534, w_130_184);
  and2 I152_573(w_152_573, w_013_358, w_025_227);
  nand2 I152_586(w_152_586, w_065_316, w_077_107);
  and2 I152_601(w_152_601, w_126_056, w_144_032);
  not1 I152_621(w_152_621, w_105_120);
  or2  I152_714(w_152_714, w_055_072, w_094_116);
  not1 I152_721(w_152_721, w_097_038);
  not1 I152_729(w_152_729, w_075_096);
  or2  I153_009(w_153_009, w_060_045, w_141_021);
  and2 I153_016(w_153_016, w_019_002, w_112_079);
  and2 I153_018(w_153_018, w_099_192, w_102_550);
  or2  I153_019(w_153_019, w_054_166, w_110_410);
  or2  I153_020(w_153_020, w_116_061, w_066_372);
  and2 I153_022(w_153_022, w_019_009, w_046_456);
  not1 I153_025(w_153_025, w_041_077);
  nand2 I153_026(w_153_026, w_060_075, w_138_246);
  or2  I153_029(w_153_029, w_145_048, w_055_234);
  nand2 I153_030(w_153_030, w_145_037, w_046_085);
  not1 I153_032(w_153_032, w_024_090);
  or2  I153_037(w_153_037, w_078_195, w_108_127);
  not1 I153_038(w_153_038, w_122_063);
  not1 I153_044(w_153_044, w_030_086);
  and2 I153_045(w_153_045, w_115_101, w_098_008);
  nand2 I153_047(w_153_047, w_005_058, w_121_125);
  or2  I153_049(w_153_049, w_017_043, w_094_370);
  not1 I153_052(w_153_052, w_105_364);
  nand2 I153_053(w_153_053, w_030_239, w_116_142);
  and2 I153_055(w_153_055, w_139_009, w_106_043);
  not1 I153_056(w_153_056, w_149_501);
  and2 I153_057(w_153_057, w_088_015, w_126_063);
  not1 I153_060(w_153_060, w_131_121);
  or2  I153_067(w_153_067, w_100_030, w_135_029);
  not1 I153_070(w_153_070, w_002_578);
  nand2 I153_072(w_153_072, w_107_304, w_111_059);
  or2  I153_073(w_153_073, w_054_412, w_017_131);
  and2 I153_085(w_153_085, w_115_036, w_014_034);
  nand2 I153_091(w_153_091, w_019_014, w_028_255);
  or2  I154_002(w_154_002, w_061_027, w_149_314);
  and2 I154_009(w_154_009, w_054_161, w_151_264);
  not1 I154_010(w_154_010, w_152_586);
  nand2 I154_025(w_154_025, w_079_029, w_148_077);
  or2  I154_030(w_154_030, w_068_136, w_007_144);
  nand2 I154_031(w_154_031, w_043_046, w_076_210);
  or2  I154_033(w_154_033, w_053_143, w_022_267);
  or2  I154_036(w_154_036, w_101_168, w_052_018);
  not1 I154_039(w_154_039, w_056_058);
  and2 I154_046(w_154_046, w_113_107, w_075_030);
  and2 I154_051(w_154_051, w_104_266, w_081_019);
  or2  I154_054(w_154_054, w_062_251, w_033_378);
  not1 I154_055(w_154_055, w_025_056);
  and2 I154_056(w_154_056, w_115_136, w_050_034);
  or2  I154_060(w_154_060, w_032_088, w_016_006);
  nand2 I154_062(w_154_062, w_091_078, w_028_018);
  not1 I154_065(w_154_065, w_117_072);
  and2 I154_075(w_154_075, w_101_049, w_125_069);
  or2  I154_078(w_154_078, w_036_018, w_082_141);
  or2  I154_080(w_154_080, w_073_374, w_100_024);
  nand2 I154_082(w_154_082, w_124_065, w_048_007);
  and2 I154_093(w_154_093, w_002_262, w_149_080);
  nand2 I154_094(w_154_094, w_094_150, w_020_372);
  nand2 I154_095(w_154_095, w_073_043, w_111_062);
  not1 I154_096(w_154_096, w_150_108);
  nand2 I154_097(w_154_097, w_002_643, w_131_212);
  and2 I154_098(w_154_098, w_126_130, w_034_064);
  not1 I154_099(w_154_099, w_136_014);
  or2  I154_103(w_154_103, w_144_190, w_143_344);
  and2 I154_110(w_154_110, w_106_081, w_049_342);
  not1 I154_112(w_154_112, w_092_264);
  and2 I154_119(w_154_119, w_037_032, w_126_135);
  not1 I154_120(w_154_120, w_146_042);
  not1 I154_121(w_154_121, w_112_054);
  or2  I154_131(w_154_131, w_071_121, w_150_008);
  or2  I155_000(w_155_000, w_002_021, w_042_369);
  or2  I155_001(w_155_001, w_000_394, w_052_046);
  or2  I155_024(w_155_024, w_072_054, w_023_142);
  or2  I155_033(w_155_033, w_072_195, w_139_014);
  and2 I155_034(w_155_034, w_110_042, w_066_406);
  not1 I155_041(w_155_041, w_046_631);
  not1 I155_045(w_155_045, w_004_167);
  and2 I155_050(w_155_050, w_074_077, w_037_330);
  nand2 I155_072(w_155_072, w_026_107, w_100_019);
  not1 I155_076(w_155_076, w_098_024);
  not1 I155_088(w_155_088, w_148_106);
  or2  I155_090(w_155_090, w_138_094, w_101_261);
  nand2 I155_102(w_155_102, w_138_248, w_061_099);
  and2 I155_103(w_155_103, w_141_107, w_057_144);
  and2 I155_109(w_155_109, w_042_192, w_049_220);
  not1 I155_122(w_155_122, w_007_023);
  not1 I155_145(w_155_145, w_122_034);
  or2  I155_148(w_155_148, w_046_263, w_008_729);
  and2 I155_149(w_155_149, w_019_014, w_097_135);
  and2 I155_180(w_155_180, w_065_606, w_131_149);
  not1 I155_192(w_155_192, w_028_106);
  and2 I155_197(w_155_197, w_051_171, w_029_055);
  or2  I155_217(w_155_217, w_119_104, w_023_106);
  not1 I155_242(w_155_242, w_041_166);
  or2  I155_252(w_155_252, w_042_281, w_099_002);
  not1 I155_276(w_155_276, w_012_073);
  nand2 I155_288(w_155_288, w_085_329, w_049_041);
  not1 I155_289(w_155_289, w_024_151);
  not1 I155_290(w_155_290, w_052_025);
  not1 I155_352(w_155_352, w_037_100);
  not1 I155_402(w_155_402, w_038_549);
  nand2 I155_403(w_155_403, w_150_300, w_073_200);
  not1 I155_405(w_155_405, w_110_425);
  nand2 I155_415(w_155_415, w_063_269, w_078_349);
  and2 I155_424(w_155_424, w_087_156, w_101_090);
  or2  I155_443(w_155_443, w_108_132, w_088_018);
  and2 I155_444(w_155_444, w_045_220, w_071_144);
  not1 I155_470(w_155_470, w_053_000);
  not1 I155_493(w_155_493, w_077_290);
  or2  I155_494(w_155_494, w_110_327, w_151_057);
  nand2 I155_508(w_155_508, w_149_367, w_001_007);
  not1 I155_531(w_155_531, w_011_570);
  or2  I156_005(w_156_005, w_052_036, w_098_035);
  and2 I156_007(w_156_007, w_015_047, w_042_415);
  or2  I156_013(w_156_013, w_003_023, w_106_044);
  not1 I156_029(w_156_029, w_089_028);
  or2  I156_032(w_156_032, w_013_573, w_011_069);
  or2  I156_041(w_156_041, w_080_120, w_043_011);
  not1 I156_044(w_156_044, w_136_020);
  or2  I156_057(w_156_057, w_039_569, w_108_188);
  nand2 I156_100(w_156_100, w_097_521, w_078_434);
  not1 I156_130(w_156_130, w_037_261);
  or2  I156_150(w_156_150, w_051_098, w_004_390);
  or2  I156_167(w_156_167, w_048_010, w_024_477);
  and2 I156_172(w_156_172, w_112_078, w_063_113);
  or2  I156_209(w_156_209, w_037_258, w_123_255);
  and2 I156_224(w_156_224, w_141_079, w_059_146);
  nand2 I156_231(w_156_231, w_055_185, w_083_017);
  and2 I156_232(w_156_232, w_012_193, w_061_103);
  nand2 I156_238(w_156_238, w_128_571, w_071_052);
  nand2 I156_242(w_156_242, w_050_237, w_057_254);
  and2 I156_261(w_156_261, w_039_324, w_038_087);
  or2  I156_289(w_156_289, w_139_020, w_078_208);
  nand2 I156_296(w_156_296, w_129_251, w_063_410);
  nand2 I156_342(w_156_342, w_028_256, w_081_003);
  nand2 I156_374(w_156_374, w_028_350, w_059_061);
  nand2 I156_386(w_156_386, w_025_000, w_011_096);
  and2 I156_428(w_156_428, w_100_053, w_058_210);
  or2  I156_430(w_156_430, w_016_001, w_105_082);
  and2 I156_467(w_156_467, w_087_408, w_110_022);
  nand2 I156_472(w_156_472, w_151_099, w_099_068);
  or2  I156_501(w_156_501, w_007_164, w_088_055);
  or2  I156_545(w_156_545, w_001_020, w_102_183);
  or2  I157_001(w_157_001, w_123_379, w_148_060);
  and2 I157_002(w_157_002, w_091_059, w_115_033);
  nand2 I157_007(w_157_007, w_154_078, w_050_384);
  not1 I157_013(w_157_013, w_114_120);
  not1 I157_021(w_157_021, w_051_014);
  or2  I157_022(w_157_022, w_026_126, w_154_094);
  or2  I157_031(w_157_031, w_058_457, w_063_387);
  not1 I157_032(w_157_032, w_052_033);
  or2  I157_036(w_157_036, w_117_058, w_035_095);
  nand2 I157_048(w_157_048, w_069_182, w_061_157);
  not1 I157_051(w_157_051, w_044_457);
  not1 I157_053(w_157_053, w_088_121);
  nand2 I157_054(w_157_054, w_016_002, w_111_039);
  not1 I157_058(w_157_058, w_089_017);
  nand2 I157_064(w_157_064, w_018_011, w_033_637);
  and2 I157_065(w_157_065, w_122_014, w_087_372);
  nand2 I157_066(w_157_066, w_149_478, w_142_587);
  and2 I157_074(w_157_074, w_026_044, w_119_012);
  not1 I157_094(w_157_094, w_080_158);
  nand2 I157_097(w_157_097, w_064_086, w_145_005);
  and2 I157_098(w_157_098, w_136_007, w_144_242);
  not1 I157_101(w_157_101, w_063_058);
  or2  I157_121(w_157_121, w_016_005, w_008_560);
  or2  I157_123(w_157_123, w_019_020, w_113_273);
  nand2 I157_124(w_157_124, w_149_063, w_104_062);
  not1 I157_126(w_157_126, w_098_028);
  and2 I157_133(w_157_133, w_105_325, w_010_151);
  nand2 I157_135(w_157_135, w_144_035, w_008_111);
  or2  I157_141(w_157_141, w_055_124, w_011_188);
  nand2 I157_148(w_157_148, w_050_009, w_130_194);
  nand2 I157_151(w_157_151, w_064_052, w_139_016);
  or2  I157_160(w_157_160, w_151_262, w_116_570);
  not1 I157_162(w_157_162, w_016_005);
  and2 I157_164(w_157_164, w_007_271, w_109_002);
  not1 I158_000(w_158_000, w_015_527);
  not1 I158_001(w_158_001, w_022_064);
  or2  I158_002(w_158_002, w_120_430, w_050_034);
  and2 I158_003(w_158_003, w_114_039, w_027_032);
  and2 I158_004(w_158_004, w_095_006, w_087_054);
  not1 I159_004(w_159_004, w_012_303);
  nand2 I159_007(w_159_007, w_098_068, w_016_004);
  or2  I159_008(w_159_008, w_138_171, w_025_101);
  nand2 I159_012(w_159_012, w_082_218, w_017_449);
  nand2 I159_013(w_159_013, w_062_100, w_056_088);
  or2  I159_018(w_159_018, w_087_037, w_046_025);
  and2 I159_024(w_159_024, w_151_013, w_124_122);
  nand2 I159_029(w_159_029, w_016_002, w_133_187);
  nand2 I159_030(w_159_030, w_121_194, w_147_040);
  not1 I159_032(w_159_032, w_155_494);
  or2  I159_037(w_159_037, w_158_000, w_142_494);
  or2  I159_039(w_159_039, w_004_015, w_148_581);
  nand2 I159_045(w_159_045, w_157_123, w_092_588);
  nand2 I159_048(w_159_048, w_029_045, w_094_432);
  not1 I159_063(w_159_063, w_129_170);
  or2  I159_065(w_159_065, w_103_045, w_013_006);
  and2 I159_074(w_159_074, w_086_022, w_038_618);
  or2  I159_077(w_159_077, w_032_226, w_036_217);
  and2 I159_078(w_159_078, w_059_364, w_119_082);
  and2 I159_079(w_159_079, w_066_315, w_129_044);
  nand2 I159_080(w_159_080, w_044_564, w_024_186);
  nand2 I159_083(w_159_083, w_077_099, w_115_061);
  not1 I159_098(w_159_098, w_027_014);
  and2 I159_101(w_159_101, w_010_455, w_074_052);
  or2  I159_108(w_159_108, w_091_088, w_099_178);
  or2  I160_039(w_160_039, w_146_124, w_073_419);
  or2  I160_049(w_160_049, w_026_328, w_014_253);
  nand2 I160_056(w_160_056, w_057_114, w_049_342);
  and2 I160_059(w_160_059, w_036_455, w_146_049);
  or2  I160_063(w_160_063, w_109_352, w_058_484);
  or2  I160_074(w_160_074, w_081_020, w_117_075);
  or2  I160_080(w_160_080, w_016_007, w_070_289);
  and2 I160_092(w_160_092, w_027_099, w_066_572);
  not1 I160_148(w_160_148, w_044_658);
  or2  I160_182(w_160_182, w_129_017, w_150_449);
  not1 I160_223(w_160_223, w_134_147);
  and2 I160_237(w_160_237, w_037_149, w_017_606);
  not1 I160_245(w_160_245, w_116_601);
  nand2 I160_299(w_160_299, w_046_229, w_108_119);
  and2 I160_382(w_160_382, w_099_174, w_006_165);
  and2 I160_394(w_160_394, w_031_260, w_092_560);
  not1 I160_398(w_160_398, w_118_036);
  nand2 I160_405(w_160_405, w_121_128, w_097_049);
  and2 I160_426(w_160_426, w_105_144, w_067_027);
  not1 I160_433(w_160_433, w_075_139);
  nand2 I160_449(w_160_449, w_051_226, w_135_528);
  and2 I160_465(w_160_465, w_076_319, w_145_005);
  and2 I160_479(w_160_479, w_065_015, w_099_133);
  and2 I160_580(w_160_580, w_095_039, w_119_053);
  and2 I160_601(w_160_601, w_040_386, w_045_006);
  nand2 I160_611(w_160_611, w_027_135, w_035_098);
  not1 I160_634(w_160_634, w_012_019);
  or2  I160_667(w_160_667, w_056_427, w_017_620);
  or2  I160_673(w_160_673, w_070_444, w_042_310);
  nand2 I160_699(w_160_699, w_007_068, w_151_048);
  not1 I160_706(w_160_706, w_157_148);
  and2 I160_753(w_160_753, w_011_336, w_039_167);
  or2  I160_793(w_160_793, w_134_114, w_076_111);
  not1 I161_009(w_161_009, w_138_023);
  or2  I161_013(w_161_013, w_081_002, w_153_045);
  not1 I161_023(w_161_023, w_047_311);
  and2 I161_026(w_161_026, w_060_033, w_060_259);
  not1 I161_035(w_161_035, w_038_370);
  nand2 I161_065(w_161_065, w_114_186, w_026_299);
  nand2 I161_071(w_161_071, w_095_001, w_094_021);
  or2  I161_074(w_161_074, w_035_126, w_160_237);
  or2  I161_079(w_161_079, w_094_475, w_132_289);
  not1 I161_093(w_161_093, w_131_144);
  not1 I161_121(w_161_121, w_066_243);
  not1 I161_133(w_161_133, w_010_224);
  and2 I161_134(w_161_134, w_153_072, w_032_398);
  or2  I161_135(w_161_135, w_075_155, w_093_497);
  not1 I161_153(w_161_153, w_156_428);
  not1 I161_155(w_161_155, w_058_681);
  not1 I161_160(w_161_160, w_067_280);
  and2 I161_183(w_161_183, w_037_286, w_021_068);
  nand2 I161_272(w_161_272, w_114_037, w_015_650);
  or2  I161_294(w_161_294, w_056_365, w_054_138);
  nand2 I161_326(w_161_326, w_143_401, w_160_063);
  and2 I161_365(w_161_365, w_032_321, w_114_116);
  and2 I161_369(w_161_369, w_101_285, w_014_014);
  not1 I161_394(w_161_394, w_148_060);
  and2 I161_446(w_161_446, w_051_195, w_058_179);
  nand2 I161_451(w_161_451, w_034_033, w_104_188);
  nand2 I161_460(w_161_460, w_028_143, w_113_034);
  or2  I161_461(w_161_461, w_063_064, w_053_126);
  or2  I161_472(w_161_472, w_048_016, w_056_145);
  not1 I161_487(w_161_487, w_043_034);
  not1 I161_514(w_161_514, w_131_000);
  and2 I161_533(w_161_533, w_100_082, w_104_053);
  or2  I161_565(w_161_565, w_074_303, w_128_580);
  or2  I161_567(w_161_567, w_149_032, w_122_009);
  or2  I161_607(w_161_607, w_051_218, w_038_132);
  and2 I162_000(w_162_000, w_092_609, w_135_184);
  not1 I162_001(w_162_001, w_036_444);
  or2  I162_002(w_162_002, w_017_038, w_033_770);
  not1 I162_003(w_162_003, w_044_335);
  not1 I162_004(w_162_004, w_077_140);
  not1 I162_006(w_162_006, w_105_220);
  not1 I162_008(w_162_008, w_149_079);
  and2 I162_013(w_162_013, w_047_040, w_004_455);
  nand2 I162_015(w_162_015, w_018_026, w_048_004);
  not1 I162_017(w_162_017, w_028_263);
  or2  I162_019(w_162_019, w_123_503, w_089_132);
  not1 I162_020(w_162_020, w_093_395);
  nand2 I162_021(w_162_021, w_092_043, w_081_011);
  not1 I162_022(w_162_022, w_116_424);
  not1 I162_023(w_162_023, w_076_072);
  not1 I162_024(w_162_024, w_159_079);
  nand2 I162_025(w_162_025, w_076_295, w_071_276);
  and2 I163_036(w_163_036, w_121_127, w_009_362);
  or2  I163_050(w_163_050, w_082_270, w_078_183);
  not1 I163_065(w_163_065, w_102_546);
  nand2 I163_077(w_163_077, w_054_178, w_022_248);
  nand2 I163_078(w_163_078, w_094_234, w_029_011);
  nand2 I163_081(w_163_081, w_097_082, w_084_008);
  and2 I163_091(w_163_091, w_047_050, w_044_643);
  nand2 I163_099(w_163_099, w_086_275, w_073_003);
  nand2 I163_132(w_163_132, w_065_256, w_063_208);
  and2 I163_133(w_163_133, w_154_010, w_007_031);
  nand2 I163_157(w_163_157, w_145_022, w_102_014);
  not1 I163_159(w_163_159, w_018_016);
  or2  I163_162(w_163_162, w_057_291, w_049_049);
  or2  I163_163(w_163_163, w_046_047, w_061_100);
  not1 I163_178(w_163_178, w_134_261);
  not1 I163_185(w_163_185, w_012_113);
  and2 I163_188(w_163_188, w_091_074, w_104_112);
  nand2 I163_189(w_163_189, w_079_040, w_016_003);
  or2  I163_221(w_163_221, w_058_581, w_153_055);
  or2  I163_225(w_163_225, w_096_005, w_103_260);
  and2 I163_228(w_163_228, w_010_560, w_029_117);
  or2  I163_243(w_163_243, w_132_217, w_088_021);
  nand2 I163_249(w_163_249, w_145_079, w_015_027);
  or2  I163_266(w_163_266, w_033_331, w_000_066);
  not1 I163_284(w_163_284, w_154_119);
  nand2 I163_307(w_163_307, w_154_098, w_153_016);
  nand2 I163_327(w_163_327, w_116_124, w_155_276);
  not1 I163_343(w_163_343, w_016_007);
  not1 I163_416(w_163_416, w_044_653);
  or2  I163_428(w_163_428, w_005_013, w_000_054);
  not1 I163_445(w_163_445, w_128_094);
  nand2 I163_478(w_163_478, w_000_711, w_129_337);
  not1 I163_486(w_163_486, w_153_032);
  or2  I163_488(w_163_488, w_038_405, w_065_165);
  or2  I163_489(w_163_489, w_140_088, w_096_004);
  nand2 I163_491(w_163_491, w_040_493, w_131_059);
  or2  I163_497(w_163_497, w_079_056, w_141_114);
  or2  I163_509(w_163_509, w_076_364, w_003_030);
  not1 I163_515(w_163_515, w_148_595);
  not1 I163_519(w_163_519, w_131_187);
  or2  I163_567(w_163_567, w_076_294, w_099_248);
  nand2 I163_574(w_163_574, w_065_609, w_131_109);
  nand2 I163_593(w_163_593, w_155_102, w_117_011);
  not1 I164_004(w_164_004, w_099_141);
  nand2 I164_005(w_164_005, w_012_188, w_068_167);
  not1 I164_023(w_164_023, w_115_131);
  nand2 I164_079(w_164_079, w_023_195, w_143_107);
  nand2 I164_085(w_164_085, w_016_005, w_142_559);
  nand2 I164_093(w_164_093, w_147_031, w_134_173);
  and2 I164_119(w_164_119, w_006_093, w_132_099);
  nand2 I164_127(w_164_127, w_132_255, w_042_339);
  or2  I164_141(w_164_141, w_129_333, w_152_337);
  or2  I164_204(w_164_204, w_079_054, w_125_318);
  or2  I164_235(w_164_235, w_043_016, w_036_037);
  nand2 I164_241(w_164_241, w_096_003, w_063_421);
  not1 I164_244(w_164_244, w_115_126);
  not1 I164_266(w_164_266, w_152_714);
  not1 I164_277(w_164_277, w_146_008);
  or2  I164_291(w_164_291, w_012_065, w_019_017);
  not1 I164_294(w_164_294, w_120_489);
  nand2 I164_302(w_164_302, w_114_119, w_081_001);
  or2  I164_339(w_164_339, w_068_275, w_108_103);
  not1 I164_348(w_164_348, w_145_077);
  and2 I164_374(w_164_374, w_034_059, w_133_117);
  or2  I164_387(w_164_387, w_133_223, w_131_254);
  not1 I164_390(w_164_390, w_016_008);
  and2 I164_395(w_164_395, w_031_377, w_029_058);
  not1 I164_424(w_164_424, w_004_361);
  and2 I164_453(w_164_453, w_151_247, w_051_222);
  not1 I164_502(w_164_502, w_026_580);
  not1 I164_588(w_164_588, w_162_022);
  and2 I164_593(w_164_593, w_010_339, w_005_120);
  nand2 I165_003(w_165_003, w_102_195, w_130_071);
  or2  I165_007(w_165_007, w_157_048, w_009_048);
  not1 I165_009(w_165_009, w_002_398);
  and2 I165_012(w_165_012, w_056_557, w_001_035);
  and2 I165_015(w_165_015, w_076_209, w_082_051);
  nand2 I165_017(w_165_017, w_032_106, w_038_567);
  and2 I165_025(w_165_025, w_146_107, w_095_042);
  nand2 I165_026(w_165_026, w_120_633, w_007_047);
  not1 I165_028(w_165_028, w_062_406);
  not1 I165_032(w_165_032, w_072_186);
  not1 I165_034(w_165_034, w_034_016);
  and2 I165_043(w_165_043, w_027_078, w_096_000);
  and2 I165_049(w_165_049, w_130_171, w_110_364);
  and2 I165_050(w_165_050, w_138_326, w_121_162);
  not1 I165_051(w_165_051, w_138_206);
  or2  I165_054(w_165_054, w_075_016, w_069_034);
  or2  I165_056(w_165_056, w_062_282, w_006_182);
  or2  I165_059(w_165_059, w_015_431, w_002_669);
  and2 I165_071(w_165_071, w_117_014, w_132_026);
  nand2 I165_079(w_165_079, w_029_074, w_060_354);
  not1 I165_088(w_165_088, w_132_281);
  or2  I165_094(w_165_094, w_071_063, w_096_004);
  nand2 I165_095(w_165_095, w_063_177, w_000_100);
  not1 I165_096(w_165_096, w_126_100);
  nand2 I165_101(w_165_101, w_044_712, w_091_157);
  not1 I165_105(w_165_105, w_095_047);
  nand2 I165_109(w_165_109, w_107_080, w_046_319);
  or2  I165_110(w_165_110, w_030_338, w_097_121);
  and2 I165_111(w_165_111, w_012_071, w_152_234);
  nand2 I165_146(w_165_146, w_027_164, w_124_056);
  or2  I165_150(w_165_150, w_060_169, w_120_223);
  not1 I165_155(w_165_155, w_106_093);
  nand2 I166_010(w_166_010, w_100_044, w_088_063);
  and2 I166_040(w_166_040, w_002_229, w_045_000);
  nand2 I166_041(w_166_041, w_112_134, w_085_001);
  or2  I166_056(w_166_056, w_016_000, w_067_037);
  nand2 I166_076(w_166_076, w_094_600, w_119_164);
  and2 I166_081(w_166_081, w_140_161, w_070_424);
  nand2 I166_095(w_166_095, w_105_216, w_073_632);
  nand2 I166_097(w_166_097, w_091_032, w_058_029);
  nand2 I166_103(w_166_103, w_147_226, w_159_004);
  and2 I166_109(w_166_109, w_117_029, w_038_551);
  or2  I166_110(w_166_110, w_085_027, w_062_083);
  nand2 I166_115(w_166_115, w_054_122, w_102_093);
  and2 I166_123(w_166_123, w_151_453, w_108_200);
  or2  I166_127(w_166_127, w_030_099, w_110_017);
  nand2 I166_138(w_166_138, w_004_218, w_087_381);
  nand2 I166_145(w_166_145, w_048_001, w_099_051);
  not1 I166_152(w_166_152, w_112_022);
  or2  I166_165(w_166_165, w_107_379, w_056_224);
  nand2 I166_199(w_166_199, w_147_003, w_078_058);
  not1 I166_202(w_166_202, w_033_200);
  not1 I166_219(w_166_219, w_080_054);
  not1 I166_248(w_166_248, w_113_198);
  not1 I166_268(w_166_268, w_032_122);
  not1 I166_279(w_166_279, w_044_033);
  or2  I166_282(w_166_282, w_035_104, w_020_315);
  nand2 I166_287(w_166_287, w_014_108, w_110_275);
  nand2 I166_288(w_166_288, w_128_268, w_100_065);
  or2  I166_299(w_166_299, w_036_241, w_138_069);
  not1 I166_305(w_166_305, w_111_034);
  and2 I166_313(w_166_313, w_151_148, w_052_002);
  not1 I166_322(w_166_322, w_055_066);
  or2  I167_005(w_167_005, w_029_038, w_040_000);
  not1 I167_014(w_167_014, w_023_063);
  not1 I167_016(w_167_016, w_058_061);
  not1 I167_022(w_167_022, w_061_219);
  not1 I167_031(w_167_031, w_086_124);
  not1 I167_040(w_167_040, w_126_024);
  and2 I167_041(w_167_041, w_137_042, w_139_021);
  and2 I167_043(w_167_043, w_155_443, w_089_100);
  nand2 I167_049(w_167_049, w_028_135, w_104_068);
  not1 I167_050(w_167_050, w_047_072);
  nand2 I167_057(w_167_057, w_161_160, w_102_316);
  not1 I167_068(w_167_068, w_063_005);
  not1 I167_078(w_167_078, w_091_042);
  or2  I167_080(w_167_080, w_081_009, w_091_122);
  or2  I167_081(w_167_081, w_086_049, w_119_018);
  not1 I167_082(w_167_082, w_046_028);
  or2  I167_099(w_167_099, w_106_108, w_045_091);
  or2  I167_100(w_167_100, w_110_124, w_058_538);
  and2 I167_107(w_167_107, w_003_071, w_111_099);
  or2  I167_108(w_167_108, w_016_005, w_064_345);
  and2 I167_122(w_167_122, w_132_231, w_049_231);
  or2  I167_131(w_167_131, w_112_085, w_036_039);
  and2 I167_140(w_167_140, w_054_137, w_014_173);
  or2  I167_145(w_167_145, w_008_495, w_100_093);
  not1 I167_152(w_167_152, w_129_078);
  and2 I167_161(w_167_163, w_167_162, w_093_028);
  or2  I167_162(w_167_164, w_092_203, w_167_163);
  not1 I167_163(w_167_165, w_167_164);
  and2 I167_164(w_167_166, w_167_183, w_167_165);
  and2 I167_165(w_167_162, w_112_039, w_167_166);
  nand2 I167_166(w_167_171, w_167_170, w_092_080);
  and2 I167_167(w_167_172, w_167_171, w_073_299);
  or2  I167_168(w_167_173, w_060_171, w_167_172);
  and2 I167_169(w_167_174, w_012_200, w_167_173);
  not1 I167_170(w_167_175, w_167_174);
  and2 I167_171(w_167_176, w_069_033, w_167_175);
  not1 I167_172(w_167_177, w_167_176);
  not1 I167_173(w_167_178, w_167_177);
  nand2 I167_174(w_167_179, w_167_178, w_148_004);
  or2  I167_175(w_167_180, w_167_179, w_028_588);
  and2 I167_176(w_167_181, w_012_289, w_167_180);
  not1 I167_177(w_167_170, w_167_166);
  and2 I167_178(w_167_183, w_097_144, w_167_181);
  and2 I168_014(w_168_014, w_012_040, w_060_118);
  or2  I168_028(w_168_028, w_078_061, w_125_497);
  nand2 I168_088(w_168_088, w_048_019, w_065_275);
  not1 I168_110(w_168_110, w_038_146);
  and2 I168_126(w_168_126, w_129_117, w_014_035);
  nand2 I168_143(w_168_143, w_038_486, w_075_019);
  and2 I168_147(w_168_147, w_067_343, w_015_618);
  not1 I168_151(w_168_151, w_124_070);
  or2  I168_152(w_168_152, w_095_002, w_129_349);
  or2  I168_159(w_168_159, w_155_041, w_122_010);
  and2 I168_171(w_168_171, w_155_531, w_004_245);
  not1 I168_216(w_168_216, w_167_099);
  not1 I168_232(w_168_232, w_010_050);
  not1 I168_266(w_168_266, w_138_078);
  not1 I168_315(w_168_315, w_125_399);
  not1 I168_354(w_168_354, w_149_484);
  and2 I168_359(w_168_359, w_125_129, w_073_624);
  nand2 I168_380(w_168_380, w_165_071, w_057_082);
  and2 I168_381(w_168_381, w_149_056, w_126_034);
  nand2 I168_419(w_168_419, w_146_303, w_044_027);
  nand2 I168_448(w_168_448, w_130_254, w_159_024);
  nand2 I168_452(w_168_452, w_006_042, w_012_147);
  and2 I168_492(w_168_492, w_005_063, w_014_192);
  or2  I168_506(w_168_506, w_100_125, w_082_066);
  and2 I168_542(w_168_542, w_074_196, w_109_053);
  not1 I169_004(w_169_004, w_026_344);
  not1 I169_008(w_169_008, w_095_006);
  nand2 I169_062(w_169_062, w_090_478, w_157_053);
  nand2 I169_101(w_169_101, w_033_355, w_039_710);
  not1 I169_103(w_169_103, w_120_083);
  or2  I169_106(w_169_106, w_060_050, w_068_008);
  not1 I169_141(w_169_141, w_047_137);
  nand2 I169_170(w_169_170, w_026_662, w_087_137);
  nand2 I169_187(w_169_187, w_014_175, w_167_005);
  and2 I169_192(w_169_192, w_141_053, w_077_310);
  or2  I169_200(w_169_200, w_033_313, w_044_452);
  and2 I169_218(w_169_218, w_150_294, w_073_537);
  or2  I169_221(w_169_221, w_034_040, w_079_051);
  nand2 I169_236(w_169_236, w_005_139, w_007_316);
  not1 I169_273(w_169_273, w_038_331);
  or2  I169_279(w_169_279, w_046_484, w_086_307);
  not1 I169_283(w_169_283, w_044_650);
  not1 I169_296(w_169_296, w_045_196);
  and2 I169_303(w_169_303, w_119_109, w_136_004);
  not1 I169_305(w_169_305, w_072_048);
  nand2 I169_318(w_169_318, w_109_009, w_025_261);
  and2 I169_323(w_169_323, w_161_026, w_113_323);
  or2  I169_333(w_169_333, w_129_065, w_114_032);
  and2 I169_344(w_169_344, w_020_170, w_155_424);
  and2 I169_365(w_169_365, w_021_214, w_083_153);
  and2 I169_380(w_169_380, w_106_160, w_045_358);
  nand2 I169_405(w_169_405, w_110_197, w_095_057);
  and2 I169_437(w_169_437, w_133_244, w_153_056);
  and2 I170_015(w_170_015, w_142_258, w_068_098);
  nand2 I170_017(w_170_017, w_098_034, w_114_150);
  not1 I170_040(w_170_040, w_102_479);
  and2 I170_053(w_170_053, w_096_002, w_092_089);
  not1 I170_085(w_170_085, w_029_044);
  not1 I170_139(w_170_139, w_143_061);
  not1 I170_172(w_170_172, w_072_190);
  not1 I170_185(w_170_185, w_104_080);
  or2  I170_194(w_170_194, w_063_101, w_115_040);
  not1 I170_198(w_170_198, w_020_280);
  nand2 I170_209(w_170_209, w_017_019, w_012_057);
  or2  I170_212(w_170_212, w_061_143, w_045_308);
  and2 I170_222(w_170_222, w_006_072, w_101_244);
  not1 I170_226(w_170_226, w_164_005);
  or2  I170_240(w_170_240, w_037_235, w_135_609);
  and2 I170_248(w_170_248, w_053_155, w_042_406);
  not1 I170_250(w_170_250, w_073_439);
  or2  I170_277(w_170_277, w_056_252, w_057_126);
  and2 I170_282(w_170_282, w_161_487, w_129_342);
  or2  I170_310(w_170_310, w_088_005, w_023_128);
  or2  I170_331(w_170_331, w_102_229, w_002_499);
  or2  I170_399(w_170_399, w_120_594, w_009_444);
  and2 I170_423(w_170_423, w_165_146, w_019_014);
  and2 I171_013(w_171_013, w_097_085, w_052_012);
  or2  I171_119(w_171_119, w_085_116, w_129_082);
  nand2 I171_124(w_171_124, w_066_556, w_062_607);
  nand2 I171_135(w_171_135, w_114_007, w_091_125);
  not1 I171_162(w_171_162, w_140_233);
  nand2 I171_176(w_171_176, w_097_139, w_151_203);
  or2  I171_192(w_171_192, w_029_103, w_089_185);
  or2  I171_195(w_171_195, w_086_158, w_141_168);
  not1 I171_221(w_171_221, w_075_135);
  not1 I171_228(w_171_228, w_057_008);
  or2  I171_252(w_171_252, w_044_335, w_107_318);
  not1 I171_263(w_171_263, w_119_099);
  not1 I171_265(w_171_265, w_012_233);
  or2  I171_303(w_171_303, w_063_139, w_165_059);
  and2 I171_322(w_171_322, w_043_011, w_105_202);
  not1 I171_333(w_171_333, w_011_563);
  nand2 I171_334(w_171_334, w_119_188, w_166_040);
  and2 I171_363(w_171_363, w_018_028, w_072_260);
  nand2 I171_384(w_171_384, w_135_200, w_094_027);
  not1 I171_408(w_171_408, w_112_107);
  and2 I171_412(w_171_412, w_014_138, w_004_288);
  or2  I171_425(w_171_425, w_041_494, w_039_552);
  not1 I171_450(w_171_450, w_086_187);
  not1 I171_470(w_171_470, w_099_075);
  or2  I171_479(w_171_479, w_121_053, w_104_040);
  and2 I171_495(w_171_495, w_012_332, w_117_063);
  and2 I171_560(w_171_560, w_162_024, w_104_216);
  and2 I171_578(w_171_578, w_090_126, w_111_061);
  nand2 I171_606(w_171_606, w_128_122, w_100_085);
  nand2 I171_611(w_171_611, w_016_004, w_047_077);
  and2 I171_654(w_171_654, w_057_023, w_050_207);
  or2  I171_706(w_171_706, w_061_338, w_038_268);
  not1 I171_711(w_171_711, w_020_364);
  not1 I171_722(w_171_722, w_124_156);
  or2  I171_731(w_171_731, w_161_607, w_035_103);
  not1 I172_000(w_172_000, w_063_076);
  and2 I172_001(w_172_001, w_015_441, w_100_125);
  nand2 I172_002(w_172_002, w_143_106, w_135_587);
  nand2 I172_003(w_172_003, w_115_251, w_022_136);
  not1 I172_005(w_172_005, w_117_028);
  not1 I172_006(w_172_006, w_050_035);
  nand2 I172_007(w_172_007, w_080_120, w_042_157);
  nand2 I172_012(w_172_012, w_063_509, w_156_467);
  nand2 I172_013(w_172_013, w_035_054, w_107_313);
  not1 I172_024(w_172_024, w_143_211);
  not1 I172_030(w_172_030, w_149_450);
  and2 I172_031(w_172_031, w_113_300, w_014_243);
  nand2 I172_033(w_172_033, w_108_024, w_013_065);
  and2 I172_035(w_172_035, w_129_351, w_068_275);
  not1 I172_039(w_172_039, w_121_084);
  not1 I172_040(w_172_040, w_126_018);
  nand2 I172_041(w_172_041, w_116_092, w_103_053);
  and2 I172_042(w_172_042, w_052_014, w_113_062);
  or2  I172_044(w_172_044, w_093_151, w_079_015);
  and2 I172_046(w_172_046, w_119_027, w_054_041);
  nand2 I172_048(w_172_048, w_142_792, w_071_148);
  and2 I172_049(w_172_049, w_004_007, w_132_422);
  or2  I172_052(w_172_052, w_113_172, w_102_022);
  not1 I172_053(w_172_053, w_156_501);
  nand2 I173_001(w_173_001, w_085_146, w_057_145);
  not1 I173_002(w_173_002, w_132_291);
  and2 I173_003(w_173_003, w_139_007, w_048_000);
  or2  I173_004(w_173_004, w_090_072, w_018_011);
  not1 I173_005(w_173_005, w_000_610);
  not1 I173_008(w_173_008, w_076_036);
  or2  I173_009(w_173_009, w_165_043, w_035_055);
  nand2 I173_011(w_173_011, w_047_132, w_098_069);
  not1 I173_012(w_173_012, w_168_419);
  or2  I173_013(w_173_013, w_075_120, w_145_075);
  nand2 I173_015(w_173_015, w_142_348, w_140_188);
  not1 I173_016(w_173_016, w_128_196);
  not1 I173_017(w_173_017, w_102_563);
  or2  I173_018(w_173_018, w_119_165, w_169_333);
  not1 I173_022(w_173_022, w_155_122);
  not1 I173_023(w_173_023, w_117_020);
  and2 I173_025(w_173_025, w_155_088, w_099_141);
  nand2 I173_026(w_173_026, w_036_322, w_131_140);
  nand2 I173_027(w_173_027, w_092_062, w_146_255);
  and2 I173_028(w_173_028, w_116_231, w_036_281);
  and2 I173_030(w_173_030, w_169_103, w_093_417);
  or2  I173_031(w_173_031, w_022_026, w_157_001);
  nand2 I174_001(w_174_001, w_043_003, w_085_246);
  or2  I174_004(w_174_004, w_159_012, w_056_499);
  or2  I174_010(w_174_010, w_129_156, w_000_041);
  nand2 I174_014(w_174_014, w_119_029, w_112_197);
  not1 I174_024(w_174_024, w_032_545);
  and2 I174_028(w_174_028, w_091_077, w_009_094);
  or2  I174_029(w_174_029, w_058_156, w_041_561);
  or2  I174_044(w_174_044, w_092_073, w_142_499);
  nand2 I174_060(w_174_060, w_135_119, w_007_006);
  not1 I174_066(w_174_066, w_074_117);
  and2 I174_072(w_174_072, w_124_242, w_096_001);
  and2 I174_075(w_174_075, w_012_319, w_090_063);
  nand2 I174_083(w_174_083, w_143_000, w_003_064);
  and2 I174_088(w_174_088, w_023_047, w_001_032);
  not1 I174_090(w_174_090, w_115_169);
  not1 I174_092(w_174_092, w_095_022);
  and2 I174_093(w_174_093, w_073_507, w_012_034);
  not1 I174_096(w_174_096, w_089_167);
  not1 I174_098(w_174_098, w_067_163);
  and2 I174_104(w_174_104, w_112_010, w_112_025);
  or2  I174_107(w_174_107, w_037_200, w_017_359);
  not1 I174_110(w_174_110, w_107_157);
  or2  I175_018(w_175_018, w_074_321, w_089_136);
  and2 I175_019(w_175_019, w_165_015, w_162_008);
  nand2 I175_022(w_175_022, w_126_117, w_071_048);
  and2 I175_025(w_175_025, w_118_041, w_036_258);
  nand2 I175_026(w_175_026, w_001_004, w_082_486);
  and2 I175_038(w_175_038, w_072_052, w_137_255);
  or2  I175_056(w_175_056, w_145_020, w_138_083);
  and2 I175_083(w_175_083, w_169_405, w_110_250);
  and2 I175_103(w_175_103, w_077_560, w_138_308);
  or2  I175_108(w_175_108, w_091_122, w_119_175);
  nand2 I175_141(w_175_141, w_075_097, w_098_074);
  nand2 I175_144(w_175_144, w_039_368, w_090_151);
  nand2 I175_156(w_175_156, w_046_496, w_039_260);
  or2  I175_167(w_175_167, w_123_505, w_015_275);
  nand2 I175_208(w_175_208, w_028_033, w_171_606);
  or2  I175_221(w_175_221, w_014_043, w_042_061);
  nand2 I175_240(w_175_240, w_163_091, w_151_116);
  not1 I175_285(w_175_285, w_122_063);
  not1 I175_373(w_175_373, w_041_279);
  not1 I175_417(w_175_417, w_134_251);
  and2 I175_422(w_175_422, w_102_047, w_109_385);
  nand2 I175_464(w_175_464, w_113_008, w_002_144);
  or2  I175_477(w_175_477, w_125_003, w_009_483);
  nand2 I175_488(w_175_488, w_140_073, w_109_279);
  and2 I175_504(w_175_504, w_084_029, w_073_688);
  or2  I175_549(w_175_549, w_144_062, w_001_003);
  not1 I175_558(w_175_558, w_009_273);
  and2 I175_594(w_175_594, w_164_390, w_166_095);
  nand2 I175_615(w_175_615, w_077_058, w_003_005);
  or2  I176_001(w_176_001, w_169_141, w_085_040);
  not1 I176_002(w_176_002, w_039_553);
  not1 I176_008(w_176_008, w_035_060);
  nand2 I176_049(w_176_049, w_033_614, w_004_238);
  or2  I176_059(w_176_059, w_161_451, w_141_128);
  not1 I176_080(w_176_080, w_013_169);
  not1 I176_085(w_176_085, w_064_215);
  or2  I176_097(w_176_097, w_090_464, w_105_249);
  and2 I176_110(w_176_110, w_174_004, w_119_063);
  or2  I176_129(w_176_129, w_009_380, w_038_538);
  not1 I176_136(w_176_136, w_173_011);
  and2 I176_138(w_176_138, w_171_195, w_078_566);
  nand2 I176_148(w_176_148, w_152_729, w_089_094);
  and2 I176_151(w_176_151, w_002_592, w_103_232);
  and2 I176_158(w_176_158, w_002_158, w_138_066);
  nand2 I176_170(w_176_170, w_078_084, w_151_175);
  and2 I177_006(w_177_006, w_001_032, w_084_032);
  not1 I177_008(w_177_008, w_047_065);
  and2 I177_014(w_177_014, w_101_243, w_171_706);
  and2 I177_024(w_177_024, w_044_154, w_092_200);
  and2 I177_025(w_177_025, w_077_245, w_119_123);
  or2  I177_036(w_177_036, w_014_088, w_032_322);
  not1 I177_085(w_177_085, w_011_474);
  or2  I177_102(w_177_102, w_167_145, w_167_049);
  not1 I177_108(w_177_108, w_032_102);
  and2 I177_160(w_177_160, w_073_484, w_165_034);
  and2 I177_166(w_177_166, w_113_158, w_081_001);
  or2  I177_178(w_177_178, w_133_344, w_157_066);
  nand2 I177_238(w_177_238, w_099_278, w_009_380);
  or2  I177_258(w_177_258, w_155_217, w_174_072);
  and2 I177_266(w_177_266, w_029_029, w_138_231);
  and2 I177_280(w_177_280, w_031_472, w_114_047);
  not1 I177_288(w_177_288, w_088_102);
  nand2 I177_307(w_177_307, w_156_242, w_003_053);
  nand2 I177_310(w_177_310, w_126_112, w_151_086);
  nand2 I177_333(w_177_333, w_073_053, w_094_527);
  and2 I177_375(w_177_375, w_051_366, w_136_007);
  and2 I177_385(w_177_385, w_110_376, w_168_354);
  not1 I177_399(w_177_399, w_047_420);
  nand2 I177_402(w_177_402, w_012_183, w_088_080);
  nand2 I177_405(w_177_405, w_116_532, w_123_122);
  nand2 I178_005(w_178_005, w_112_187, w_063_114);
  not1 I178_006(w_178_006, w_010_186);
  and2 I178_009(w_178_009, w_159_077, w_024_452);
  not1 I178_015(w_178_015, w_125_332);
  or2  I178_028(w_178_028, w_022_024, w_038_532);
  not1 I178_036(w_178_036, w_148_398);
  or2  I178_043(w_178_043, w_119_050, w_011_344);
  nand2 I178_049(w_178_049, w_142_365, w_063_181);
  or2  I178_054(w_178_054, w_175_464, w_117_078);
  and2 I178_067(w_178_067, w_043_018, w_105_123);
  nand2 I178_075(w_178_075, w_029_039, w_032_331);
  nand2 I178_076(w_178_076, w_065_542, w_052_011);
  and2 I178_077(w_178_077, w_117_062, w_024_096);
  not1 I178_095(w_178_095, w_055_192);
  nand2 I178_097(w_178_097, w_056_231, w_117_050);
  and2 I178_099(w_178_099, w_093_442, w_109_279);
  not1 I178_102(w_178_102, w_006_229);
  and2 I178_107(w_178_107, w_165_101, w_153_070);
  and2 I178_113(w_178_115, w_178_114, w_178_131);
  and2 I178_114(w_178_116, w_014_238, w_178_115);
  not1 I178_115(w_178_114, w_178_116);
  or2  I178_116(w_178_121, w_178_120, w_132_059);
  and2 I178_117(w_178_122, w_178_121, w_077_044);
  nand2 I178_118(w_178_123, w_029_004, w_178_122);
  nand2 I178_119(w_178_124, w_178_123, w_146_291);
  and2 I178_120(w_178_125, w_178_124, w_136_031);
  not1 I178_121(w_178_126, w_178_125);
  or2  I178_122(w_178_127, w_178_126, w_017_055);
  not1 I178_123(w_178_128, w_178_127);
  and2 I178_124(w_178_129, w_178_128, w_005_137);
  not1 I178_125(w_178_120, w_178_115);
  and2 I178_126(w_178_131, w_091_095, w_178_129);
  not1 I179_023(w_179_023, w_163_488);
  not1 I179_039(w_179_039, w_011_083);
  or2  I179_044(w_179_044, w_037_332, w_053_096);
  not1 I179_079(w_179_079, w_023_117);
  or2  I179_140(w_179_140, w_054_116, w_079_003);
  not1 I179_141(w_179_141, w_154_056);
  nand2 I179_159(w_179_159, w_167_107, w_067_347);
  nand2 I179_164(w_179_164, w_168_171, w_087_065);
  not1 I179_184(w_179_184, w_126_064);
  or2  I179_188(w_179_188, w_069_120, w_042_130);
  not1 I179_203(w_179_203, w_043_047);
  or2  I179_204(w_179_204, w_133_085, w_076_158);
  not1 I179_416(w_179_416, w_117_051);
  nand2 I179_423(w_179_423, w_058_306, w_093_086);
  nand2 I179_507(w_179_507, w_146_198, w_037_104);
  not1 I179_579(w_179_579, w_068_267);
  or2  I179_583(w_179_583, w_033_613, w_043_001);
  or2  I179_620(w_179_620, w_103_121, w_110_239);
  not1 I179_710(w_179_710, w_006_092);
  not1 I179_721(w_179_721, w_153_072);
  and2 I179_737(w_179_737, w_109_011, w_057_194);
  nand2 I179_745(w_179_745, w_076_173, w_125_031);
  and2 I179_767(w_179_767, w_102_436, w_001_027);
  nand2 I179_768(w_179_768, w_133_201, w_101_238);
  and2 I179_769(w_178_118, w_104_216, w_178_114);
  nand2 I180_001(w_180_001, w_166_299, w_090_405);
  or2  I180_002(w_180_002, w_120_695, w_043_039);
  and2 I180_003(w_180_003, w_054_166, w_025_106);
  or2  I180_007(w_180_007, w_139_011, w_105_091);
  not1 I180_008(w_180_008, w_092_391);
  and2 I180_009(w_180_009, w_109_264, w_153_091);
  nand2 I180_010(w_180_010, w_178_118, w_001_023);
  not1 I180_011(w_180_011, w_039_539);
  or2  I180_012(w_180_012, w_106_181, w_097_331);
  or2  I180_013(w_180_013, w_139_004, w_135_110);
  or2  I180_014(w_180_014, w_095_029, w_083_046);
  and2 I180_015(w_180_015, w_047_318, w_061_311);
  or2  I180_016(w_180_016, w_086_332, w_100_125);
  not1 I180_019(w_180_019, w_158_001);
  nand2 I180_020(w_180_020, w_113_211, w_060_097);
  not1 I180_021(w_180_021, w_015_099);
  nand2 I180_023(w_180_023, w_090_168, w_117_055);
  not1 I180_024(w_180_024, w_179_188);
  and2 I180_025(w_180_025, w_115_125, w_025_110);
  or2  I180_026(w_180_026, w_068_308, w_043_022);
  or2  I181_002(w_181_002, w_049_140, w_035_101);
  nand2 I181_039(w_181_039, w_030_077, w_046_300);
  or2  I181_048(w_181_048, w_108_145, w_067_363);
  or2  I181_058(w_181_058, w_017_611, w_126_047);
  nand2 I181_064(w_181_064, w_106_072, w_004_491);
  not1 I181_118(w_181_118, w_006_030);
  or2  I181_123(w_181_123, w_086_098, w_135_240);
  not1 I181_132(w_181_132, w_123_187);
  not1 I181_142(w_181_142, w_141_168);
  not1 I181_147(w_181_147, w_132_056);
  and2 I181_153(w_181_153, w_102_442, w_044_535);
  not1 I181_169(w_181_169, w_067_253);
  or2  I181_195(w_181_195, w_084_029, w_027_191);
  not1 I181_205(w_181_205, w_025_218);
  not1 I181_208(w_181_208, w_055_285);
  and2 I181_249(w_181_249, w_070_179, w_137_085);
  nand2 I181_265(w_181_265, w_032_312, w_089_006);
  and2 I182_002(w_182_002, w_067_175, w_141_056);
  not1 I182_004(w_182_004, w_005_121);
  or2  I182_005(w_182_005, w_082_053, w_005_026);
  nand2 I182_007(w_182_007, w_032_136, w_133_313);
  nand2 I182_009(w_182_009, w_015_642, w_136_049);
  nand2 I182_010(w_182_010, w_103_056, w_014_260);
  not1 I182_011(w_182_011, w_085_084);
  nand2 I182_013(w_182_013, w_077_000, w_105_331);
  or2  I182_015(w_182_015, w_005_015, w_127_008);
  and2 I182_016(w_182_016, w_014_281, w_083_163);
  and2 I182_017(w_182_017, w_004_061, w_074_320);
  or2  I182_018(w_182_018, w_159_048, w_135_163);
  and2 I182_021(w_182_021, w_023_062, w_030_352);
  nand2 I182_023(w_182_023, w_146_309, w_071_031);
  or2  I182_024(w_182_024, w_152_428, w_093_393);
  and2 I182_025(w_182_025, w_148_015, w_042_062);
  nand2 I182_026(w_182_026, w_136_031, w_054_148);
  or2  I183_005(w_183_005, w_008_459, w_129_256);
  or2  I183_008(w_183_008, w_148_609, w_077_409);
  nand2 I183_011(w_183_011, w_044_159, w_094_195);
  and2 I183_018(w_183_018, w_074_176, w_150_056);
  nand2 I183_025(w_183_025, w_037_103, w_034_065);
  and2 I183_031(w_183_031, w_166_219, w_173_016);
  and2 I183_039(w_183_039, w_162_008, w_112_084);
  and2 I183_041(w_183_041, w_136_013, w_076_087);
  not1 I183_073(w_183_073, w_035_050);
  and2 I183_092(w_183_092, w_143_076, w_040_630);
  or2  I183_103(w_183_103, w_128_327, w_119_082);
  or2  I183_111(w_183_111, w_176_110, w_142_442);
  and2 I183_118(w_183_118, w_000_292, w_029_051);
  nand2 I183_119(w_183_119, w_034_008, w_095_057);
  or2  I183_131(w_183_131, w_095_026, w_081_013);
  not1 I183_133(w_183_133, w_019_017);
  or2  I183_139(w_183_139, w_020_430, w_074_179);
  not1 I183_164(w_183_164, w_073_413);
  and2 I183_183(w_183_183, w_131_073, w_182_017);
  and2 I183_193(w_183_193, w_009_308, w_102_042);
  not1 I183_194(w_183_194, w_176_080);
  not1 I183_202(w_183_202, w_063_073);
  nand2 I183_243(w_183_243, w_122_126, w_029_070);
  nand2 I183_244(w_183_244, w_094_083, w_117_079);
  nand2 I183_270(w_183_270, w_098_052, w_139_009);
  and2 I184_000(w_184_000, w_122_072, w_135_438);
  nand2 I184_007(w_184_007, w_011_113, w_146_071);
  not1 I184_011(w_184_011, w_136_002);
  and2 I184_019(w_184_019, w_008_356, w_046_712);
  not1 I184_025(w_184_025, w_162_003);
  and2 I184_029(w_184_029, w_055_059, w_100_085);
  and2 I184_032(w_184_032, w_105_016, w_055_200);
  or2  I184_033(w_184_033, w_014_214, w_121_045);
  or2  I184_038(w_184_038, w_098_053, w_021_137);
  and2 I184_041(w_184_041, w_171_124, w_003_048);
  not1 I184_049(w_184_049, w_073_734);
  and2 I184_052(w_184_052, w_034_050, w_049_290);
  and2 I184_056(w_184_056, w_023_034, w_114_106);
  or2  I184_065(w_184_065, w_008_275, w_044_013);
  not1 I184_073(w_184_073, w_021_140);
  or2  I184_112(w_184_112, w_105_213, w_027_139);
  and2 I184_130(w_184_130, w_060_080, w_106_069);
  and2 I184_132(w_184_132, w_068_086, w_157_021);
  and2 I185_023(w_185_023, w_140_165, w_010_488);
  nand2 I185_027(w_185_027, w_109_284, w_087_069);
  nand2 I185_039(w_185_039, w_041_106, w_144_061);
  or2  I185_049(w_185_049, w_080_086, w_089_232);
  not1 I185_059(w_185_059, w_089_215);
  nand2 I185_069(w_185_069, w_175_167, w_085_161);
  and2 I185_072(w_185_072, w_134_405, w_150_231);
  or2  I185_076(w_185_076, w_094_376, w_142_792);
  or2  I185_090(w_185_090, w_083_021, w_155_508);
  or2  I185_094(w_185_094, w_166_010, w_064_130);
  not1 I185_100(w_185_100, w_078_497);
  not1 I185_103(w_185_103, w_007_152);
  or2  I185_104(w_185_104, w_078_093, w_127_041);
  nand2 I185_108(w_185_108, w_070_389, w_170_017);
  nand2 I185_109(w_185_109, w_000_569, w_009_064);
  not1 I185_112(w_185_112, w_021_055);
  and2 I185_130(w_185_130, w_147_097, w_020_034);
  not1 I185_137(w_185_137, w_062_643);
  not1 I185_140(w_185_140, w_095_002);
  or2  I185_185(w_185_185, w_093_178, w_153_057);
  not1 I185_198(w_185_198, w_122_020);
  not1 I185_202(w_185_202, w_090_415);
  nand2 I185_209(w_185_209, w_147_203, w_086_175);
  or2  I185_218(w_185_220, w_185_219, w_046_232);
  and2 I185_219(w_185_221, w_044_048, w_185_220);
  or2  I185_220(w_185_222, w_185_221, w_160_673);
  or2  I185_221(w_185_223, w_141_143, w_185_222);
  nand2 I185_222(w_185_224, w_185_223, w_034_004);
  and2 I185_223(w_185_225, w_085_353, w_185_224);
  nand2 I185_224(w_185_226, w_124_134, w_185_225);
  nand2 I185_225(w_185_227, w_066_584, w_185_226);
  not1 I185_226(w_185_228, w_185_227);
  and2 I185_227(w_185_229, w_185_228, w_069_237);
  nand2 I185_228(w_185_219, w_185_229, w_112_144);
  or2  I186_042(w_186_042, w_110_362, w_039_033);
  not1 I186_055(w_186_055, w_087_162);
  nand2 I186_084(w_186_084, w_136_058, w_063_432);
  and2 I186_093(w_186_093, w_163_567, w_180_026);
  not1 I186_095(w_186_095, w_003_025);
  nand2 I186_099(w_186_099, w_015_431, w_082_502);
  not1 I186_131(w_186_131, w_065_060);
  and2 I186_140(w_186_140, w_099_150, w_049_389);
  not1 I186_177(w_186_177, w_132_077);
  nand2 I186_197(w_186_197, w_142_603, w_121_209);
  or2  I186_205(w_186_205, w_161_155, w_041_038);
  and2 I186_208(w_186_208, w_024_009, w_022_186);
  nand2 I186_212(w_186_212, w_055_088, w_118_082);
  or2  I186_223(w_186_223, w_167_122, w_168_147);
  nand2 I186_231(w_186_231, w_063_250, w_001_032);
  or2  I186_235(w_186_235, w_114_152, w_043_032);
  nand2 I186_257(w_186_257, w_155_145, w_149_506);
  not1 I186_262(w_186_262, w_107_329);
  nand2 I186_295(w_186_295, w_138_100, w_043_047);
  and2 I186_322(w_186_322, w_128_010, w_029_020);
  nand2 I186_336(w_186_336, w_059_278, w_065_555);
  or2  I186_361(w_186_361, w_185_094, w_108_057);
  or2  I186_440(w_186_440, w_156_342, w_046_467);
  nand2 I186_450(w_186_450, w_173_004, w_003_026);
  or2  I186_467(w_186_467, w_122_035, w_068_081);
  not1 I186_537(w_186_537, w_052_043);
  and2 I186_575(w_185_231, w_171_578, w_185_219);
  nand2 I187_001(w_187_001, w_059_550, w_008_757);
  not1 I187_002(w_187_002, w_185_231);
  or2  I187_004(w_187_004, w_180_009, w_106_105);
  not1 I187_006(w_187_006, w_139_024);
  nand2 I187_009(w_187_009, w_001_026, w_084_028);
  and2 I187_010(w_187_010, w_162_003, w_161_160);
  nand2 I187_011(w_187_011, w_154_131, w_057_182);
  and2 I187_012(w_187_012, w_155_050, w_131_113);
  and2 I187_013(w_187_013, w_125_138, w_160_049);
  and2 I187_014(w_187_014, w_070_209, w_009_076);
  nand2 I187_015(w_187_015, w_109_114, w_067_010);
  not1 I187_016(w_187_016, w_047_291);
  and2 I187_017(w_187_017, w_021_004, w_117_060);
  and2 I187_019(w_187_019, w_137_045, w_116_192);
  nand2 I187_020(w_187_020, w_089_289, w_170_282);
  nand2 I187_023(w_187_023, w_021_273, w_068_337);
  or2  I187_026(w_187_026, w_065_338, w_095_056);
  not1 I187_028(w_187_028, w_169_303);
  nand2 I187_029(w_187_029, w_143_568, w_097_105);
  and2 I187_030(w_187_030, w_165_088, w_159_029);
  not1 I187_032(w_187_032, w_167_031);
  and2 I187_033(w_187_033, w_087_243, w_052_039);
  or2  I187_039(w_187_039, w_023_122, w_067_255);
  and2 I187_041(w_187_041, w_142_040, w_052_024);
  or2  I188_003(w_188_003, w_173_002, w_171_450);
  or2  I188_007(w_188_007, w_121_160, w_093_060);
  and2 I188_036(w_188_036, w_156_100, w_171_495);
  nand2 I188_039(w_188_039, w_012_037, w_151_108);
  and2 I188_062(w_188_062, w_169_273, w_008_241);
  and2 I188_091(w_188_091, w_114_144, w_095_036);
  not1 I188_107(w_188_107, w_062_483);
  not1 I188_146(w_188_146, w_003_065);
  and2 I188_158(w_188_158, w_175_417, w_012_345);
  nand2 I188_184(w_188_184, w_052_012, w_045_067);
  nand2 I188_225(w_188_225, w_016_005, w_110_277);
  and2 I188_281(w_188_281, w_134_066, w_049_162);
  not1 I188_393(w_188_393, w_129_278);
  and2 I188_437(w_188_437, w_109_003, w_079_052);
  nand2 I188_592(w_188_592, w_106_044, w_008_616);
  and2 I188_646(w_188_646, w_000_259, w_125_057);
  not1 I189_023(w_189_023, w_183_008);
  not1 I189_025(w_189_025, w_045_055);
  nand2 I189_026(w_189_026, w_118_099, w_131_304);
  and2 I189_056(w_189_056, w_052_011, w_084_044);
  and2 I189_092(w_189_092, w_151_284, w_036_299);
  nand2 I189_119(w_189_119, w_120_244, w_083_138);
  nand2 I189_157(w_189_157, w_003_075, w_084_039);
  or2  I189_175(w_189_175, w_011_099, w_150_150);
  not1 I189_220(w_189_220, w_058_321);
  or2  I189_298(w_189_298, w_074_258, w_061_105);
  or2  I189_319(w_189_319, w_100_096, w_134_251);
  or2  I189_367(w_189_367, w_008_208, w_154_009);
  and2 I189_443(w_189_443, w_060_123, w_067_024);
  nand2 I189_445(w_189_445, w_110_459, w_065_426);
  or2  I189_446(w_189_446, w_096_005, w_004_500);
  nand2 I189_463(w_189_463, w_161_326, w_013_443);
  nand2 I189_471(w_189_471, w_130_212, w_093_409);
  or2  I189_478(w_189_478, w_056_108, w_039_280);
  nand2 I189_484(w_189_484, w_139_013, w_096_003);
  or2  I189_513(w_189_513, w_121_121, w_067_347);
  nand2 I189_546(w_189_546, w_085_152, w_090_380);
  or2  I189_619(w_189_621, w_189_620, w_061_467);
  nand2 I189_620(w_189_622, w_189_621, w_069_081);
  and2 I189_621(w_189_623, w_162_013, w_189_622);
  or2  I189_622(w_189_620, w_015_449, w_189_623);
  or2  I190_000(w_190_000, w_041_511, w_047_330);
  or2  I190_001(w_190_001, w_116_238, w_047_305);
  not1 I190_005(w_190_005, w_170_015);
  nand2 I190_008(w_190_008, w_065_603, w_110_282);
  and2 I190_009(w_190_009, w_016_002, w_095_000);
  nand2 I190_014(w_190_014, w_115_179, w_051_195);
  and2 I190_029(w_190_029, w_146_090, w_096_003);
  or2  I190_034(w_190_034, w_113_033, w_115_018);
  or2  I190_036(w_190_036, w_061_188, w_065_569);
  and2 I190_040(w_190_040, w_123_481, w_081_018);
  not1 I190_041(w_190_041, w_099_278);
  and2 I190_053(w_190_053, w_063_223, w_172_000);
  not1 I190_066(w_190_066, w_011_634);
  nand2 I190_067(w_190_067, w_152_118, w_046_414);
  not1 I190_073(w_190_073, w_147_175);
  or2  I190_074(w_190_074, w_109_293, w_044_373);
  or2  I190_093(w_190_093, w_043_047, w_023_090);
  or2  I190_095(w_190_095, w_076_362, w_131_147);
  not1 I190_096(w_190_096, w_138_104);
  nand2 I190_100(w_190_100, w_126_038, w_034_060);
  nand2 I190_103(w_190_103, w_170_040, w_184_000);
  nand2 I190_112(w_190_112, w_077_420, w_007_160);
  or2  I190_116(w_190_116, w_166_041, w_110_047);
  not1 I191_008(w_191_008, w_061_172);
  not1 I191_011(w_191_011, w_148_553);
  and2 I191_026(w_191_026, w_068_131, w_166_268);
  nand2 I191_027(w_191_027, w_160_245, w_020_108);
  or2  I191_033(w_191_033, w_084_018, w_103_248);
  or2  I191_034(w_191_034, w_134_451, w_080_369);
  not1 I191_045(w_191_045, w_080_173);
  and2 I191_047(w_191_047, w_042_117, w_115_240);
  and2 I191_051(w_191_051, w_162_025, w_076_140);
  not1 I191_052(w_191_052, w_156_041);
  and2 I191_062(w_191_062, w_091_081, w_119_087);
  nand2 I191_065(w_191_065, w_177_024, w_002_472);
  not1 I191_069(w_191_069, w_132_333);
  or2  I191_074(w_191_074, w_039_073, w_024_028);
  not1 I191_076(w_191_076, w_139_004);
  and2 I191_082(w_191_082, w_173_005, w_023_162);
  not1 I191_092(w_191_092, w_177_399);
  nand2 I191_134(w_191_134, w_016_006, w_005_120);
  not1 I191_136(w_191_136, w_095_027);
  nand2 I191_163(w_191_163, w_102_025, w_140_190);
  not1 I191_210(w_191_210, w_092_471);
  nand2 I191_215(w_191_215, w_033_322, w_026_606);
  nand2 I191_229(w_191_229, w_035_031, w_170_250);
  and2 I191_232(w_191_232, w_049_189, w_113_250);
  or2  I191_240(w_191_240, w_163_574, w_017_191);
  not1 I191_245(w_191_245, w_162_021);
  or2  I191_262(w_191_262, w_070_510, w_102_333);
  and2 I191_275(w_191_275, w_022_053, w_042_121);
  and2 I191_286(w_191_286, w_054_146, w_011_490);
  or2  I191_306(w_191_306, w_152_161, w_066_348);
  and2 I191_309(w_191_309, w_026_544, w_187_033);
  and2 I191_331(w_191_331, w_166_115, w_171_412);
  or2  I191_336(w_191_336, w_010_124, w_109_131);
  nand2 I191_362(w_191_362, w_147_118, w_002_024);
  or2  I192_008(w_192_008, w_099_172, w_132_155);
  or2  I192_009(w_192_009, w_096_005, w_091_088);
  not1 I192_010(w_192_010, w_059_462);
  not1 I192_017(w_192_017, w_064_310);
  or2  I192_019(w_192_019, w_067_211, w_063_088);
  not1 I192_031(w_192_031, w_071_209);
  not1 I192_041(w_192_041, w_178_054);
  nand2 I192_045(w_192_045, w_088_041, w_000_308);
  or2  I192_059(w_192_059, w_045_212, w_121_058);
  nand2 I192_063(w_192_063, w_087_149, w_044_030);
  not1 I192_065(w_192_065, w_043_018);
  not1 I192_079(w_192_079, w_032_478);
  nand2 I192_082(w_192_082, w_143_116, w_103_015);
  nand2 I192_099(w_192_099, w_001_004, w_132_031);
  or2  I192_113(w_192_113, w_050_045, w_010_225);
  or2  I192_114(w_192_114, w_068_221, w_038_467);
  not1 I192_119(w_192_119, w_154_093);
  or2  I192_134(w_192_134, w_123_174, w_060_359);
  and2 I192_138(w_192_138, w_114_112, w_073_514);
  or2  I192_145(w_192_145, w_071_300, w_191_008);
  not1 I192_146(w_192_146, w_102_252);
  nand2 I192_148(w_192_148, w_006_216, w_052_006);
  not1 I192_153(w_192_153, w_067_201);
  or2  I192_163(w_192_163, w_191_051, w_018_018);
  not1 I192_164(w_192_164, w_005_077);
  not1 I192_165(w_192_165, w_112_145);
  nand2 I192_172(w_192_172, w_097_090, w_150_003);
  and2 I192_175(w_192_175, w_168_380, w_104_273);
  not1 I192_176(w_192_176, w_105_241);
  and2 I192_179(w_192_179, w_169_296, w_185_100);
  nand2 I192_189(w_192_189, w_173_017, w_069_236);
  nand2 I192_195(w_192_197, w_192_196, w_002_522);
  and2 I192_196(w_192_198, w_104_280, w_192_197);
  or2  I192_197(w_192_199, w_056_609, w_192_198);
  nand2 I192_198(w_192_200, w_192_199, w_128_233);
  and2 I192_199(w_192_201, w_059_248, w_192_200);
  and2 I192_200(w_192_202, w_152_073, w_192_201);
  not1 I192_201(w_192_203, w_192_202);
  or2  I192_202(w_192_204, w_072_053, w_192_203);
  and2 I192_203(w_192_205, w_192_204, w_160_667);
  and2 I192_204(w_192_206, w_004_220, w_192_205);
  and2 I192_205(w_192_207, w_192_206, w_058_148);
  and2 I192_206(w_192_196, w_192_207, w_067_133);
  or2  I193_006(w_193_006, w_032_395, w_042_305);
  or2  I193_014(w_193_014, w_067_126, w_143_004);
  nand2 I193_021(w_193_021, w_146_057, w_155_290);
  and2 I193_033(w_193_033, w_035_115, w_141_059);
  or2  I193_067(w_193_067, w_083_043, w_142_095);
  and2 I193_080(w_193_080, w_056_692, w_081_012);
  or2  I193_085(w_193_085, w_104_009, w_019_000);
  or2  I193_087(w_193_087, w_153_038, w_095_004);
  nand2 I193_091(w_193_091, w_163_132, w_178_043);
  nand2 I193_097(w_193_097, w_058_447, w_025_139);
  nand2 I193_106(w_193_106, w_032_076, w_017_112);
  or2  I193_131(w_193_131, w_150_333, w_012_028);
  and2 I193_136(w_193_136, w_139_009, w_003_057);
  nand2 I193_137(w_193_137, w_133_362, w_020_378);
  nand2 I193_151(w_193_151, w_178_036, w_087_247);
  and2 I193_169(w_193_169, w_080_257, w_172_041);
  or2  I193_183(w_193_183, w_007_143, w_103_264);
  and2 I193_184(w_193_184, w_170_248, w_152_008);
  nand2 I193_190(w_193_190, w_026_711, w_063_173);
  or2  I193_199(w_193_199, w_123_036, w_024_026);
  nand2 I193_233(w_193_233, w_135_136, w_025_026);
  nand2 I193_272(w_193_272, w_024_404, w_019_005);
  not1 I193_296(w_193_296, w_061_062);
  or2  I193_299(w_193_299, w_114_226, w_090_542);
  nand2 I193_312(w_193_312, w_091_153, w_085_070);
  or2  I193_327(w_193_327, w_015_091, w_039_518);
  not1 I193_345(w_193_345, w_014_221);
  not1 I193_350(w_193_350, w_040_044);
  not1 I194_021(w_194_021, w_148_447);
  nand2 I194_057(w_194_057, w_038_549, w_163_225);
  and2 I194_077(w_194_077, w_010_216, w_046_698);
  and2 I194_078(w_194_078, w_066_154, w_067_356);
  nand2 I194_096(w_194_096, w_138_073, w_113_181);
  and2 I194_098(w_194_098, w_009_229, w_116_407);
  nand2 I194_102(w_194_102, w_010_159, w_022_365);
  nand2 I194_117(w_194_117, w_017_541, w_082_541);
  nand2 I194_132(w_194_132, w_140_031, w_068_349);
  nand2 I194_136(w_194_136, w_131_566, w_086_270);
  or2  I194_142(w_194_142, w_107_097, w_004_453);
  and2 I194_170(w_194_170, w_006_086, w_057_262);
  nand2 I194_173(w_194_173, w_157_065, w_027_122);
  or2  I194_174(w_194_174, w_155_103, w_004_389);
  and2 I194_178(w_194_178, w_038_589, w_113_318);
  nand2 I194_187(w_194_187, w_075_137, w_080_212);
  not1 I194_221(w_194_221, w_032_448);
  not1 I194_238(w_194_238, w_080_245);
  not1 I194_241(w_194_241, w_081_007);
  and2 I194_246(w_194_246, w_059_501, w_012_110);
  and2 I194_262(w_194_262, w_146_005, w_061_057);
  not1 I194_298(w_194_298, w_076_036);
  and2 I194_304(w_194_304, w_182_015, w_154_046);
  and2 I194_314(w_194_314, w_147_165, w_157_032);
  and2 I194_325(w_194_325, w_011_426, w_129_198);
  and2 I195_003(w_195_003, w_115_162, w_120_569);
  not1 I195_006(w_195_006, w_149_082);
  nand2 I195_007(w_195_007, w_019_014, w_015_585);
  not1 I195_023(w_195_023, w_114_106);
  or2  I195_030(w_195_030, w_076_115, w_109_285);
  or2  I195_035(w_195_035, w_111_023, w_020_092);
  and2 I195_044(w_195_044, w_084_006, w_097_224);
  or2  I195_046(w_195_046, w_084_020, w_175_026);
  and2 I195_054(w_195_054, w_089_191, w_170_310);
  and2 I195_067(w_195_067, w_024_280, w_185_039);
  not1 I195_072(w_195_072, w_013_062);
  and2 I195_074(w_195_074, w_121_039, w_185_112);
  and2 I195_075(w_195_075, w_129_072, w_057_228);
  and2 I195_081(w_195_081, w_154_112, w_056_723);
  or2  I195_084(w_195_084, w_053_135, w_003_055);
  not1 I195_100(w_195_100, w_053_071);
  not1 I195_107(w_195_107, w_086_024);
  not1 I195_121(w_195_121, w_155_252);
  or2  I195_128(w_195_128, w_031_556, w_049_116);
  nand2 I195_129(w_195_129, w_087_215, w_121_189);
  and2 I195_139(w_195_139, w_012_324, w_152_221);
  or2  I195_140(w_195_140, w_087_051, w_097_504);
  not1 I195_141(w_195_141, w_030_325);
  or2  I195_148(w_195_148, w_022_196, w_113_047);
  or2  I195_177(w_195_177, w_183_118, w_110_039);
  nand2 I195_194(w_195_194, w_126_013, w_000_123);
  not1 I195_205(w_195_205, w_093_178);
  nand2 I195_208(w_195_208, w_035_017, w_160_426);
  not1 I195_209(w_195_209, w_185_076);
  nand2 I195_216(w_195_216, w_039_050, w_180_009);
  or2  I195_228(w_195_228, w_146_044, w_131_285);
  or2  I195_232(w_195_232, w_154_080, w_147_168);
  not1 I195_233(w_195_233, w_108_166);
  nand2 I195_236(w_195_236, w_139_014, w_154_131);
  nand2 I195_241(w_195_241, w_104_021, w_037_248);
  nand2 I196_007(w_196_007, w_055_082, w_010_715);
  nand2 I196_016(w_196_016, w_096_002, w_064_125);
  or2  I196_023(w_196_023, w_017_357, w_065_040);
  not1 I196_040(w_196_040, w_117_038);
  nand2 I196_072(w_196_072, w_067_125, w_193_184);
  or2  I196_075(w_196_075, w_112_182, w_092_480);
  and2 I196_079(w_196_079, w_052_044, w_068_170);
  and2 I196_095(w_196_095, w_190_008, w_043_003);
  nand2 I196_101(w_196_101, w_014_068, w_043_009);
  nand2 I196_111(w_196_111, w_065_425, w_166_282);
  and2 I196_136(w_196_136, w_151_259, w_069_088);
  and2 I196_141(w_196_141, w_002_626, w_093_041);
  or2  I196_149(w_196_149, w_079_055, w_030_125);
  nand2 I196_154(w_196_154, w_113_146, w_187_020);
  and2 I196_163(w_196_163, w_179_203, w_195_075);
  or2  I196_173(w_196_173, w_000_716, w_140_093);
  not1 I196_196(w_196_196, w_186_467);
  or2  I196_210(w_196_210, w_101_247, w_118_104);
  not1 I196_212(w_196_212, w_103_210);
  not1 I196_217(w_196_217, w_013_540);
  and2 I196_254(w_196_254, w_026_669, w_032_025);
  or2  I197_017(w_197_017, w_098_016, w_173_030);
  or2  I197_060(w_197_060, w_149_466, w_074_251);
  nand2 I197_064(w_197_064, w_019_004, w_114_015);
  and2 I197_098(w_197_098, w_113_209, w_164_291);
  nand2 I197_114(w_197_114, w_063_361, w_102_345);
  or2  I197_141(w_197_141, w_171_408, w_063_142);
  not1 I197_146(w_197_146, w_028_078);
  or2  I197_152(w_197_152, w_076_255, w_104_162);
  nand2 I197_160(w_197_160, w_017_236, w_090_232);
  or2  I197_161(w_197_161, w_072_235, w_091_119);
  and2 I197_194(w_197_194, w_138_205, w_140_137);
  not1 I197_223(w_197_223, w_138_250);
  nand2 I197_228(w_197_228, w_143_501, w_132_395);
  and2 I197_247(w_197_247, w_172_053, w_122_060);
  nand2 I197_248(w_197_248, w_048_002, w_179_620);
  or2  I197_312(w_197_312, w_041_532, w_111_091);
  and2 I197_396(w_197_396, w_115_134, w_101_176);
  not1 I197_445(w_197_445, w_172_024);
  and2 I198_006(w_198_006, w_064_329, w_100_100);
  and2 I198_014(w_198_014, w_110_139, w_153_052);
  not1 I198_017(w_198_017, w_098_004);
  and2 I198_021(w_198_021, w_099_229, w_001_020);
  not1 I198_024(w_198_024, w_032_042);
  or2  I198_030(w_198_030, w_167_081, w_005_094);
  and2 I198_044(w_198_044, w_019_002, w_052_032);
  not1 I198_046(w_198_046, w_118_093);
  and2 I198_052(w_198_052, w_086_055, w_070_508);
  not1 I198_053(w_198_053, w_188_437);
  and2 I198_054(w_198_054, w_061_221, w_083_110);
  or2  I198_056(w_198_056, w_183_131, w_014_064);
  or2  I198_057(w_198_057, w_021_096, w_154_121);
  nand2 I198_059(w_198_059, w_116_077, w_013_044);
  or2  I198_060(w_198_060, w_004_265, w_045_271);
  nand2 I198_062(w_198_062, w_123_087, w_147_099);
  nand2 I198_076(w_198_076, w_120_578, w_123_053);
  not1 I198_078(w_198_078, w_025_121);
  not1 I199_040(w_199_040, w_154_096);
  or2  I199_048(w_199_048, w_090_536, w_016_006);
  and2 I199_054(w_199_054, w_057_004, w_101_258);
  or2  I199_073(w_199_073, w_066_182, w_170_212);
  nand2 I199_076(w_199_076, w_163_157, w_195_129);
  and2 I199_106(w_199_106, w_164_141, w_011_140);
  or2  I199_156(w_199_156, w_047_134, w_124_273);
  or2  I199_159(w_199_159, w_114_197, w_174_093);
  and2 I199_173(w_199_173, w_069_218, w_022_290);
  not1 I199_178(w_199_178, w_119_135);
  or2  I199_235(w_199_235, w_119_177, w_070_199);
  and2 I199_240(w_199_240, w_080_113, w_181_249);
  and2 I199_253(w_199_253, w_151_184, w_170_198);
  nand2 I199_266(w_199_266, w_154_119, w_042_180);
  or2  I199_267(w_199_267, w_144_169, w_178_095);
  not1 I199_280(w_199_280, w_181_118);
  nand2 I199_294(w_199_294, w_112_189, w_087_106);
  nand2 I199_338(w_199_338, w_089_155, w_139_006);
  not1 I199_373(w_199_373, w_141_002);
  nand2 I200_002(w_200_002, w_023_038, w_140_094);
  nand2 I200_005(w_200_005, w_016_006, w_165_025);
  nand2 I200_021(w_200_021, w_173_030, w_022_297);
  or2  I200_028(w_200_028, w_140_188, w_099_071);
  and2 I200_045(w_200_045, w_177_178, w_046_184);
  or2  I200_061(w_200_061, w_146_191, w_041_081);
  and2 I200_089(w_200_089, w_020_327, w_142_772);
  or2  I200_106(w_200_106, w_196_154, w_138_160);
  or2  I200_117(w_200_117, w_106_025, w_157_151);
  and2 I200_127(w_200_127, w_147_216, w_195_216);
  nand2 I200_128(w_200_128, w_189_056, w_109_374);
  not1 I200_178(w_200_178, w_095_057);
  not1 I200_183(w_200_183, w_085_219);
  and2 I200_188(w_200_188, w_085_059, w_120_169);
  nand2 I200_211(w_200_211, w_125_193, w_195_081);
  not1 I200_214(w_200_214, w_160_182);
  not1 I200_216(w_200_216, w_114_144);
  not1 I200_234(w_200_234, w_160_299);
  nand2 I200_254(w_200_254, w_121_199, w_186_042);
  and2 I200_282(w_200_282, w_109_217, w_094_271);
  nand2 I200_359(w_200_359, w_195_233, w_144_206);
  and2 I200_407(w_200_407, w_193_350, w_049_304);
  nand2 I200_429(w_200_429, w_165_028, w_067_353);
  and2 I200_436(w_200_436, w_127_015, w_159_080);
  or2  I200_440(w_200_440, w_004_264, w_183_018);
  not1 I200_448(w_200_448, w_005_073);
  or2  I200_498(w_200_498, w_108_095, w_082_128);
  or2  I201_007(w_201_007, w_037_132, w_086_095);
  not1 I201_009(w_201_009, w_043_000);
  not1 I201_026(w_201_026, w_140_074);
  and2 I201_027(w_201_027, w_190_014, w_062_308);
  and2 I201_035(w_201_035, w_054_490, w_130_049);
  not1 I201_057(w_201_057, w_091_143);
  not1 I201_062(w_201_062, w_019_001);
  and2 I201_081(w_201_081, w_079_045, w_043_042);
  or2  I201_141(w_201_141, w_168_152, w_011_249);
  or2  I201_148(w_201_148, w_196_210, w_020_466);
  not1 I201_174(w_201_174, w_194_142);
  or2  I201_190(w_201_190, w_174_098, w_056_033);
  and2 I201_193(w_201_193, w_064_312, w_055_103);
  and2 I201_203(w_201_203, w_020_577, w_163_228);
  and2 I201_226(w_201_226, w_132_204, w_178_005);
  or2  I201_268(w_201_268, w_130_033, w_153_009);
  nand2 I201_280(w_201_280, w_177_014, w_022_392);
  or2  I201_286(w_201_286, w_033_119, w_164_348);
  nand2 I201_346(w_201_346, w_144_190, w_021_068);
  nand2 I201_409(w_201_409, w_013_001, w_169_437);
  not1 I201_422(w_201_422, w_050_446);
  and2 I201_502(w_201_502, w_101_272, w_137_351);
  and2 I202_014(w_202_014, w_106_012, w_187_012);
  not1 I202_017(w_202_017, w_035_014);
  nand2 I202_022(w_202_022, w_040_019, w_160_699);
  and2 I202_029(w_202_029, w_079_050, w_139_010);
  and2 I202_033(w_202_033, w_128_417, w_074_128);
  nand2 I202_040(w_202_040, w_178_107, w_037_168);
  or2  I202_055(w_202_055, w_129_090, w_156_057);
  and2 I202_064(w_202_064, w_094_387, w_112_104);
  not1 I202_066(w_202_066, w_100_055);
  nand2 I202_077(w_202_077, w_101_135, w_154_051);
  nand2 I202_078(w_202_078, w_045_307, w_006_131);
  not1 I202_079(w_202_079, w_163_491);
  not1 I202_085(w_202_085, w_138_283);
  nand2 I202_089(w_202_089, w_160_580, w_198_060);
  or2  I202_095(w_202_095, w_135_196, w_144_006);
  or2  I202_105(w_202_105, w_129_133, w_080_202);
  and2 I202_111(w_202_111, w_009_353, w_070_109);
  and2 I202_116(w_202_116, w_137_183, w_150_041);
  not1 I202_119(w_202_119, w_152_108);
  or2  I202_149(w_202_149, w_153_073, w_187_029);
  not1 I202_153(w_202_153, w_154_120);
  or2  I202_165(w_202_165, w_081_004, w_050_537);
  not1 I202_184(w_202_184, w_195_046);
  not1 I202_186(w_202_186, w_027_170);
  not1 I202_196(w_202_196, w_097_179);
  not1 I202_198(w_202_198, w_155_076);
  and2 I202_218(w_202_218, w_080_464, w_085_306);
  nand2 I202_223(w_202_223, w_059_111, w_027_113);
  not1 I202_231(w_202_231, w_070_435);
  not1 I202_252(w_202_252, w_094_299);
  not1 I202_267(w_202_267, w_138_047);
  or2  I202_276(w_202_276, w_143_081, w_021_167);
  and2 I202_278(w_202_278, w_001_027, w_019_020);
  nand2 I202_286(w_202_286, w_014_041, w_039_088);
  or2  I202_292(w_202_292, w_141_016, w_032_239);
  not1 I202_295(w_202_295, w_080_433);
  and2 I203_015(w_203_015, w_028_413, w_144_447);
  and2 I203_016(w_203_016, w_191_262, w_175_083);
  not1 I203_027(w_203_027, w_104_370);
  and2 I203_032(w_203_032, w_182_009, w_124_109);
  not1 I203_045(w_203_045, w_141_012);
  nand2 I203_062(w_203_062, w_143_598, w_018_024);
  and2 I203_074(w_203_074, w_192_163, w_106_146);
  not1 I203_083(w_203_083, w_175_558);
  nand2 I203_090(w_203_090, w_069_089, w_202_079);
  or2  I203_143(w_203_143, w_194_298, w_051_326);
  or2  I203_184(w_203_184, w_193_136, w_092_154);
  not1 I203_198(w_203_198, w_112_056);
  not1 I203_246(w_203_246, w_010_544);
  nand2 I203_259(w_203_259, w_091_170, w_184_065);
  or2  I203_271(w_203_271, w_117_066, w_028_325);
  not1 I203_297(w_203_297, w_089_151);
  nand2 I203_339(w_203_339, w_077_292, w_188_158);
  or2  I203_368(w_203_368, w_192_148, w_144_185);
  not1 I203_375(w_203_375, w_120_612);
  or2  I203_430(w_203_430, w_171_176, w_058_330);
  and2 I203_433(w_203_433, w_137_202, w_003_044);
  not1 I203_444(w_203_444, w_128_130);
  not1 I203_473(w_203_473, w_060_025);
  not1 I203_478(w_203_478, w_005_119);
  not1 I204_011(w_204_011, w_202_153);
  nand2 I204_027(w_204_027, w_169_323, w_099_256);
  and2 I204_043(w_204_043, w_129_100, w_053_055);
  and2 I204_056(w_204_056, w_121_141, w_126_027);
  and2 I204_135(w_204_135, w_041_234, w_005_071);
  or2  I204_218(w_204_218, w_049_111, w_178_054);
  or2  I204_280(w_204_280, w_058_505, w_102_451);
  nand2 I204_323(w_204_323, w_070_210, w_089_126);
  and2 I204_386(w_204_386, w_013_509, w_117_054);
  nand2 I204_388(w_204_388, w_155_192, w_091_073);
  or2  I204_473(w_204_473, w_022_174, w_057_092);
  and2 I204_493(w_204_493, w_187_017, w_060_019);
  not1 I204_510(w_204_510, w_105_218);
  or2  I204_651(w_204_651, w_123_459, w_135_003);
  or2  I205_000(w_205_000, w_052_030, w_045_129);
  or2  I205_007(w_205_007, w_132_130, w_112_165);
  not1 I205_034(w_205_034, w_085_024);
  or2  I205_035(w_205_035, w_170_399, w_014_114);
  or2  I205_053(w_205_053, w_151_178, w_161_155);
  nand2 I205_066(w_205_066, w_145_012, w_190_095);
  or2  I205_076(w_205_076, w_028_126, w_041_276);
  not1 I205_122(w_205_122, w_082_142);
  or2  I205_153(w_205_153, w_055_138, w_022_351);
  not1 I205_173(w_205_173, w_069_173);
  not1 I205_186(w_205_186, w_088_036);
  nand2 I205_199(w_205_199, w_119_003, w_166_165);
  not1 I205_216(w_205_216, w_041_482);
  not1 I205_217(w_205_217, w_129_180);
  and2 I205_245(w_205_245, w_092_580, w_121_174);
  nand2 I205_285(w_205_285, w_043_042, w_172_049);
  or2  I205_309(w_205_309, w_114_036, w_100_038);
  nand2 I205_317(w_205_317, w_083_190, w_049_322);
  and2 I205_330(w_205_330, w_188_062, w_117_000);
  nand2 I205_353(w_205_353, w_027_064, w_137_235);
  not1 I205_367(w_205_367, w_010_188);
  or2  I205_453(w_205_453, w_087_160, w_181_058);
  nand2 I205_459(w_205_459, w_035_013, w_021_113);
  and2 I205_462(w_205_462, w_114_003, w_140_010);
  not1 I205_504(w_205_504, w_162_004);
  and2 I205_519(w_205_519, w_038_146, w_104_047);
  not1 I205_537(w_205_537, w_185_090);
  nand2 I206_002(w_206_002, w_046_436, w_137_034);
  or2  I206_009(w_206_009, w_037_263, w_037_076);
  not1 I206_010(w_206_010, w_016_002);
  and2 I206_038(w_206_038, w_094_336, w_044_574);
  not1 I206_046(w_206_046, w_180_002);
  or2  I206_047(w_206_047, w_045_197, w_158_002);
  nand2 I206_058(w_206_058, w_188_281, w_166_152);
  and2 I206_070(w_206_070, w_150_127, w_186_197);
  not1 I206_082(w_206_082, w_126_153);
  not1 I206_086(w_206_086, w_098_004);
  and2 I206_087(w_206_087, w_085_255, w_145_052);
  or2  I206_119(w_206_119, w_135_398, w_154_036);
  and2 I206_139(w_206_139, w_003_037, w_115_089);
  not1 I206_144(w_206_144, w_135_487);
  not1 I206_145(w_206_145, w_171_479);
  or2  I206_157(w_206_157, w_176_138, w_008_232);
  or2  I206_203(w_206_203, w_025_164, w_152_236);
  not1 I207_026(w_207_026, w_172_039);
  or2  I207_049(w_207_049, w_105_200, w_090_042);
  nand2 I207_050(w_207_050, w_166_076, w_067_154);
  and2 I207_069(w_207_069, w_104_091, w_051_275);
  not1 I207_086(w_207_086, w_093_088);
  not1 I207_110(w_207_110, w_158_004);
  or2  I207_119(w_207_119, w_154_065, w_160_074);
  nand2 I207_144(w_207_144, w_201_286, w_158_001);
  nand2 I207_152(w_207_152, w_023_162, w_044_290);
  or2  I207_189(w_207_189, w_204_388, w_042_156);
  not1 I207_198(w_207_198, w_015_478);
  not1 I207_202(w_207_202, w_102_421);
  or2  I207_233(w_207_233, w_164_266, w_142_421);
  and2 I207_263(w_207_263, w_202_077, w_131_040);
  not1 I207_378(w_207_378, w_179_768);
  and2 I207_463(w_207_463, w_060_027, w_187_041);
  or2  I207_468(w_207_468, w_017_197, w_146_044);
  nand2 I207_546(w_207_546, w_011_030, w_175_488);
  or2  I208_021(w_208_021, w_111_021, w_026_455);
  and2 I208_026(w_208_026, w_196_210, w_086_173);
  or2  I208_027(w_208_027, w_161_023, w_102_609);
  and2 I208_035(w_208_035, w_185_209, w_157_022);
  or2  I208_053(w_208_053, w_059_168, w_159_045);
  and2 I208_072(w_208_072, w_087_182, w_118_061);
  and2 I208_083(w_208_083, w_166_305, w_199_173);
  not1 I208_122(w_208_122, w_183_005);
  and2 I208_133(w_208_133, w_091_157, w_063_483);
  or2  I208_161(w_208_161, w_129_095, w_147_029);
  nand2 I208_169(w_208_169, w_127_018, w_020_018);
  nand2 I208_175(w_208_175, w_162_024, w_197_396);
  or2  I208_214(w_208_214, w_073_143, w_029_026);
  and2 I208_225(w_208_225, w_142_101, w_108_087);
  and2 I208_231(w_208_231, w_130_260, w_064_214);
  not1 I208_238(w_208_238, w_089_111);
  or2  I208_244(w_208_244, w_178_067, w_179_507);
  not1 I208_259(w_208_259, w_077_262);
  and2 I208_268(w_208_268, w_025_003, w_098_058);
  nand2 I208_273(w_208_273, w_153_067, w_122_012);
  nand2 I208_277(w_208_277, w_155_034, w_023_091);
  or2  I208_354(w_208_354, w_061_256, w_093_162);
  nand2 I208_400(w_208_400, w_154_036, w_138_214);
  nand2 I208_408(w_208_408, w_195_030, w_159_074);
  and2 I209_007(w_209_007, w_025_145, w_031_103);
  or2  I209_012(w_209_012, w_194_246, w_163_266);
  and2 I209_018(w_209_018, w_047_124, w_057_076);
  or2  I209_033(w_209_033, w_141_175, w_098_020);
  nand2 I209_043(w_209_043, w_030_327, w_106_138);
  and2 I209_054(w_209_054, w_068_348, w_040_432);
  nand2 I209_057(w_209_057, w_120_051, w_042_432);
  or2  I209_062(w_209_062, w_098_009, w_188_646);
  and2 I209_063(w_209_063, w_153_060, w_195_074);
  nand2 I209_065(w_209_065, w_006_053, w_127_038);
  not1 I209_087(w_209_087, w_106_012);
  and2 I209_106(w_209_106, w_087_154, w_027_204);
  or2  I209_139(w_209_139, w_161_071, w_072_001);
  and2 I209_140(w_209_140, w_138_037, w_162_003);
  or2  I209_145(w_209_145, w_048_007, w_164_204);
  not1 I209_176(w_209_176, w_031_070);
  not1 I209_182(w_209_182, w_108_073);
  or2  I209_209(w_209_209, w_046_575, w_192_045);
  or2  I209_255(w_209_255, w_048_017, w_117_074);
  not1 I209_263(w_209_263, w_077_022);
  not1 I209_281(w_209_281, w_086_189);
  nand2 I209_299(w_209_299, w_080_131, w_150_068);
  not1 I209_314(w_209_314, w_026_466);
  or2  I209_322(w_209_322, w_059_396, w_044_652);
  or2  I209_342(w_209_342, w_189_478, w_036_244);
  or2  I209_345(w_209_345, w_073_209, w_070_568);
  not1 I210_003(w_210_003, w_152_601);
  nand2 I210_014(w_210_014, w_127_052, w_208_268);
  and2 I210_019(w_210_019, w_160_706, w_034_054);
  not1 I210_020(w_210_020, w_061_065);
  nand2 I210_028(w_210_028, w_199_054, w_181_048);
  and2 I210_030(w_210_030, w_032_496, w_139_023);
  not1 I210_040(w_210_040, w_109_127);
  and2 I210_044(w_210_044, w_033_231, w_053_158);
  or2  I210_061(w_210_061, w_011_550, w_104_197);
  nand2 I210_064(w_210_064, w_052_045, w_114_176);
  not1 I210_093(w_210_093, w_183_164);
  not1 I210_098(w_210_098, w_087_127);
  not1 I210_101(w_210_101, w_062_239);
  or2  I210_102(w_210_102, w_194_096, w_172_048);
  not1 I210_107(w_210_107, w_057_250);
  nand2 I210_124(w_210_124, w_190_103, w_050_257);
  nand2 I210_132(w_210_132, w_151_302, w_095_038);
  nand2 I210_139(w_210_139, w_004_076, w_207_463);
  or2  I210_142(w_210_142, w_024_483, w_120_126);
  nand2 I211_003(w_211_003, w_191_092, w_122_021);
  not1 I211_004(w_211_004, w_071_058);
  and2 I211_005(w_211_005, w_070_579, w_020_554);
  nand2 I211_006(w_211_006, w_063_194, w_203_246);
  and2 I211_012(w_211_012, w_040_616, w_182_023);
  nand2 I211_014(w_211_014, w_205_317, w_183_103);
  and2 I211_017(w_211_017, w_013_154, w_186_295);
  nand2 I211_018(w_211_018, w_116_412, w_138_157);
  and2 I211_019(w_211_019, w_178_099, w_014_088);
  nand2 I211_021(w_211_021, w_016_004, w_024_286);
  not1 I211_023(w_211_023, w_106_129);
  not1 I211_026(w_211_026, w_202_218);
  not1 I211_027(w_211_027, w_049_267);
  not1 I211_028(w_211_028, w_181_002);
  nand2 I211_033(w_211_033, w_101_294, w_016_004);
  and2 I211_034(w_211_034, w_161_079, w_146_210);
  or2  I211_036(w_211_036, w_080_319, w_125_586);
  not1 I211_037(w_211_037, w_110_041);
  and2 I211_038(w_211_040, w_211_039, w_112_180);
  and2 I211_039(w_211_041, w_002_046, w_211_040);
  or2  I211_040(w_211_042, w_211_041, w_082_240);
  not1 I211_041(w_211_043, w_211_042);
  nand2 I211_042(w_211_044, w_211_043, w_042_127);
  not1 I211_043(w_211_045, w_211_044);
  not1 I211_044(w_211_046, w_211_045);
  nand2 I211_045(w_211_047, w_211_046, w_155_109);
  not1 I211_046(w_211_048, w_211_047);
  and2 I211_047(w_211_049, w_149_207, w_211_048);
  or2  I211_048(w_211_039, w_211_049, w_205_459);
  nand2 I212_003(w_212_003, w_194_174, w_042_423);
  nand2 I212_006(w_212_006, w_099_262, w_079_015);
  nand2 I212_009(w_212_009, w_175_025, w_174_088);
  or2  I212_019(w_212_019, w_119_149, w_084_045);
  and2 I212_034(w_212_034, w_032_109, w_058_607);
  not1 I212_048(w_212_048, w_094_159);
  nand2 I212_052(w_212_052, w_074_259, w_066_061);
  not1 I212_061(w_212_061, w_209_057);
  nand2 I212_064(w_212_064, w_144_219, w_056_551);
  and2 I212_067(w_212_067, w_163_428, w_210_064);
  and2 I212_073(w_212_073, w_147_113, w_148_043);
  or2  I212_087(w_212_087, w_163_416, w_120_167);
  and2 I212_092(w_212_092, w_058_287, w_186_197);
  and2 I212_117(w_212_117, w_119_119, w_007_454);
  nand2 I212_120(w_212_120, w_044_658, w_088_011);
  not1 I212_124(w_212_124, w_142_517);
  not1 I212_162(w_212_162, w_114_058);
  not1 I212_163(w_212_163, w_210_102);
  not1 I212_165(w_212_165, w_106_123);
  nand2 I212_170(w_212_170, w_132_087, w_137_190);
  and2 I212_182(w_212_182, w_173_030, w_208_244);
  and2 I212_189(w_212_189, w_055_057, w_205_153);
  and2 I212_190(w_212_190, w_161_472, w_070_028);
  not1 I212_202(w_212_202, w_101_139);
  or2  I212_204(w_212_204, w_135_488, w_057_137);
  nand2 I212_218(w_212_218, w_134_204, w_076_046);
  and2 I212_226(w_212_226, w_116_153, w_090_191);
  and2 I212_229(w_211_051, w_075_013, w_211_039);
  and2 I213_005(w_213_005, w_077_052, w_116_345);
  or2  I213_007(w_213_007, w_009_056, w_006_207);
  nand2 I213_013(w_213_013, w_173_030, w_020_068);
  or2  I213_015(w_213_015, w_026_061, w_030_168);
  not1 I213_017(w_213_017, w_098_059);
  and2 I213_046(w_213_046, w_164_023, w_096_002);
  or2  I213_052(w_213_052, w_132_219, w_004_017);
  or2  I213_070(w_213_070, w_050_121, w_191_027);
  not1 I213_078(w_213_078, w_196_163);
  nand2 I213_079(w_213_079, w_043_015, w_193_233);
  not1 I213_085(w_213_085, w_011_117);
  or2  I213_086(w_213_086, w_055_080, w_107_121);
  nand2 I213_179(w_213_179, w_151_034, w_071_020);
  not1 I213_194(w_213_194, w_194_078);
  nand2 I213_241(w_213_241, w_180_024, w_040_475);
  nand2 I213_303(w_213_303, w_072_144, w_120_353);
  or2  I213_315(w_213_315, w_102_181, w_134_448);
  or2  I213_339(w_213_339, w_125_297, w_022_234);
  or2  I213_358(w_213_358, w_040_514, w_015_458);
  or2  I213_368(w_213_368, w_116_260, w_027_020);
  not1 I213_392(w_213_392, w_115_131);
  not1 I213_414(w_213_414, w_129_111);
  nand2 I213_419(w_213_419, w_163_519, w_038_065);
  not1 I213_466(w_213_466, w_158_000);
  not1 I213_479(w_213_479, w_173_013);
  nand2 I213_513(w_213_513, w_053_106, w_088_119);
  or2  I213_541(w_213_541, w_083_021, w_045_321);
  nand2 I213_577(w_213_577, w_024_534, w_031_457);
  nand2 I213_600(w_213_600, w_211_051, w_065_250);
  or2  I213_605(w_213_605, w_107_252, w_109_331);
  and2 I213_665(w_213_665, w_014_124, w_075_043);
  and2 I214_010(w_214_010, w_001_009, w_017_344);
  and2 I214_016(w_214_016, w_041_535, w_179_184);
  or2  I214_021(w_214_021, w_211_006, w_197_146);
  not1 I214_055(w_214_055, w_138_120);
  nand2 I214_148(w_214_148, w_130_046, w_046_463);
  and2 I214_166(w_214_166, w_053_044, w_117_053);
  nand2 I214_175(w_214_175, w_002_625, w_207_263);
  and2 I214_181(w_214_181, w_105_163, w_057_094);
  or2  I214_201(w_214_201, w_141_008, w_099_113);
  or2  I214_203(w_214_203, w_080_176, w_202_292);
  or2  I214_206(w_214_206, w_100_022, w_123_471);
  not1 I214_225(w_214_225, w_022_117);
  and2 I214_280(w_214_280, w_079_033, w_171_425);
  and2 I214_371(w_214_371, w_209_043, w_191_047);
  or2  I214_381(w_214_381, w_196_212, w_134_076);
  or2  I214_448(w_214_448, w_084_029, w_017_214);
  not1 I214_457(w_214_457, w_192_010);
  not1 I214_518(w_214_518, w_020_051);
  nand2 I214_550(w_214_550, w_143_066, w_153_047);
  or2  I214_577(w_214_577, w_085_299, w_171_731);
  not1 I214_593(w_214_595, w_214_594);
  or2  I214_594(w_214_596, w_214_616, w_214_595);
  not1 I214_595(w_214_597, w_214_596);
  not1 I214_596(w_214_598, w_214_597);
  nand2 I214_597(w_214_599, w_202_022, w_214_598);
  and2 I214_598(w_214_600, w_003_075, w_214_599);
  not1 I214_599(w_214_594, w_214_600);
  not1 I214_600(w_214_605, w_214_604);
  or2  I214_601(w_214_606, w_127_004, w_214_605);
  or2  I214_602(w_214_607, w_214_606, w_149_138);
  and2 I214_603(w_214_608, w_214_607, w_038_538);
  not1 I214_604(w_214_609, w_214_608);
  and2 I214_605(w_214_610, w_214_609, w_086_343);
  not1 I214_606(w_214_611, w_214_610);
  not1 I214_607(w_214_612, w_214_611);
  and2 I214_608(w_214_613, w_214_612, w_106_089);
  and2 I214_609(w_214_614, w_155_289, w_214_613);
  not1 I214_610(w_214_604, w_214_596);
  and2 I214_611(w_214_616, w_208_238, w_214_614);
  nand2 I215_015(w_215_015, w_213_665, w_095_023);
  nand2 I215_024(w_215_024, w_134_218, w_201_035);
  or2  I215_025(w_215_025, w_079_021, w_018_010);
  not1 I215_038(w_215_038, w_187_011);
  nand2 I215_049(w_215_049, w_199_156, w_097_553);
  or2  I215_099(w_215_099, w_140_216, w_133_373);
  not1 I215_106(w_215_106, w_203_045);
  not1 I215_124(w_215_124, w_067_134);
  or2  I215_138(w_215_138, w_052_012, w_090_535);
  and2 I215_139(w_215_139, w_122_041, w_133_290);
  not1 I215_166(w_215_166, w_160_148);
  not1 I215_197(w_215_197, w_084_011);
  and2 I215_203(w_215_203, w_080_360, w_012_106);
  and2 I215_206(w_215_206, w_070_437, w_047_341);
  or2  I215_211(w_215_211, w_082_247, w_128_191);
  not1 I215_246(w_215_246, w_185_185);
  not1 I215_249(w_215_249, w_196_111);
  not1 I215_286(w_215_286, w_032_307);
  not1 I215_335(w_215_335, w_172_012);
  not1 I215_344(w_215_344, w_040_616);
  nand2 I215_346(w_215_346, w_066_558, w_063_026);
  not1 I215_429(w_215_429, w_104_033);
  or2  I215_434(w_215_434, w_026_459, w_028_390);
  not1 I215_438(w_215_438, w_045_017);
  or2  I215_487(w_215_487, w_165_049, w_169_187);
  and2 I215_494(w_215_494, w_200_216, w_147_116);
  not1 I215_532(w_215_532, w_161_074);
  and2 I215_533(w_215_533, w_136_005, w_010_151);
  nand2 I216_002(w_216_002, w_056_049, w_159_039);
  nand2 I216_034(w_216_034, w_082_540, w_003_014);
  nand2 I216_044(w_216_044, w_213_086, w_136_047);
  and2 I216_048(w_216_048, w_053_017, w_099_148);
  nand2 I216_088(w_216_088, w_036_255, w_179_767);
  not1 I216_105(w_216_105, w_048_004);
  nand2 I216_149(w_216_149, w_157_051, w_111_062);
  nand2 I216_169(w_216_169, w_139_004, w_070_155);
  nand2 I216_203(w_216_203, w_191_210, w_032_502);
  and2 I216_234(w_216_234, w_106_170, w_177_160);
  nand2 I216_236(w_216_236, w_060_366, w_129_087);
  nand2 I216_253(w_216_253, w_071_095, w_081_014);
  not1 I216_262(w_216_262, w_082_291);
  nand2 I216_281(w_216_281, w_078_329, w_206_009);
  nand2 I216_290(w_216_290, w_096_003, w_166_287);
  and2 I216_301(w_216_301, w_001_012, w_100_061);
  not1 I216_308(w_216_308, w_132_152);
  not1 I216_340(w_216_340, w_027_096);
  not1 I216_345(w_216_345, w_094_120);
  and2 I216_352(w_216_352, w_082_070, w_030_235);
  or2  I216_357(w_216_357, w_197_228, w_081_015);
  nand2 I216_362(w_216_362, w_035_030, w_002_621);
  or2  I216_376(w_216_376, w_153_018, w_021_016);
  or2  I216_377(w_216_377, w_023_205, w_141_079);
  nand2 I216_410(w_216_410, w_123_112, w_205_245);
  not1 I217_001(w_217_001, w_017_091);
  and2 I217_006(w_217_006, w_209_342, w_133_000);
  nand2 I217_008(w_217_008, w_115_209, w_131_480);
  nand2 I217_014(w_217_014, w_066_141, w_215_532);
  or2  I217_018(w_217_018, w_033_475, w_161_065);
  not1 I217_020(w_217_020, w_059_218);
  and2 I217_023(w_217_023, w_111_027, w_020_163);
  or2  I217_031(w_217_031, w_180_011, w_032_508);
  and2 I217_034(w_217_034, w_150_296, w_135_194);
  nand2 I217_049(w_217_049, w_066_433, w_105_052);
  and2 I217_051(w_217_051, w_136_060, w_205_285);
  or2  I217_054(w_217_054, w_000_527, w_001_007);
  not1 I217_060(w_217_060, w_137_176);
  nand2 I217_061(w_217_061, w_135_086, w_081_011);
  not1 I217_064(w_217_064, w_179_141);
  or2  I217_068(w_217_068, w_100_063, w_215_211);
  and2 I217_074(w_217_074, w_013_415, w_162_003);
  or2  I217_078(w_217_078, w_167_022, w_137_443);
  nand2 I217_083(w_217_083, w_114_069, w_172_003);
  not1 I218_080(w_218_080, w_048_014);
  nand2 I218_124(w_218_124, w_149_590, w_207_198);
  and2 I218_178(w_218_178, w_124_291, w_040_358);
  and2 I218_180(w_218_180, w_144_045, w_097_205);
  nand2 I218_189(w_218_189, w_106_000, w_040_278);
  or2  I218_195(w_218_195, w_035_092, w_153_053);
  and2 I218_261(w_218_261, w_074_334, w_146_275);
  not1 I218_334(w_218_334, w_104_284);
  not1 I218_338(w_218_338, w_137_099);
  and2 I218_380(w_218_380, w_207_110, w_177_333);
  and2 I218_576(w_218_576, w_158_001, w_075_133);
  nand2 I218_584(w_218_584, w_200_359, w_061_270);
  nand2 I218_595(w_218_595, w_110_260, w_212_092);
  or2  I218_599(w_218_599, w_114_181, w_102_424);
  and2 I218_660(w_218_660, w_015_079, w_047_018);
  or2  I218_671(w_218_671, w_080_098, w_104_000);
  not1 I218_698(w_218_698, w_038_590);
  nand2 I218_701(w_218_701, w_093_180, w_151_156);
  or2  I218_725(w_218_725, w_201_226, w_037_277);
  or2  I218_775(w_218_777, w_128_426, w_218_776);
  and2 I218_776(w_218_778, w_185_202, w_218_777);
  not1 I218_777(w_218_779, w_218_778);
  or2  I218_778(w_218_780, w_218_779, w_013_443);
  and2 I218_779(w_218_781, w_218_780, w_055_220);
  and2 I218_780(w_218_782, w_183_139, w_218_781);
  and2 I218_781(w_218_783, w_218_782, w_218_802);
  and2 I218_782(w_218_784, w_218_783, w_130_088);
  and2 I218_783(w_218_785, w_218_784, w_141_000);
  or2  I218_784(w_218_776, w_218_785, w_161_607);
  not1 I218_785(w_218_790, w_218_789);
  and2 I218_786(w_218_791, w_218_790, w_013_184);
  nand2 I218_787(w_218_792, w_218_791, w_216_377);
  not1 I218_788(w_218_793, w_218_792);
  not1 I218_789(w_218_794, w_218_793);
  nand2 I218_790(w_218_795, w_021_014, w_218_794);
  nand2 I218_791(w_218_796, w_171_334, w_218_795);
  or2  I218_792(w_218_797, w_005_173, w_218_796);
  or2  I218_793(w_218_798, w_072_102, w_218_797);
  or2  I218_794(w_218_799, w_193_091, w_218_798);
  and2 I218_795(w_218_800, w_218_799, w_138_304);
  not1 I218_796(w_218_789, w_218_783);
  and2 I218_797(w_218_802, w_041_692, w_218_800);
  and2 I219_005(w_219_005, w_131_149, w_103_289);
  and2 I219_008(w_219_008, w_096_005, w_134_073);
  and2 I219_067(w_219_067, w_182_026, w_050_333);
  and2 I219_090(w_219_090, w_034_031, w_204_043);
  or2  I219_242(w_219_242, w_024_045, w_185_109);
  nand2 I219_244(w_219_244, w_089_098, w_052_001);
  not1 I219_265(w_219_265, w_145_046);
  nand2 I219_340(w_219_340, w_185_137, w_186_208);
  not1 I219_413(w_219_413, w_058_536);
  nand2 I219_439(w_219_439, w_089_206, w_139_009);
  and2 I219_522(w_219_522, w_095_054, w_090_036);
  nand2 I219_604(w_219_604, w_063_149, w_037_146);
  and2 I219_626(w_219_626, w_065_246, w_182_025);
  nand2 I219_636(w_219_636, w_177_025, w_080_029);
  nand2 I219_644(w_219_644, w_118_031, w_058_216);
  not1 I219_656(w_219_656, w_007_113);
  or2  I219_668(w_219_668, w_032_541, w_051_250);
  not1 I219_738(w_219_738, w_069_242);
  or2  I220_119(w_220_119, w_145_002, w_153_049);
  or2  I220_142(w_220_142, w_103_287, w_062_352);
  or2  I220_186(w_220_186, w_190_041, w_105_351);
  nand2 I220_195(w_220_195, w_092_484, w_218_380);
  not1 I220_197(w_220_197, w_202_029);
  and2 I220_231(w_220_231, w_128_067, w_138_056);
  not1 I220_248(w_220_248, w_001_024);
  not1 I220_263(w_220_263, w_205_035);
  nand2 I220_265(w_220_265, w_030_052, w_182_002);
  and2 I220_290(w_220_290, w_088_005, w_089_086);
  and2 I220_322(w_220_322, w_132_393, w_177_238);
  nand2 I220_337(w_220_337, w_166_145, w_200_211);
  or2  I220_340(w_220_340, w_202_116, w_156_232);
  not1 I220_346(w_220_346, w_139_010);
  not1 I220_350(w_220_350, w_100_092);
  nand2 I220_367(w_220_367, w_065_453, w_059_589);
  nand2 I220_371(w_220_371, w_147_175, w_182_023);
  or2  I220_377(w_220_377, w_201_203, w_140_202);
  and2 I220_380(w_220_380, w_076_479, w_146_273);
  or2  I221_018(w_221_018, w_183_193, w_106_124);
  not1 I221_033(w_221_033, w_127_047);
  not1 I221_044(w_221_044, w_031_001);
  or2  I221_054(w_221_054, w_003_031, w_152_002);
  or2  I221_063(w_221_063, w_044_540, w_149_018);
  not1 I221_067(w_221_067, w_117_024);
  nand2 I221_069(w_221_069, w_066_246, w_161_369);
  not1 I221_071(w_221_071, w_088_093);
  not1 I221_125(w_221_125, w_062_401);
  not1 I221_143(w_221_143, w_156_296);
  nand2 I221_159(w_221_159, w_053_046, w_089_142);
  or2  I221_175(w_221_175, w_073_183, w_057_160);
  or2  I221_190(w_221_190, w_033_583, w_088_043);
  not1 I221_207(w_221_207, w_197_152);
  and2 I221_213(w_221_213, w_094_009, w_153_085);
  nand2 I221_225(w_221_225, w_180_019, w_201_009);
  nand2 I222_026(w_222_026, w_017_134, w_159_083);
  not1 I222_032(w_222_032, w_130_469);
  and2 I222_120(w_222_120, w_115_055, w_120_345);
  nand2 I222_141(w_222_141, w_019_005, w_211_019);
  or2  I222_163(w_222_163, w_141_000, w_216_034);
  or2  I222_185(w_222_185, w_131_054, w_201_280);
  or2  I222_226(w_222_226, w_201_026, w_035_056);
  nand2 I222_236(w_222_236, w_133_249, w_169_305);
  and2 I222_255(w_222_255, w_006_154, w_205_537);
  or2  I222_315(w_222_315, w_096_001, w_026_231);
  not1 I222_321(w_222_321, w_178_077);
  and2 I222_422(w_222_422, w_147_160, w_085_272);
  not1 I222_469(w_222_469, w_084_010);
  or2  I222_521(w_222_521, w_172_044, w_160_433);
  nand2 I222_623(w_222_623, w_213_513, w_100_071);
  and2 I222_628(w_222_628, w_000_097, w_073_602);
  nand2 I223_016(w_223_016, w_174_029, w_006_171);
  and2 I223_027(w_223_027, w_149_438, w_066_115);
  and2 I223_040(w_223_040, w_074_108, w_167_040);
  nand2 I223_047(w_223_047, w_010_553, w_058_515);
  nand2 I223_073(w_223_073, w_195_107, w_054_252);
  and2 I223_075(w_223_075, w_145_027, w_057_271);
  not1 I223_079(w_223_079, w_127_026);
  or2  I223_140(w_223_140, w_134_071, w_168_088);
  not1 I223_141(w_223_141, w_104_311);
  not1 I223_145(w_223_145, w_104_029);
  not1 I223_146(w_223_146, w_069_174);
  not1 I223_151(w_223_151, w_197_161);
  or2  I223_156(w_223_156, w_121_027, w_108_002);
  nand2 I223_166(w_223_166, w_004_279, w_064_150);
  nand2 I223_184(w_223_184, w_038_321, w_127_017);
  nand2 I223_201(w_223_201, w_055_219, w_168_110);
  nand2 I223_202(w_223_202, w_164_277, w_071_094);
  or2  I223_209(w_223_209, w_009_507, w_165_095);
  or2  I223_218(w_223_218, w_103_143, w_152_045);
  or2  I223_235(w_223_235, w_104_004, w_008_683);
  nand2 I223_241(w_223_241, w_028_392, w_213_007);
  and2 I223_267(w_223_267, w_136_044, w_187_001);
  nand2 I223_284(w_223_284, w_134_017, w_134_396);
  not1 I224_024(w_224_024, w_009_264);
  not1 I224_036(w_224_036, w_166_103);
  nand2 I224_049(w_224_049, w_168_542, w_149_179);
  not1 I224_069(w_224_069, w_120_241);
  or2  I224_083(w_224_083, w_156_224, w_177_307);
  or2  I224_095(w_224_095, w_179_164, w_140_188);
  not1 I224_104(w_224_104, w_152_198);
  nand2 I224_113(w_224_113, w_030_372, w_220_367);
  nand2 I224_114(w_224_114, w_141_139, w_147_022);
  and2 I224_156(w_224_156, w_129_067, w_092_070);
  and2 I224_178(w_224_178, w_112_121, w_028_142);
  and2 I224_210(w_224_210, w_187_014, w_015_637);
  and2 I224_241(w_224_241, w_106_065, w_130_511);
  and2 I224_256(w_224_256, w_084_002, w_162_004);
  not1 I224_303(w_224_303, w_124_061);
  not1 I224_331(w_224_331, w_073_095);
  nand2 I224_353(w_224_353, w_083_193, w_186_450);
  or2  I224_386(w_224_386, w_085_029, w_124_286);
  nand2 I224_401(w_224_401, w_169_279, w_046_583);
  not1 I224_405(w_224_405, w_163_163);
  and2 I224_421(w_224_421, w_215_025, w_061_182);
  not1 I224_494(w_224_494, w_110_147);
  or2  I224_524(w_224_524, w_149_600, w_100_115);
  nand2 I225_010(w_225_010, w_017_197, w_150_361);
  not1 I225_019(w_225_019, w_118_094);
  nand2 I225_033(w_225_033, w_081_013, w_045_362);
  nand2 I225_051(w_225_051, w_056_597, w_100_092);
  not1 I225_053(w_225_053, w_152_089);
  nand2 I225_059(w_225_059, w_220_263, w_173_015);
  or2  I225_062(w_225_062, w_209_087, w_115_037);
  and2 I225_086(w_225_086, w_002_301, w_051_279);
  and2 I225_102(w_225_102, w_150_159, w_217_083);
  not1 I225_104(w_225_104, w_191_163);
  or2  I225_112(w_225_112, w_166_127, w_104_057);
  not1 I225_142(w_225_142, w_059_309);
  not1 I225_154(w_225_154, w_095_030);
  and2 I225_168(w_225_168, w_144_302, w_210_003);
  nand2 I225_180(w_225_180, w_007_421, w_219_340);
  and2 I225_194(w_225_194, w_164_339, w_044_175);
  nand2 I225_204(w_225_204, w_091_133, w_031_130);
  or2  I225_220(w_225_220, w_217_064, w_224_210);
  not1 I225_227(w_225_227, w_175_422);
  and2 I225_240(w_225_240, w_117_016, w_057_086);
  and2 I226_019(w_226_019, w_217_060, w_206_119);
  nand2 I226_077(w_226_077, w_083_007, w_160_382);
  nand2 I226_092(w_226_092, w_174_072, w_019_006);
  or2  I226_138(w_226_138, w_182_021, w_061_302);
  and2 I226_152(w_226_152, w_041_110, w_051_381);
  not1 I226_171(w_226_171, w_051_031);
  and2 I226_189(w_226_189, w_054_214, w_183_183);
  or2  I226_190(w_226_190, w_029_082, w_172_030);
  or2  I226_199(w_226_199, w_136_051, w_177_385);
  and2 I226_219(w_226_219, w_107_183, w_113_081);
  and2 I226_222(w_226_222, w_024_195, w_031_509);
  and2 I226_310(w_226_310, w_174_107, w_127_054);
  and2 I226_393(w_226_393, w_126_078, w_113_114);
  nand2 I226_401(w_226_401, w_111_023, w_017_451);
  not1 I226_455(w_226_455, w_010_592);
  and2 I226_475(w_226_475, w_156_007, w_177_166);
  not1 I226_497(w_226_497, w_053_108);
  and2 I226_556(w_226_558, w_026_226, w_226_557);
  and2 I226_557(w_226_559, w_226_558, w_063_341);
  not1 I226_558(w_226_557, w_226_559);
  not1 I227_026(w_227_026, w_212_204);
  or2  I227_036(w_227_036, w_188_007, w_063_262);
  not1 I227_062(w_227_062, w_033_753);
  and2 I227_160(w_227_160, w_093_200, w_029_015);
  not1 I227_163(w_227_163, w_060_161);
  nand2 I227_173(w_227_173, w_128_174, w_081_004);
  not1 I227_209(w_227_209, w_119_162);
  and2 I227_231(w_227_231, w_121_039, w_066_181);
  not1 I227_269(w_227_269, w_098_038);
  nand2 I227_278(w_227_278, w_215_197, w_054_344);
  nand2 I227_339(w_227_339, w_117_014, w_132_260);
  nand2 I227_403(w_227_403, w_049_161, w_168_452);
  not1 I227_475(w_227_475, w_148_536);
  and2 I227_485(w_227_485, w_162_023, w_116_497);
  and2 I227_513(w_227_513, w_099_188, w_050_479);
  nand2 I227_584(w_227_584, w_081_011, w_040_132);
  and2 I227_597(w_227_597, w_098_009, w_153_038);
  and2 I227_612(w_227_612, w_072_092, w_220_263);
  not1 I227_620(w_227_620, w_195_205);
  nand2 I227_647(w_227_647, w_010_226, w_154_093);
  nand2 I227_658(w_227_658, w_011_052, w_110_075);
  and2 I228_005(w_228_005, w_011_317, w_072_113);
  not1 I228_011(w_228_011, w_102_619);
  nand2 I228_013(w_228_013, w_025_202, w_060_020);
  not1 I228_039(w_228_039, w_192_145);
  nand2 I228_050(w_228_050, w_056_038, w_043_030);
  and2 I228_066(w_228_066, w_019_013, w_227_620);
  nand2 I228_105(w_228_105, w_004_041, w_042_367);
  nand2 I228_123(w_228_123, w_141_059, w_024_413);
  not1 I228_146(w_228_146, w_201_007);
  not1 I228_214(w_228_214, w_082_576);
  and2 I228_343(w_228_343, w_187_010, w_192_082);
  and2 I228_374(w_228_374, w_052_034, w_146_182);
  and2 I228_466(w_228_466, w_044_139, w_127_053);
  nand2 I228_533(w_228_533, w_225_227, w_014_055);
  and2 I228_578(w_228_578, w_203_074, w_178_107);
  or2  I228_580(w_228_580, w_015_314, w_215_429);
  not1 I228_584(w_228_584, w_031_122);
  and2 I228_588(w_228_588, w_068_309, w_160_793);
  nand2 I228_625(w_228_625, w_096_001, w_216_044);
  nand2 I228_627(w_228_627, w_129_372, w_186_336);
  or2  I229_000(w_229_000, w_226_189, w_173_003);
  nand2 I229_003(w_229_003, w_001_003, w_155_148);
  or2  I229_015(w_229_015, w_221_054, w_217_078);
  or2  I229_034(w_229_034, w_110_242, w_199_073);
  not1 I229_035(w_229_035, w_171_119);
  nand2 I229_041(w_229_041, w_117_048, w_140_009);
  nand2 I229_046(w_229_046, w_023_129, w_213_339);
  not1 I229_086(w_229_086, w_021_074);
  nand2 I229_136(w_229_136, w_192_079, w_055_110);
  and2 I229_192(w_229_192, w_208_400, w_146_324);
  or2  I229_247(w_229_247, w_171_470, w_218_124);
  and2 I229_268(w_229_268, w_059_286, w_051_279);
  not1 I229_285(w_229_285, w_045_177);
  not1 I229_323(w_229_323, w_140_189);
  not1 I229_455(w_229_455, w_198_078);
  or2  I230_007(w_230_007, w_077_479, w_091_166);
  and2 I230_010(w_230_010, w_129_135, w_017_589);
  and2 I230_024(w_230_024, w_221_063, w_099_274);
  not1 I230_027(w_230_027, w_128_345);
  or2  I230_037(w_230_037, w_059_167, w_185_108);
  and2 I230_038(w_230_038, w_202_079, w_046_234);
  or2  I230_055(w_230_055, w_092_551, w_200_183);
  or2  I230_060(w_230_060, w_038_043, w_223_146);
  or2  I230_077(w_230_077, w_198_054, w_046_599);
  or2  I230_080(w_230_080, w_005_009, w_071_085);
  or2  I230_095(w_230_095, w_051_170, w_035_090);
  not1 I230_157(w_230_157, w_057_007);
  nand2 I230_197(w_230_197, w_213_368, w_000_528);
  nand2 I230_215(w_230_215, w_109_213, w_165_079);
  not1 I230_233(w_230_233, w_069_076);
  nand2 I230_266(w_230_266, w_225_019, w_114_198);
  and2 I230_298(w_230_298, w_116_365, w_163_065);
  or2  I230_320(w_230_322, w_230_321, w_155_149);
  or2  I230_321(w_230_323, w_181_208, w_230_322);
  or2  I230_322(w_230_324, w_090_052, w_230_323);
  and2 I230_323(w_230_325, w_004_090, w_230_324);
  nand2 I230_324(w_230_326, w_230_325, w_226_497);
  nand2 I230_325(w_230_327, w_230_326, w_230_344);
  not1 I230_326(w_230_328, w_230_327);
  and2 I230_327(w_230_329, w_230_328, w_009_560);
  nand2 I230_328(w_230_321, w_191_065, w_230_329);
  nand2 I230_329(w_230_334, w_230_333, w_151_080);
  nand2 I230_330(w_230_335, w_134_151, w_230_334);
  or2  I230_331(w_230_336, w_143_374, w_230_335);
  nand2 I230_332(w_230_337, w_046_450, w_230_336);
  not1 I230_333(w_230_338, w_230_337);
  or2  I230_334(w_230_339, w_230_338, w_081_019);
  and2 I230_335(w_230_340, w_212_073, w_230_339);
  nand2 I230_336(w_230_341, w_230_340, w_133_081);
  and2 I230_337(w_230_342, w_230_341, w_082_196);
  not1 I230_338(w_230_333, w_230_327);
  and2 I230_339(w_230_344, w_163_515, w_230_342);
  and2 I231_001(w_231_001, w_023_041, w_216_236);
  nand2 I231_003(w_231_003, w_023_065, w_138_051);
  or2  I231_009(w_231_009, w_018_022, w_201_193);
  not1 I231_056(w_231_056, w_042_385);
  and2 I231_064(w_231_064, w_218_584, w_146_085);
  nand2 I231_157(w_231_157, w_075_033, w_230_197);
  and2 I231_160(w_231_160, w_073_592, w_046_599);
  and2 I231_198(w_231_198, w_073_284, w_017_056);
  not1 I231_199(w_231_199, w_224_353);
  nand2 I231_220(w_231_220, w_165_088, w_011_374);
  nand2 I231_321(w_231_321, w_187_013, w_094_469);
  or2  I231_322(w_231_322, w_164_424, w_104_062);
  nand2 I231_427(w_231_427, w_096_003, w_221_175);
  and2 I231_463(w_231_463, w_158_003, w_028_245);
  or2  I231_464(w_231_464, w_101_156, w_033_775);
  and2 I231_530(w_231_530, w_045_063, w_180_019);
  nand2 I231_532(w_231_532, w_030_183, w_219_090);
  not1 I231_537(w_231_537, w_223_075);
  and2 I231_545(w_231_545, w_196_079, w_150_000);
  nand2 I231_579(w_231_579, w_035_083, w_196_101);
  or2  I232_035(w_232_035, w_131_087, w_069_153);
  not1 I232_050(w_232_050, w_171_135);
  nand2 I232_069(w_232_069, w_092_377, w_001_006);
  nand2 I232_077(w_232_077, w_161_567, w_200_178);
  not1 I232_079(w_232_079, w_094_373);
  or2  I232_084(w_232_084, w_175_285, w_121_054);
  nand2 I232_103(w_232_103, w_020_092, w_186_235);
  and2 I232_125(w_232_125, w_082_112, w_148_010);
  and2 I232_150(w_232_150, w_190_040, w_225_112);
  not1 I232_166(w_232_166, w_134_163);
  and2 I232_172(w_232_172, w_075_079, w_057_171);
  not1 I232_190(w_232_190, w_022_167);
  not1 I232_237(w_232_237, w_088_032);
  nand2 I232_295(w_232_295, w_136_063, w_208_161);
  nand2 I232_318(w_232_318, w_053_004, w_040_098);
  not1 I232_332(w_232_332, w_096_005);
  or2  I232_376(w_232_376, w_023_170, w_182_024);
  nand2 I232_381(w_232_381, w_035_085, w_043_026);
  and2 I232_399(w_232_399, w_099_058, w_140_015);
  not1 I232_456(w_232_456, w_179_140);
  not1 I232_457(w_232_457, w_133_235);
  or2  I232_478(w_232_478, w_085_080, w_129_175);
  or2  I232_479(w_232_479, w_144_406, w_055_106);
  nand2 I232_503(w_232_503, w_222_321, w_096_005);
  and2 I232_507(w_232_509, w_232_508, w_232_529);
  and2 I232_508(w_232_510, w_232_509, w_052_011);
  and2 I232_509(w_232_511, w_232_510, w_092_516);
  nand2 I232_510(w_232_512, w_012_039, w_232_511);
  and2 I232_511(w_232_513, w_230_010, w_232_512);
  not1 I232_512(w_232_508, w_232_513);
  nand2 I232_513(w_232_518, w_053_083, w_232_517);
  not1 I232_514(w_232_519, w_232_518);
  nand2 I232_515(w_232_520, w_232_519, w_126_058);
  not1 I232_516(w_232_521, w_232_520);
  or2  I232_517(w_232_522, w_232_521, w_038_340);
  not1 I232_518(w_232_523, w_232_522);
  nand2 I232_519(w_232_524, w_227_513, w_232_523);
  nand2 I232_520(w_232_525, w_173_018, w_232_524);
  nand2 I232_521(w_232_526, w_148_576, w_232_525);
  and2 I232_522(w_232_527, w_024_300, w_232_526);
  not1 I232_523(w_232_517, w_232_509);
  and2 I232_524(w_232_529, w_179_039, w_232_527);
  nand2 I233_001(w_233_001, w_010_373, w_094_610);
  nand2 I233_012(w_233_012, w_107_047, w_100_080);
  and2 I233_037(w_233_037, w_136_032, w_114_003);
  and2 I233_038(w_233_038, w_144_473, w_017_008);
  and2 I233_068(w_233_068, w_120_506, w_007_155);
  and2 I233_088(w_233_088, w_197_312, w_221_143);
  nand2 I233_101(w_233_101, w_194_178, w_201_027);
  nand2 I233_168(w_233_168, w_073_117, w_042_095);
  and2 I233_169(w_233_169, w_093_133, w_088_028);
  nand2 I233_171(w_233_171, w_174_110, w_206_139);
  or2  I233_204(w_233_204, w_073_379, w_131_308);
  nand2 I233_234(w_233_234, w_113_289, w_153_060);
  not1 I233_239(w_233_239, w_107_100);
  nand2 I233_249(w_233_249, w_206_058, w_063_374);
  or2  I233_326(w_233_326, w_193_080, w_174_044);
  nand2 I233_353(w_233_353, w_025_194, w_105_372);
  and2 I233_378(w_233_378, w_226_393, w_046_238);
  not1 I233_386(w_233_386, w_121_050);
  not1 I234_038(w_234_038, w_045_388);
  or2  I234_086(w_234_086, w_114_138, w_158_001);
  not1 I234_111(w_234_111, w_192_019);
  or2  I234_145(w_234_145, w_008_595, w_151_200);
  not1 I234_147(w_234_147, w_226_199);
  nand2 I234_153(w_234_153, w_126_115, w_193_151);
  and2 I234_159(w_234_159, w_081_014, w_070_365);
  nand2 I234_182(w_234_182, w_097_012, w_184_032);
  nand2 I234_195(w_234_195, w_046_351, w_160_237);
  or2  I234_254(w_234_254, w_172_052, w_011_419);
  and2 I234_309(w_234_309, w_035_049, w_130_377);
  or2  I234_326(w_234_326, w_007_043, w_171_252);
  nand2 I234_403(w_234_403, w_157_036, w_062_465);
  or2  I234_429(w_234_429, w_034_007, w_178_049);
  not1 I235_018(w_235_018, w_023_111);
  not1 I235_034(w_235_034, w_070_121);
  and2 I235_046(w_235_046, w_068_052, w_147_063);
  or2  I235_056(w_235_056, w_171_722, w_210_044);
  not1 I235_062(w_235_062, w_203_027);
  nand2 I235_066(w_235_066, w_105_079, w_186_084);
  not1 I235_070(w_235_070, w_067_076);
  not1 I235_079(w_235_079, w_052_041);
  or2  I235_083(w_235_083, w_207_378, w_044_303);
  and2 I235_101(w_235_101, w_008_028, w_196_196);
  not1 I235_112(w_235_112, w_192_176);
  nand2 I235_114(w_235_114, w_037_287, w_028_260);
  or2  I235_115(w_235_115, w_149_081, w_207_546);
  or2  I235_121(w_235_121, w_108_067, w_206_144);
  or2  I235_141(w_235_141, w_045_131, w_124_252);
  or2  I235_177(w_235_177, w_170_085, w_055_076);
  or2  I235_181(w_235_181, w_149_207, w_099_019);
  or2  I235_206(w_235_206, w_027_119, w_068_041);
  and2 I236_010(w_236_010, w_224_024, w_144_125);
  nand2 I236_028(w_236_028, w_034_035, w_060_033);
  and2 I236_046(w_236_046, w_080_185, w_175_504);
  and2 I236_097(w_236_097, w_035_037, w_159_018);
  nand2 I236_132(w_236_132, w_153_029, w_138_051);
  not1 I236_159(w_236_159, w_203_090);
  nand2 I236_166(w_236_166, w_191_215, w_129_041);
  or2  I236_199(w_236_199, w_131_048, w_177_280);
  or2  I237_000(w_237_000, w_174_028, w_132_313);
  not1 I237_012(w_237_012, w_164_085);
  nand2 I237_033(w_237_033, w_113_341, w_105_267);
  not1 I237_062(w_237_062, w_084_028);
  or2  I237_063(w_237_063, w_187_016, w_200_440);
  or2  I237_074(w_237_074, w_206_082, w_148_123);
  not1 I237_081(w_237_081, w_206_038);
  or2  I237_084(w_237_084, w_034_046, w_216_281);
  nand2 I237_107(w_237_107, w_145_030, w_186_257);
  nand2 I237_111(w_237_111, w_057_123, w_205_519);
  or2  I237_128(w_237_128, w_095_042, w_181_142);
  nand2 I237_130(w_237_130, w_030_252, w_016_007);
  not1 I237_131(w_237_131, w_211_034);
  or2  I237_134(w_237_134, w_036_154, w_228_627);
  or2  I238_000(w_238_000, w_011_309, w_170_222);
  nand2 I238_010(w_238_010, w_169_236, w_114_114);
  and2 I238_021(w_238_021, w_115_178, w_231_464);
  and2 I238_052(w_238_052, w_159_030, w_159_108);
  and2 I238_105(w_238_105, w_189_443, w_184_019);
  and2 I238_120(w_238_120, w_148_684, w_183_133);
  nand2 I238_141(w_238_141, w_090_222, w_001_007);
  and2 I238_150(w_238_150, w_163_050, w_112_143);
  and2 I238_189(w_238_189, w_078_102, w_099_205);
  or2  I238_195(w_238_195, w_216_345, w_140_062);
  or2  I238_235(w_238_235, w_128_115, w_202_278);
  not1 I238_264(w_238_264, w_036_144);
  nand2 I238_395(w_238_395, w_080_289, w_228_533);
  and2 I238_412(w_238_412, w_015_351, w_147_214);
  not1 I238_429(w_238_429, w_108_021);
  and2 I238_449(w_238_449, w_237_130, w_020_018);
  nand2 I239_000(w_239_000, w_065_666, w_090_564);
  and2 I240_005(w_240_005, w_215_494, w_123_251);
  not1 I240_019(w_240_019, w_203_339);
  nand2 I240_024(w_240_024, w_162_017, w_051_262);
  not1 I240_026(w_240_026, w_038_368);
  not1 I240_038(w_240_038, w_166_109);
  and2 I240_047(w_240_047, w_018_026, w_084_045);
  not1 I240_055(w_240_055, w_045_300);
  not1 I240_056(w_240_056, w_192_189);
  not1 I240_072(w_240_072, w_224_036);
  or2  I240_076(w_240_076, w_154_030, w_173_012);
  nand2 I240_090(w_240_090, w_193_272, w_006_118);
  and2 I240_098(w_240_098, w_058_065, w_069_213);
  and2 I240_101(w_240_101, w_212_064, w_193_097);
  nand2 I240_104(w_240_104, w_041_721, w_022_347);
  and2 I240_109(w_240_109, w_125_308, w_075_078);
  or2  I240_114(w_240_114, w_060_288, w_128_295);
  and2 I240_125(w_240_125, w_018_008, w_126_119);
  nand2 I240_142(w_240_142, w_061_063, w_047_367);
  or2  I240_147(w_240_147, w_144_346, w_115_178);
  nand2 I240_159(w_240_159, w_041_189, w_147_062);
  and2 I240_171(w_240_171, w_200_028, w_108_073);
  or2  I240_184(w_240_184, w_039_066, w_123_097);
  and2 I241_000(w_241_000, w_154_056, w_220_186);
  not1 I241_002(w_241_002, w_235_206);
  or2  I241_008(w_241_008, w_050_626, w_218_195);
  or2  I241_010(w_241_010, w_216_149, w_220_290);
  or2  I241_011(w_241_011, w_240_184, w_093_239);
  and2 I241_021(w_241_021, w_173_025, w_122_000);
  or2  I241_029(w_241_029, w_176_136, w_125_079);
  and2 I241_030(w_241_030, w_006_015, w_069_097);
  nand2 I241_031(w_241_031, w_000_762, w_002_533);
  nand2 I241_032(w_241_032, w_072_131, w_033_670);
  nand2 I241_033(w_241_033, w_071_058, w_043_021);
  nand2 I241_055(w_241_055, w_180_014, w_027_095);
  or2  I241_058(w_241_058, w_000_402, w_017_227);
  or2  I241_059(w_241_059, w_185_198, w_222_120);
  nand2 I241_068(w_241_068, w_017_598, w_064_012);
  or2  I241_081(w_241_081, w_200_117, w_091_137);
  or2  I241_085(w_241_085, w_191_008, w_232_077);
  and2 I242_000(w_242_000, w_133_159, w_190_040);
  nand2 I242_002(w_242_002, w_222_628, w_059_094);
  nand2 I242_006(w_242_006, w_157_133, w_132_398);
  and2 I242_058(w_242_058, w_060_116, w_224_421);
  and2 I242_077(w_242_077, w_049_237, w_007_205);
  and2 I242_082(w_242_082, w_195_128, w_005_077);
  and2 I242_090(w_242_090, w_192_179, w_218_671);
  or2  I242_093(w_242_093, w_155_403, w_130_239);
  nand2 I242_122(w_242_122, w_046_101, w_166_248);
  and2 I242_132(w_242_132, w_109_233, w_074_033);
  not1 I242_133(w_242_133, w_203_473);
  nand2 I242_134(w_242_134, w_069_230, w_206_046);
  and2 I242_153(w_242_153, w_021_271, w_190_000);
  and2 I242_162(w_242_162, w_158_001, w_205_007);
  or2  I242_163(w_242_163, w_230_215, w_162_008);
  not1 I243_015(w_243_015, w_135_286);
  and2 I243_057(w_243_057, w_219_242, w_026_231);
  and2 I243_072(w_243_072, w_129_226, w_121_009);
  or2  I243_109(w_243_109, w_083_151, w_053_156);
  nand2 I243_111(w_243_111, w_046_516, w_122_055);
  not1 I243_143(w_243_143, w_052_036);
  or2  I243_150(w_243_150, w_151_321, w_019_016);
  nand2 I243_160(w_243_160, w_035_081, w_138_058);
  not1 I243_181(w_243_181, w_021_242);
  nand2 I243_268(w_243_268, w_047_419, w_080_362);
  not1 I243_297(w_243_297, w_043_008);
  and2 I244_000(w_244_000, w_169_200, w_045_220);
  or2  I244_026(w_244_026, w_157_002, w_123_139);
  nand2 I244_053(w_244_053, w_158_003, w_002_218);
  nand2 I244_071(w_244_071, w_209_176, w_033_250);
  and2 I244_081(w_244_081, w_104_290, w_051_009);
  nand2 I244_111(w_244_111, w_140_096, w_087_043);
  or2  I244_117(w_244_117, w_129_120, w_180_012);
  or2  I244_136(w_244_136, w_147_032, w_064_072);
  nand2 I244_185(w_244_185, w_076_447, w_126_055);
  nand2 I244_200(w_244_200, w_201_346, w_220_197);
  nand2 I244_205(w_244_205, w_082_309, w_232_457);
  or2  I244_216(w_244_216, w_086_067, w_193_183);
  or2  I244_220(w_244_220, w_239_000, w_011_401);
  and2 I244_229(w_244_229, w_136_054, w_106_067);
  nand2 I244_238(w_244_238, w_114_220, w_034_018);
  or2  I244_244(w_244_244, w_094_296, w_037_221);
  or2  I244_246(w_244_248, w_244_247, w_119_142);
  nand2 I244_247(w_244_249, w_244_248, w_161_461);
  not1 I244_248(w_244_250, w_244_249);
  or2  I244_249(w_244_251, w_135_156, w_244_250);
  and2 I244_250(w_244_252, w_149_619, w_244_251);
  or2  I244_251(w_244_247, w_198_017, w_244_252);
  nand2 I245_035(w_245_035, w_013_178, w_217_008);
  nand2 I245_153(w_245_153, w_092_229, w_135_429);
  or2  I245_155(w_245_155, w_082_106, w_114_148);
  not1 I245_188(w_245_188, w_066_112);
  nand2 I245_262(w_245_262, w_009_219, w_212_003);
  nand2 I245_339(w_245_339, w_150_067, w_128_152);
  and2 I245_347(w_245_347, w_065_259, w_069_080);
  and2 I245_397(w_245_397, w_190_073, w_042_264);
  nand2 I245_398(w_245_398, w_209_106, w_106_066);
  and2 I245_436(w_245_436, w_018_014, w_083_085);
  and2 I245_448(w_245_448, w_076_062, w_167_043);
  or2  I245_465(w_245_465, w_067_305, w_047_006);
  nand2 I245_507(w_245_507, w_228_588, w_151_130);
  nand2 I245_624(w_245_624, w_237_081, w_011_005);
  and2 I245_660(w_245_660, w_092_563, w_194_238);
  and2 I245_696(w_245_696, w_110_273, w_139_018);
  or2  I245_730(w_245_730, w_231_545, w_013_131);
  nand2 I245_735(w_245_735, w_134_138, w_152_153);
  and2 I245_774(w_244_254, w_171_192, w_244_247);
  or2  I246_014(w_246_014, w_045_235, w_071_097);
  not1 I246_074(w_246_074, w_156_238);
  or2  I246_075(w_246_075, w_127_070, w_037_115);
  not1 I246_079(w_246_079, w_002_595);
  and2 I246_092(w_246_092, w_131_472, w_232_069);
  and2 I246_107(w_246_107, w_036_231, w_028_438);
  or2  I246_119(w_246_119, w_131_345, w_047_288);
  not1 I246_124(w_246_124, w_118_000);
  nand2 I246_286(w_246_286, w_074_046, w_172_012);
  or2  I246_289(w_246_289, w_014_169, w_198_053);
  or2  I246_307(w_246_307, w_175_144, w_041_275);
  and2 I246_482(w_246_482, w_024_528, w_178_049);
  or2  I246_485(w_246_485, w_136_049, w_146_001);
  and2 I246_520(w_246_520, w_120_439, w_190_034);
  or2  I246_521(w_246_521, w_056_051, w_119_070);
  not1 I246_573(w_246_573, w_200_188);
  not1 I246_593(w_246_593, w_244_254);
  or2  I246_607(w_246_607, w_223_027, w_080_063);
  nand2 I246_608(w_246_608, w_209_007, w_211_004);
  or2  I247_000(w_247_000, w_036_141, w_106_098);
  not1 I247_021(w_247_021, w_107_181);
  and2 I247_035(w_247_035, w_051_237, w_037_212);
  and2 I247_076(w_247_076, w_232_237, w_208_259);
  and2 I247_079(w_247_079, w_198_060, w_202_066);
  nand2 I247_107(w_247_107, w_042_199, w_187_026);
  and2 I247_131(w_247_131, w_236_132, w_002_321);
  nand2 I247_135(w_247_135, w_158_004, w_150_253);
  or2  I247_140(w_247_140, w_085_087, w_002_210);
  not1 I247_142(w_247_142, w_085_096);
  not1 I247_147(w_247_147, w_228_580);
  and2 I247_154(w_247_154, w_230_007, w_041_614);
  and2 I247_159(w_247_159, w_195_228, w_232_050);
  nand2 I247_161(w_247_161, w_035_045, w_186_322);
  nand2 I247_162(w_247_162, w_078_560, w_062_268);
  or2  I247_163(w_247_163, w_173_031, w_159_098);
  nand2 I247_170(w_247_170, w_023_019, w_123_096);
  nand2 I247_181(w_247_181, w_078_465, w_186_177);
  or2  I247_183(w_247_183, w_180_003, w_121_129);
  and2 I247_184(w_247_184, w_089_221, w_129_205);
  not1 I248_025(w_248_025, w_195_054);
  nand2 I248_028(w_248_028, w_194_325, w_107_161);
  and2 I248_034(w_248_034, w_061_407, w_247_140);
  and2 I248_039(w_248_039, w_123_153, w_163_284);
  nand2 I248_042(w_248_042, w_041_300, w_198_060);
  nand2 I248_045(w_248_045, w_056_238, w_233_171);
  and2 I248_063(w_248_063, w_208_273, w_190_005);
  or2  I248_087(w_248_087, w_051_342, w_144_182);
  or2  I248_099(w_248_099, w_172_044, w_119_146);
  nand2 I248_111(w_248_111, w_153_022, w_080_290);
  or2  I248_130(w_248_130, w_047_255, w_124_078);
  not1 I248_136(w_248_136, w_192_165);
  and2 I248_142(w_248_142, w_209_139, w_006_074);
  not1 I249_069(w_249_069, w_067_373);
  or2  I249_150(w_249_150, w_169_344, w_068_138);
  and2 I249_152(w_249_152, w_248_045, w_185_059);
  or2  I249_169(w_249_169, w_192_172, w_248_087);
  nand2 I249_187(w_249_187, w_146_256, w_129_245);
  nand2 I249_191(w_249_191, w_209_054, w_226_455);
  not1 I249_202(w_249_202, w_225_102);
  and2 I249_268(w_249_268, w_020_028, w_140_024);
  nand2 I249_280(w_249_280, w_172_042, w_150_324);
  not1 I249_333(w_249_333, w_013_458);
  or2  I249_340(w_249_340, w_064_093, w_219_604);
  and2 I250_012(w_250_012, w_071_151, w_142_181);
  not1 I250_239(w_250_239, w_238_120);
  not1 I250_252(w_250_252, w_046_545);
  or2  I250_287(w_250_287, w_148_417, w_246_607);
  or2  I250_288(w_250_288, w_005_234, w_186_095);
  or2  I250_292(w_250_292, w_079_060, w_085_205);
  and2 I250_327(w_250_327, w_193_199, w_065_185);
  and2 I250_367(w_250_367, w_135_019, w_145_027);
  not1 I250_513(w_250_513, w_092_292);
  not1 I250_548(w_250_548, w_011_265);
  or2  I250_588(w_250_588, w_215_024, w_172_002);
  not1 I250_605(w_250_605, w_030_324);
  not1 I250_609(w_250_609, w_119_082);
  and2 I251_013(w_251_013, w_208_133, w_125_079);
  or2  I251_017(w_251_017, w_155_352, w_062_554);
  nand2 I251_028(w_251_028, w_198_076, w_218_189);
  and2 I251_035(w_251_035, w_197_223, w_018_022);
  not1 I251_037(w_251_037, w_234_326);
  nand2 I251_047(w_251_047, w_087_358, w_013_229);
  nand2 I251_048(w_251_048, w_097_502, w_249_191);
  nand2 I251_064(w_251_064, w_215_138, w_091_154);
  or2  I251_075(w_251_075, w_024_099, w_110_132);
  or2  I251_081(w_251_081, w_236_166, w_232_399);
  and2 I251_089(w_251_089, w_198_059, w_037_212);
  not1 I251_097(w_251_097, w_174_014);
  not1 I251_109(w_251_109, w_080_478);
  or2  I251_112(w_251_112, w_008_071, w_014_248);
  and2 I251_130(w_251_130, w_110_090, w_144_373);
  nand2 I251_131(w_251_131, w_083_127, w_241_068);
  and2 I251_133(w_251_133, w_178_009, w_104_007);
  nand2 I252_012(w_252_012, w_057_002, w_161_009);
  not1 I252_044(w_252_044, w_026_139);
  and2 I252_065(w_252_065, w_037_155, w_161_514);
  or2  I252_088(w_252_088, w_178_036, w_109_486);
  nand2 I252_103(w_252_103, w_138_261, w_241_011);
  nand2 I252_124(w_252_124, w_137_061, w_163_077);
  not1 I252_229(w_252_229, w_220_340);
  nand2 I252_242(w_252_242, w_069_143, w_124_244);
  or2  I252_247(w_252_247, w_004_397, w_072_070);
  not1 I252_272(w_252_272, w_172_007);
  or2  I252_275(w_252_275, w_122_067, w_026_007);
  not1 I252_280(w_252_280, w_222_315);
  not1 I252_301(w_252_301, w_221_069);
  or2  I252_306(w_252_306, w_010_660, w_011_141);
  and2 I252_331(w_252_331, w_086_093, w_180_025);
  nand2 I252_363(w_252_363, w_157_013, w_105_264);
  and2 I252_368(w_252_368, w_068_276, w_077_597);
  not1 I252_386(w_252_386, w_123_302);
  nand2 I252_394(w_252_394, w_218_701, w_222_026);
  or2  I252_428(w_252_430, w_252_429, w_023_007);
  and2 I252_429(w_252_431, w_247_107, w_252_430);
  nand2 I252_430(w_252_432, w_252_431, w_126_068);
  nand2 I252_431(w_252_433, w_077_011, w_252_432);
  not1 I252_432(w_252_434, w_252_433);
  not1 I252_433(w_252_435, w_252_434);
  and2 I252_434(w_252_436, w_252_435, w_209_314);
  and2 I252_435(w_252_437, w_252_436, w_188_592);
  nand2 I252_436(w_252_429, w_252_437, w_250_327);
  and2 I253_002(w_253_002, w_246_075, w_201_174);
  and2 I253_008(w_253_008, w_038_143, w_225_142);
  not1 I253_023(w_253_023, w_201_081);
  and2 I253_053(w_253_053, w_228_039, w_184_041);
  not1 I253_059(w_253_059, w_110_154);
  not1 I253_060(w_253_060, w_171_654);
  and2 I253_074(w_253_074, w_175_108, w_144_306);
  and2 I253_143(w_253_143, w_060_098, w_006_192);
  nand2 I253_150(w_253_150, w_028_240, w_094_514);
  and2 I253_163(w_253_163, w_193_312, w_192_065);
  or2  I253_198(w_253_198, w_082_150, w_127_000);
  nand2 I253_221(w_253_221, w_149_612, w_169_008);
  nand2 I253_318(w_253_318, w_156_044, w_187_006);
  or2  I253_344(w_253_344, w_164_235, w_241_002);
  and2 I253_361(w_253_361, w_110_294, w_035_022);
  and2 I253_363(w_253_363, w_237_134, w_177_036);
  not1 I253_415(w_253_415, w_213_577);
  not1 I254_000(w_254_000, w_085_051);
  or2  I254_020(w_254_020, w_136_040, w_057_243);
  not1 I254_028(w_254_028, w_127_007);
  not1 I254_031(w_254_031, w_043_032);
  and2 I254_037(w_254_037, w_040_488, w_090_306);
  not1 I254_053(w_254_053, w_016_005);
  or2  I254_054(w_254_054, w_130_220, w_054_508);
  and2 I254_057(w_254_057, w_056_016, w_085_167);
  or2  I254_058(w_254_058, w_021_238, w_029_081);
  nand2 I254_061(w_254_061, w_015_061, w_142_209);
  nand2 I254_062(w_254_062, w_253_008, w_155_444);
  or2  I254_065(w_254_065, w_021_056, w_030_377);
  or2  I254_073(w_254_073, w_253_002, w_097_471);
  nand2 I254_084(w_254_084, w_143_652, w_223_284);
  not1 I254_095(w_254_095, w_135_078);
  nand2 I254_104(w_254_106, w_254_105, w_013_523);
  nand2 I254_105(w_254_107, w_222_315, w_254_106);
  or2  I254_106(w_254_108, w_165_096, w_254_107);
  nand2 I254_107(w_254_109, w_045_258, w_254_108);
  or2  I254_108(w_254_110, w_254_109, w_169_106);
  nand2 I254_109(w_254_111, w_254_110, w_079_036);
  nand2 I254_110(w_254_112, w_254_111, w_149_126);
  and2 I254_111(w_254_113, w_241_010, w_254_112);
  not1 I254_112(w_254_105, w_254_113);
  nand2 I255_024(w_255_024, w_240_159, w_003_050);
  not1 I255_035(w_255_035, w_117_088);
  not1 I255_042(w_255_042, w_059_066);
  not1 I255_062(w_255_062, w_067_318);
  and2 I255_076(w_255_076, w_069_029, w_168_492);
  and2 I255_078(w_255_078, w_208_021, w_195_141);
  not1 I255_081(w_255_081, w_123_297);
  and2 I255_089(w_255_089, w_021_191, w_153_052);
  nand2 I255_103(w_255_103, w_009_096, w_108_159);
  and2 I255_105(w_255_105, w_058_352, w_188_039);
  not1 I256_021(w_256_021, w_092_009);
  not1 I256_028(w_256_028, w_000_524);
  and2 I256_060(w_256_060, w_162_015, w_117_079);
  and2 I256_089(w_256_089, w_023_093, w_229_247);
  or2  I256_097(w_256_097, w_130_408, w_053_109);
  or2  I256_310(w_256_310, w_077_178, w_127_067);
  not1 I256_477(w_256_477, w_173_001);
  and2 I256_484(w_256_484, w_042_043, w_209_299);
  and2 I256_490(w_256_490, w_126_028, w_048_000);
  nand2 I256_515(w_256_515, w_203_368, w_231_537);
  or2  I256_550(w_256_550, w_076_459, w_002_493);
  not1 I256_646(w_256_646, w_108_086);
  not1 I256_689(w_256_689, w_208_027);
  and2 I257_054(w_257_054, w_204_027, w_202_017);
  not1 I257_075(w_257_075, w_133_143);
  not1 I257_101(w_257_101, w_008_625);
  or2  I257_110(w_257_110, w_172_031, w_036_255);
  or2  I257_112(w_257_112, w_183_119, w_009_159);
  not1 I257_143(w_257_143, w_093_339);
  nand2 I257_190(w_257_190, w_172_040, w_029_025);
  or2  I257_243(w_257_243, w_113_316, w_180_024);
  nand2 I257_257(w_257_257, w_097_153, w_000_183);
  not1 I257_293(w_257_293, w_100_086);
  not1 I257_318(w_257_318, w_189_220);
  nand2 I258_026(w_258_026, w_081_014, w_017_251);
  not1 I258_032(w_258_032, w_059_702);
  not1 I258_103(w_258_103, w_195_140);
  or2  I258_138(w_258_138, w_198_052, w_017_107);
  not1 I258_153(w_258_153, w_224_049);
  not1 I258_193(w_258_193, w_064_229);
  nand2 I258_240(w_258_240, w_232_376, w_137_075);
  and2 I258_247(w_258_247, w_008_009, w_014_189);
  not1 I258_390(w_258_390, w_019_014);
  not1 I258_411(w_258_411, w_028_551);
  or2  I258_449(w_258_449, w_109_169, w_016_006);
  or2  I258_481(w_258_481, w_143_554, w_170_139);
  not1 I259_038(w_259_038, w_216_169);
  and2 I259_084(w_259_084, w_120_681, w_041_306);
  or2  I259_131(w_259_131, w_064_004, w_228_105);
  or2  I259_224(w_259_224, w_088_117, w_195_121);
  nand2 I259_316(w_259_316, w_057_055, w_131_092);
  or2  I259_338(w_259_338, w_245_397, w_128_035);
  not1 I259_345(w_259_345, w_187_016);
  nand2 I259_457(w_259_457, w_160_449, w_252_088);
  or2  I259_469(w_259_469, w_058_589, w_101_166);
  or2  I259_472(w_259_472, w_115_019, w_163_497);
  and2 I259_506(w_259_506, w_128_000, w_018_036);
  not1 I259_543(w_259_543, w_059_489);
  nand2 I259_551(w_259_551, w_251_109, w_009_229);
  nand2 I260_001(w_260_001, w_155_090, w_215_038);
  nand2 I260_017(w_260_017, w_092_331, w_193_014);
  nand2 I260_027(w_260_027, w_015_103, w_203_184);
  not1 I260_030(w_260_030, w_071_299);
  or2  I260_035(w_260_035, w_205_216, w_190_112);
  nand2 I260_058(w_260_058, w_218_080, w_178_097);
  and2 I260_061(w_260_061, w_042_377, w_076_375);
  or2  I260_082(w_260_082, w_201_502, w_250_239);
  nand2 I260_101(w_260_101, w_004_140, w_201_422);
  and2 I260_108(w_260_108, w_247_021, w_096_001);
  or2  I260_151(w_260_151, w_213_070, w_032_150);
  and2 I260_159(w_260_159, w_214_055, w_054_542);
  or2  I260_161(w_260_161, w_036_085, w_230_055);
  and2 I260_164(w_260_164, w_194_102, w_231_463);
  nand2 I260_166(w_260_166, w_251_133, w_117_038);
  not1 I260_183(w_260_183, w_095_051);
  nand2 I260_199(w_260_199, w_227_173, w_008_249);
  and2 I260_201(w_260_201, w_251_112, w_213_358);
  not1 I260_281(w_260_283, w_260_282);
  not1 I260_282(w_260_284, w_260_283);
  or2  I260_283(w_260_285, w_040_054, w_260_284);
  or2  I260_284(w_260_286, w_260_285, w_021_144);
  not1 I260_285(w_260_287, w_260_286);
  and2 I260_286(w_260_288, w_253_053, w_260_287);
  and2 I260_287(w_260_282, w_260_304, w_260_288);
  and2 I260_288(w_260_293, w_047_147, w_260_292);
  and2 I260_289(w_260_294, w_260_293, w_205_066);
  not1 I260_290(w_260_295, w_260_294);
  not1 I260_291(w_260_296, w_260_295);
  not1 I260_292(w_260_297, w_260_296);
  nand2 I260_293(w_260_298, w_098_015, w_260_297);
  or2  I260_294(w_260_299, w_127_073, w_260_298);
  and2 I260_295(w_260_300, w_143_014, w_260_299);
  not1 I260_296(w_260_301, w_260_300);
  and2 I260_297(w_260_302, w_162_023, w_260_301);
  not1 I260_298(w_260_292, w_260_282);
  and2 I260_299(w_260_304, w_180_026, w_260_302);
  nand2 I261_000(w_261_000, w_185_049, w_027_093);
  or2  I261_005(w_261_005, w_160_634, w_202_198);
  not1 I261_008(w_261_008, w_235_034);
  not1 I261_015(w_261_015, w_247_000);
  and2 I261_022(w_261_022, w_096_002, w_017_104);
  or2  I261_029(w_261_029, w_129_329, w_214_203);
  and2 I261_032(w_261_032, w_082_059, w_199_178);
  nand2 I261_034(w_261_034, w_051_282, w_004_297);
  or2  I261_041(w_261_041, w_259_084, w_129_204);
  or2  I261_044(w_261_044, w_005_157, w_120_177);
  or2  I261_061(w_261_061, w_066_040, w_013_346);
  nand2 I261_100(w_261_100, w_200_254, w_036_207);
  not1 I262_001(w_262_001, w_000_435);
  and2 I262_002(w_262_002, w_194_314, w_132_129);
  or2  I262_010(w_262_010, w_128_026, w_180_011);
  nand2 I262_044(w_262_044, w_227_647, w_181_039);
  and2 I262_068(w_262_068, w_044_435, w_037_110);
  or2  I262_073(w_262_073, w_252_044, w_026_173);
  or2  I262_202(w_262_202, w_249_333, w_139_024);
  and2 I262_223(w_262_223, w_208_214, w_100_113);
  and2 I262_267(w_262_267, w_102_329, w_024_048);
  or2  I262_321(w_262_321, w_080_065, w_128_022);
  not1 I262_371(w_262_371, w_062_516);
  nand2 I262_381(w_262_381, w_001_001, w_038_429);
  not1 I262_389(w_262_389, w_231_321);
  not1 I263_001(w_263_001, w_158_002);
  and2 I263_007(w_263_007, w_223_140, w_240_142);
  not1 I263_022(w_263_022, w_179_079);
  and2 I263_028(w_263_028, w_120_348, w_113_262);
  nand2 I263_030(w_263_030, w_002_058, w_204_510);
  not1 I263_049(w_263_049, w_057_137);
  nand2 I263_062(w_263_062, w_195_044, w_209_065);
  or2  I263_078(w_263_078, w_254_062, w_000_381);
  nand2 I263_083(w_263_083, w_045_270, w_216_203);
  or2  I263_101(w_263_101, w_242_058, w_210_040);
  and2 I263_104(w_263_104, w_246_289, w_192_163);
  and2 I263_106(w_263_106, w_182_024, w_126_117);
  and2 I263_119(w_263_119, w_143_019, w_184_029);
  not1 I263_120(w_263_120, w_021_189);
  not1 I263_133(w_263_133, w_031_386);
  not1 I264_157(w_264_157, w_065_344);
  nand2 I264_159(w_264_159, w_169_221, w_089_167);
  not1 I264_161(w_264_161, w_229_015);
  and2 I264_233(w_264_233, w_159_063, w_202_040);
  nand2 I264_266(w_264_266, w_139_001, w_008_216);
  nand2 I264_273(w_264_273, w_073_203, w_098_012);
  nand2 I264_310(w_264_310, w_103_136, w_082_303);
  and2 I264_470(w_264_470, w_228_578, w_034_063);
  nand2 I264_553(w_264_553, w_097_225, w_027_168);
  or2  I264_599(w_264_599, w_124_330, w_259_338);
  or2  I264_666(w_264_666, w_048_012, w_120_305);
  not1 I264_743(w_264_743, w_221_159);
  nand2 I265_029(w_265_029, w_020_023, w_064_180);
  not1 I265_064(w_265_064, w_012_274);
  and2 I265_073(w_265_073, w_068_206, w_064_286);
  or2  I265_120(w_265_120, w_193_006, w_097_507);
  or2  I265_171(w_265_171, w_243_160, w_172_006);
  not1 I265_197(w_265_197, w_229_003);
  and2 I265_237(w_265_237, w_256_490, w_009_066);
  nand2 I265_327(w_265_327, w_131_037, w_077_590);
  not1 I265_418(w_265_418, w_079_048);
  not1 I265_450(w_265_450, w_217_018);
  not1 I265_453(w_265_453, w_223_156);
  nand2 I265_491(w_265_491, w_130_195, w_200_005);
  or2  I265_507(w_265_507, w_015_416, w_033_380);
  or2  I265_641(w_265_641, w_100_080, w_078_050);
  or2  I265_645(w_265_645, w_002_427, w_016_001);
  nand2 I265_694(w_265_694, w_135_257, w_067_083);
  or2  I266_043(w_266_043, w_195_067, w_178_102);
  and2 I266_124(w_266_124, w_121_011, w_009_042);
  not1 I266_160(w_266_160, w_042_052);
  nand2 I266_176(w_266_176, w_244_244, w_119_106);
  not1 I266_247(w_266_247, w_122_014);
  nand2 I266_250(w_266_250, w_081_003, w_122_086);
  nand2 I266_307(w_266_307, w_017_480, w_206_203);
  and2 I266_324(w_266_324, w_167_016, w_051_028);
  or2  I266_330(w_266_330, w_234_147, w_015_068);
  not1 I266_438(w_266_438, w_049_348);
  not1 I266_533(w_266_533, w_175_056);
  or2  I266_620(w_266_622, w_093_420, w_266_621);
  not1 I266_621(w_266_623, w_266_622);
  not1 I266_622(w_266_624, w_266_623);
  not1 I266_623(w_266_625, w_266_624);
  and2 I266_624(w_266_626, w_266_625, w_266_645);
  or2  I266_625(w_266_627, w_266_626, w_072_012);
  and2 I266_626(w_266_628, w_215_249, w_266_627);
  or2  I266_627(w_266_629, w_266_628, w_099_057);
  and2 I266_628(w_266_630, w_266_629, w_070_384);
  and2 I266_629(w_266_631, w_266_630, w_061_452);
  nand2 I266_630(w_266_621, w_266_631, w_134_218);
  or2  I266_631(w_266_636, w_266_635, w_011_009);
  not1 I266_632(w_266_637, w_266_636);
  and2 I266_633(w_266_638, w_266_637, w_012_187);
  and2 I266_634(w_266_639, w_240_056, w_266_638);
  or2  I266_635(w_266_640, w_119_189, w_266_639);
  or2  I266_636(w_266_641, w_266_640, w_027_113);
  and2 I266_637(w_266_642, w_266_641, w_096_000);
  and2 I266_638(w_266_643, w_266_642, w_148_670);
  not1 I266_639(w_266_635, w_266_626);
  and2 I266_640(w_266_645, w_168_216, w_266_643);
  or2  I267_014(w_267_014, w_219_008, w_233_068);
  nand2 I267_023(w_267_023, w_069_093, w_032_174);
  or2  I267_041(w_267_041, w_091_119, w_212_087);
  and2 I267_054(w_267_054, w_079_003, w_126_041);
  not1 I267_055(w_267_055, w_194_102);
  not1 I267_065(w_267_065, w_039_657);
  and2 I267_067(w_267_067, w_042_389, w_113_218);
  and2 I267_083(w_267_083, w_175_018, w_171_303);
  not1 I267_085(w_267_085, w_039_029);
  nand2 I267_103(w_267_103, w_075_120, w_123_367);
  not1 I267_114(w_267_114, w_255_105);
  not1 I267_131(w_267_131, w_117_057);
  nand2 I267_146(w_267_146, w_028_140, w_262_044);
  or2  I267_155(w_267_155, w_073_554, w_050_602);
  or2  I267_183(w_267_183, w_067_069, w_212_009);
  nand2 I267_216(w_267_216, w_162_006, w_101_124);
  and2 I267_217(w_267_217, w_189_157, w_215_487);
  nand2 I267_248(w_267_248, w_057_239, w_189_546);
  or2  I267_276(w_267_276, w_245_436, w_168_151);
  or2  I267_298(w_267_298, w_001_021, w_043_030);
  nand2 I268_021(w_268_021, w_031_076, w_262_001);
  and2 I268_035(w_268_035, w_191_331, w_229_455);
  not1 I268_038(w_268_038, w_249_169);
  not1 I268_058(w_268_058, w_150_009);
  and2 I268_079(w_268_079, w_197_194, w_081_007);
  not1 I268_113(w_268_113, w_249_187);
  not1 I268_152(w_268_152, w_017_262);
  nand2 I268_213(w_268_213, w_016_000, w_210_142);
  nand2 I268_214(w_268_214, w_225_104, w_146_302);
  and2 I268_216(w_268_216, w_012_088, w_262_389);
  nand2 I268_237(w_268_237, w_203_430, w_062_430);
  and2 I268_261(w_268_261, w_149_302, w_013_369);
  not1 I268_268(w_268_268, w_160_059);
  or2  I269_019(w_269_019, w_119_001, w_259_316);
  and2 I269_030(w_269_030, w_118_043, w_015_272);
  or2  I269_070(w_269_070, w_030_326, w_115_000);
  or2  I269_122(w_269_122, w_215_015, w_188_393);
  or2  I269_159(w_269_159, w_240_026, w_148_499);
  nand2 I269_171(w_269_171, w_114_067, w_024_503);
  or2  I269_276(w_269_276, w_202_186, w_225_010);
  nand2 I269_356(w_269_356, w_042_340, w_008_376);
  or2  I269_363(w_269_363, w_076_102, w_078_571);
  or2  I269_382(w_269_382, w_063_238, w_182_004);
  or2  I269_405(w_269_405, w_246_119, w_131_557);
  not1 I269_414(w_269_414, w_248_034);
  and2 I269_434(w_269_434, w_054_082, w_216_088);
  nand2 I269_441(w_269_441, w_150_318, w_040_268);
  or2  I269_493(w_269_493, w_137_272, w_081_020);
  and2 I269_564(w_269_564, w_197_445, w_146_036);
  nand2 I269_565(w_269_565, w_032_283, w_214_518);
  nand2 I270_017(w_270_017, w_220_371, w_119_162);
  nand2 I270_037(w_270_037, w_060_308, w_098_013);
  or2  I270_046(w_270_046, w_024_436, w_161_153);
  nand2 I270_217(w_270_217, w_140_042, w_121_144);
  nand2 I270_228(w_270_228, w_269_434, w_081_001);
  not1 I270_284(w_270_284, w_080_033);
  and2 I270_335(w_270_335, w_177_405, w_051_378);
  nand2 I271_011(w_271_011, w_187_041, w_053_034);
  nand2 I271_021(w_271_021, w_056_244, w_148_565);
  not1 I271_030(w_271_030, w_036_192);
  and2 I271_072(w_271_072, w_073_493, w_137_188);
  and2 I271_142(w_271_142, w_227_269, w_079_015);
  nand2 I271_188(w_271_188, w_092_151, w_250_287);
  or2  I271_354(w_271_354, w_147_202, w_020_042);
  not1 I271_416(w_271_416, w_003_027);
  or2  I271_470(w_271_470, w_004_000, w_251_028);
  nand2 I271_532(w_271_532, w_090_086, w_155_402);
  and2 I271_555(w_271_555, w_126_154, w_101_038);
  nand2 I271_575(w_271_575, w_102_368, w_156_209);
  not1 I271_602(w_271_602, w_087_292);
  nand2 I271_637(w_271_637, w_226_092, w_101_006);
  or2  I271_740(w_271_740, w_032_310, w_240_072);
  not1 I272_005(w_272_005, w_091_151);
  and2 I272_009(w_272_009, w_154_062, w_161_394);
  and2 I272_018(w_272_018, w_187_015, w_240_076);
  and2 I272_021(w_272_021, w_085_074, w_099_001);
  or2  I272_024(w_272_024, w_020_196, w_221_213);
  or2  I272_026(w_272_026, w_196_196, w_261_008);
  nand2 I272_028(w_272_028, w_154_060, w_031_236);
  nand2 I272_030(w_272_030, w_053_033, w_212_170);
  or2  I272_031(w_272_031, w_161_093, w_004_144);
  not1 I272_038(w_272_038, w_038_325);
  not1 I272_039(w_272_039, w_036_319);
  and2 I272_040(w_272_040, w_103_002, w_062_518);
  and2 I272_043(w_272_043, w_026_179, w_216_362);
  not1 I273_042(w_273_042, w_252_275);
  or2  I273_054(w_273_054, w_219_626, w_244_200);
  not1 I273_065(w_273_065, w_259_131);
  not1 I273_075(w_273_075, w_108_035);
  nand2 I273_092(w_273_092, w_128_157, w_074_159);
  or2  I273_093(w_273_093, w_264_161, w_075_062);
  not1 I273_105(w_273_105, w_123_532);
  or2  I273_112(w_273_112, w_012_268, w_261_022);
  or2  I273_133(w_273_135, w_152_167, w_273_134);
  or2  I273_134(w_273_136, w_273_135, w_084_004);
  and2 I273_135(w_273_137, w_273_136, w_058_664);
  and2 I273_136(w_273_138, w_273_137, w_245_398);
  not1 I273_137(w_273_139, w_273_138);
  not1 I273_138(w_273_140, w_273_139);
  or2  I273_139(w_273_141, w_155_493, w_273_140);
  and2 I273_140(w_273_142, w_273_141, w_005_166);
  and2 I273_141(w_273_134, w_207_069, w_273_142);
  nand2 I274_029(w_274_029, w_118_023, w_239_000);
  not1 I274_055(w_274_055, w_244_205);
  and2 I274_100(w_274_100, w_182_005, w_130_264);
  or2  I274_104(w_274_104, w_098_045, w_062_689);
  or2  I274_115(w_274_115, w_232_381, w_189_319);
  not1 I274_126(w_274_126, w_227_584);
  not1 I274_130(w_274_130, w_176_001);
  not1 I274_143(w_274_143, w_207_189);
  not1 I274_144(w_274_144, w_042_232);
  and2 I274_149(w_274_149, w_225_154, w_114_134);
  and2 I274_170(w_274_170, w_211_014, w_263_104);
  nand2 I274_171(w_274_171, w_054_305, w_038_602);
  nand2 I274_188(w_274_188, w_024_284, w_232_295);
  not1 I274_221(w_274_221, w_065_387);
  and2 I274_232(w_274_232, w_084_047, w_268_213);
  or2  I274_238(w_274_238, w_238_141, w_215_203);
  not1 I275_049(w_275_049, w_099_123);
  or2  I275_090(w_275_090, w_081_020, w_078_306);
  and2 I275_133(w_275_133, w_176_148, w_003_079);
  or2  I275_135(w_275_135, w_139_021, w_191_134);
  or2  I275_291(w_275_291, w_201_409, w_219_005);
  nand2 I275_489(w_275_489, w_128_051, w_263_030);
  or2  I275_598(w_275_598, w_008_244, w_004_091);
  or2  I275_603(w_275_603, w_020_184, w_256_060);
  and2 I275_605(w_275_605, w_168_506, w_217_001);
  or2  I275_619(w_275_619, w_097_102, w_142_101);
  not1 I275_722(w_275_722, w_024_105);
  or2  I276_030(w_276_030, w_115_190, w_124_052);
  or2  I276_050(w_276_050, w_252_301, w_074_041);
  nand2 I276_110(w_276_110, w_199_338, w_150_003);
  and2 I276_142(w_276_142, w_239_000, w_122_030);
  nand2 I276_170(w_276_170, w_044_248, w_079_055);
  or2  I276_185(w_276_185, w_080_440, w_270_046);
  not1 I276_196(w_276_196, w_244_000);
  nand2 I276_200(w_276_200, w_052_009, w_143_300);
  not1 I276_264(w_276_264, w_165_017);
  or2  I276_296(w_276_296, w_082_135, w_025_180);
  and2 I276_326(w_276_326, w_135_062, w_235_112);
  and2 I276_331(w_276_331, w_195_007, w_035_121);
  not1 I276_349(w_276_349, w_168_448);
  nand2 I276_350(w_276_350, w_143_530, w_134_116);
  and2 I276_367(w_276_367, w_129_295, w_220_337);
  or2  I277_013(w_277_013, w_202_267, w_188_036);
  nand2 I277_020(w_277_020, w_047_311, w_202_223);
  or2  I277_038(w_277_038, w_009_000, w_014_056);
  nand2 I277_067(w_277_067, w_162_013, w_024_509);
  and2 I277_123(w_277_123, w_007_237, w_240_055);
  not1 I277_137(w_277_137, w_177_266);
  not1 I277_143(w_277_143, w_185_027);
  not1 I277_203(w_277_203, w_010_174);
  and2 I277_258(w_277_258, w_168_159, w_188_184);
  not1 I277_268(w_277_268, w_149_015);
  nand2 I277_293(w_277_293, w_051_126, w_171_221);
  or2  I277_315(w_277_315, w_079_024, w_084_001);
  or2  I277_317(w_277_317, w_083_093, w_139_027);
  nand2 I277_364(w_277_364, w_048_002, w_197_114);
  nand2 I277_373(w_277_373, w_153_020, w_223_202);
  nand2 I277_381(w_277_381, w_174_083, w_143_111);
  nand2 I278_045(w_278_045, w_058_238, w_232_172);
  not1 I278_057(w_278_057, w_039_396);
  and2 I278_060(w_278_060, w_001_026, w_262_223);
  and2 I278_100(w_278_100, w_264_553, w_007_198);
  nand2 I278_116(w_278_116, w_213_085, w_199_294);
  or2  I278_174(w_278_174, w_130_254, w_090_472);
  nand2 I279_026(w_279_026, w_133_374, w_192_119);
  and2 I279_068(w_279_068, w_157_074, w_048_013);
  not1 I279_069(w_279_069, w_202_078);
  and2 I279_124(w_279_124, w_222_236, w_118_050);
  nand2 I279_127(w_279_127, w_205_504, w_166_138);
  nand2 I279_138(w_279_138, w_128_297, w_032_597);
  nand2 I279_139(w_279_139, w_017_232, w_199_267);
  or2  I279_153(w_279_153, w_161_135, w_035_046);
  and2 I279_160(w_279_160, w_029_001, w_122_026);
  and2 I279_171(w_279_171, w_183_031, w_091_085);
  nand2 I279_228(w_279_228, w_038_162, w_085_294);
  nand2 I279_253(w_279_253, w_260_164, w_190_029);
  not1 I279_302(w_279_302, w_132_206);
  or2  I280_019(w_280_019, w_222_141, w_158_001);
  nand2 I280_098(w_280_098, w_120_072, w_209_063);
  not1 I280_258(w_280_258, w_004_180);
  nand2 I280_259(w_280_259, w_272_005, w_219_244);
  and2 I280_282(w_280_282, w_151_366, w_179_023);
  or2  I280_306(w_280_306, w_189_157, w_141_154);
  not1 I280_444(w_280_444, w_187_028);
  nand2 I280_448(w_280_448, w_110_092, w_220_265);
  or2  I280_503(w_280_503, w_233_234, w_157_141);
  and2 I280_559(w_280_559, w_237_033, w_187_032);
  not1 I280_652(w_280_652, w_191_286);
  and2 I280_682(w_280_682, w_090_275, w_109_259);
  or2  I280_687(w_280_687, w_215_166, w_111_018);
  and2 I281_044(w_281_044, w_267_023, w_186_055);
  and2 I281_089(w_281_089, w_067_344, w_198_046);
  and2 I281_119(w_281_119, w_034_020, w_078_150);
  and2 I281_133(w_281_133, w_008_011, w_017_453);
  and2 I281_212(w_281_212, w_069_227, w_011_599);
  not1 I281_237(w_281_237, w_093_006);
  or2  I281_283(w_281_283, w_234_086, w_092_447);
  not1 I281_307(w_281_307, w_030_251);
  or2  I281_365(w_281_365, w_175_022, w_185_069);
  and2 I281_389(w_281_389, w_044_587, w_266_176);
  nand2 I281_462(w_281_462, w_006_236, w_155_470);
  and2 I281_551(w_281_551, w_056_176, w_212_124);
  nand2 I281_616(w_281_616, w_248_130, w_168_143);
  and2 I281_627(w_281_627, w_190_053, w_026_188);
  nand2 I281_643(w_281_643, w_265_453, w_085_340);
  and2 I281_710(w_281_710, w_266_250, w_068_074);
  and2 I281_740(w_281_740, w_213_079, w_148_038);
  or2  I282_031(w_282_031, w_199_280, w_239_000);
  not1 I282_109(w_282_109, w_274_115);
  nand2 I282_110(w_282_110, w_233_353, w_187_017);
  nand2 I282_137(w_282_137, w_084_015, w_107_256);
  not1 I282_141(w_282_141, w_258_103);
  nand2 I282_150(w_282_150, w_226_019, w_190_096);
  not1 I282_166(w_282_166, w_208_053);
  and2 I282_206(w_282_206, w_115_191, w_080_023);
  not1 I282_227(w_282_227, w_193_085);
  or2  I282_236(w_282_236, w_137_104, w_202_149);
  nand2 I282_246(w_282_246, w_265_197, w_089_128);
  not1 I282_250(w_282_250, w_197_060);
  and2 I282_265(w_282_265, w_234_038, w_122_066);
  not1 I282_291(w_282_291, w_032_295);
  not1 I282_298(w_282_298, w_008_240);
  or2  I282_327(w_282_327, w_160_405, w_040_464);
  nand2 I282_367(w_282_367, w_180_008, w_128_055);
  not1 I282_384(w_282_386, w_282_385);
  not1 I282_385(w_282_387, w_282_386);
  and2 I282_386(w_282_388, w_282_387, w_200_429);
  nand2 I282_387(w_282_385, w_282_388, w_282_397);
  and2 I282_388(w_282_393, w_282_392, w_192_138);
  and2 I282_389(w_282_394, w_282_393, w_044_110);
  and2 I282_390(w_282_395, w_214_448, w_282_394);
  not1 I282_391(w_282_392, w_282_385);
  and2 I282_392(w_282_397, w_048_009, w_282_395);
  not1 I283_003(w_283_003, w_095_054);
  or2  I283_038(w_283_038, w_083_163, w_163_221);
  and2 I283_043(w_283_043, w_120_558, w_013_065);
  not1 I283_064(w_283_064, w_114_069);
  or2  I283_094(w_283_094, w_136_033, w_015_162);
  not1 I283_126(w_283_126, w_201_148);
  and2 I283_131(w_283_131, w_016_006, w_211_028);
  and2 I283_137(w_283_137, w_130_391, w_099_037);
  and2 I283_138(w_283_138, w_027_142, w_202_119);
  and2 I283_216(w_283_216, w_126_041, w_199_266);
  or2  I283_219(w_283_219, w_016_005, w_282_250);
  and2 I283_272(w_283_272, w_252_331, w_045_169);
  or2  I283_329(w_283_329, w_234_153, w_280_682);
  not1 I283_338(w_283_338, w_056_462);
  or2  I283_379(w_283_379, w_036_002, w_044_000);
  nand2 I284_005(w_284_005, w_193_299, w_169_004);
  or2  I284_014(w_284_014, w_185_130, w_208_122);
  not1 I284_015(w_284_015, w_212_165);
  not1 I284_022(w_284_022, w_283_338);
  and2 I284_024(w_284_024, w_271_470, w_077_150);
  nand2 I284_029(w_284_029, w_084_007, w_232_035);
  or2  I284_039(w_284_039, w_115_021, w_209_263);
  or2  I284_040(w_284_040, w_091_088, w_217_051);
  or2  I284_049(w_284_049, w_136_014, w_163_478);
  not1 I284_054(w_284_054, w_145_039);
  nand2 I284_080(w_284_080, w_213_046, w_059_430);
  and2 I284_081(w_284_081, w_268_261, w_030_275);
  nand2 I284_102(w_284_102, w_042_184, w_169_062);
  not1 I284_113(w_284_113, w_088_065);
  and2 I284_123(w_284_123, w_238_150, w_236_159);
  not1 I284_129(w_284_129, w_132_115);
  nand2 I284_142(w_284_142, w_204_280, w_098_024);
  or2  I284_145(w_284_145, w_208_408, w_229_192);
  not1 I285_011(w_285_011, w_095_052);
  not1 I285_037(w_285_037, w_043_036);
  nand2 I285_041(w_285_041, w_218_338, w_134_072);
  nand2 I285_057(w_285_057, w_129_276, w_142_638);
  not1 I285_091(w_285_091, w_093_123);
  and2 I285_104(w_285_104, w_172_024, w_096_002);
  not1 I285_184(w_285_184, w_099_173);
  not1 I285_353(w_285_353, w_095_040);
  nand2 I285_393(w_285_393, w_171_322, w_157_007);
  or2  I285_460(w_285_460, w_282_109, w_235_083);
  nand2 I285_689(w_285_689, w_277_381, w_137_162);
  and2 I285_774(w_285_774, w_037_223, w_105_251);
  nand2 I286_037(w_286_037, w_128_318, w_139_025);
  or2  I286_074(w_286_074, w_233_326, w_029_094);
  not1 I286_130(w_286_130, w_146_213);
  not1 I286_132(w_286_132, w_141_011);
  or2  I286_136(w_286_136, w_111_021, w_220_377);
  or2  I286_186(w_286_186, w_028_120, w_167_152);
  not1 I286_190(w_286_190, w_120_332);
  and2 I286_275(w_286_275, w_270_228, w_223_184);
  not1 I286_362(w_286_362, w_054_284);
  and2 I286_377(w_286_377, w_048_012, w_215_099);
  and2 I286_380(w_286_380, w_261_005, w_187_009);
  or2  I286_393(w_286_393, w_071_294, w_196_023);
  nand2 I287_019(w_287_019, w_132_076, w_050_573);
  and2 I287_020(w_287_020, w_031_472, w_025_172);
  and2 I287_064(w_287_064, w_208_026, w_032_232);
  nand2 I287_125(w_287_125, w_000_076, w_282_227);
  and2 I287_180(w_287_180, w_112_085, w_206_086);
  not1 I287_274(w_287_274, w_231_427);
  or2  I287_279(w_287_279, w_031_340, w_049_358);
  not1 I287_315(w_287_315, w_106_107);
  or2  I287_334(w_287_334, w_172_040, w_276_185);
  or2  I287_335(w_287_335, w_011_583, w_232_150);
  or2  I287_354(w_287_354, w_214_201, w_120_159);
  not1 I287_369(w_287_369, w_219_668);
  nand2 I287_394(w_287_394, w_163_185, w_189_026);
  not1 I288_068(w_288_068, w_098_017);
  not1 I288_070(w_288_070, w_155_405);
  or2  I288_087(w_288_087, w_127_065, w_258_240);
  and2 I288_158(w_288_158, w_203_062, w_253_150);
  and2 I288_167(w_288_167, w_185_023, w_076_262);
  not1 I288_194(w_288_194, w_156_167);
  nand2 I288_198(w_288_198, w_221_207, w_167_080);
  or2  I288_278(w_288_278, w_234_195, w_038_484);
  and2 I288_288(w_288_288, w_128_608, w_168_232);
  and2 I288_420(w_288_420, w_212_120, w_189_367);
  or2  I288_422(w_288_422, w_023_087, w_087_205);
  or2  I288_478(w_288_478, w_114_015, w_088_013);
  not1 I288_509(w_288_511, w_288_510);
  and2 I288_510(w_288_512, w_288_511, w_288_526);
  and2 I288_511(w_288_510, w_093_504, w_288_512);
  not1 I288_512(w_288_517, w_288_516);
  not1 I288_513(w_288_518, w_288_517);
  and2 I288_514(w_288_519, w_180_016, w_288_518);
  and2 I288_515(w_288_520, w_152_511, w_288_519);
  nand2 I288_516(w_288_521, w_266_330, w_288_520);
  nand2 I288_517(w_288_522, w_068_082, w_288_521);
  and2 I288_518(w_288_523, w_288_522, w_007_051);
  and2 I288_519(w_288_524, w_265_171, w_288_523);
  not1 I288_520(w_288_516, w_288_512);
  and2 I288_521(w_288_526, w_254_028, w_288_524);
  not1 I289_103(w_289_103, w_106_075);
  not1 I289_121(w_289_121, w_064_093);
  and2 I289_166(w_289_166, w_056_012, w_148_087);
  nand2 I289_257(w_289_257, w_100_078, w_143_581);
  not1 I289_417(w_289_417, w_256_646);
  not1 I289_574(w_289_574, w_000_189);
  nand2 I290_004(w_290_004, w_264_233, w_143_479);
  and2 I290_005(w_290_005, w_108_087, w_231_530);
  nand2 I290_048(w_290_048, w_035_029, w_102_116);
  not1 I290_086(w_290_086, w_246_608);
  or2  I290_100(w_290_100, w_271_575, w_264_159);
  or2  I290_103(w_290_103, w_063_229, w_189_023);
  and2 I290_106(w_290_106, w_260_061, w_265_694);
  not1 I290_117(w_290_117, w_035_043);
  not1 I290_118(w_290_118, w_078_050);
  and2 I290_128(w_290_128, w_077_035, w_164_453);
  not1 I290_157(w_290_159, w_290_158);
  nand2 I290_158(w_290_160, w_290_159, w_175_615);
  or2  I290_159(w_290_161, w_290_160, w_289_166);
  nand2 I290_160(w_290_162, w_126_139, w_290_161);
  not1 I290_161(w_290_163, w_290_162);
  nand2 I290_162(w_290_164, w_286_132, w_290_163);
  nand2 I290_163(w_290_165, w_096_005, w_290_164);
  and2 I290_164(w_290_166, w_290_165, w_089_072);
  and2 I290_165(w_290_167, w_290_166, w_129_140);
  and2 I290_166(w_290_158, w_050_177, w_290_167);
  or2  I291_001(w_291_001, w_211_026, w_245_262);
  or2  I291_007(w_291_007, w_126_092, w_238_412);
  not1 I291_022(w_291_022, w_267_248);
  nand2 I291_030(w_291_030, w_042_034, w_004_241);
  and2 I291_043(w_291_043, w_166_097, w_117_050);
  not1 I291_044(w_291_044, w_224_303);
  not1 I291_063(w_291_063, w_218_725);
  and2 I291_071(w_291_071, w_150_394, w_072_123);
  nand2 I291_073(w_291_073, w_154_082, w_271_740);
  or2  I291_082(w_291_082, w_078_177, w_284_015);
  or2  I291_085(w_291_085, w_098_041, w_005_156);
  not1 I291_099(w_291_099, w_262_267);
  or2  I291_108(w_291_108, w_148_353, w_094_056);
  or2  I291_110(w_291_110, w_178_028, w_032_491);
  nand2 I291_123(w_291_123, w_152_008, w_151_011);
  not1 I291_129(w_291_129, w_137_032);
  and2 I292_033(w_292_033, w_190_067, w_286_074);
  or2  I292_298(w_292_298, w_140_020, w_275_722);
  and2 I292_309(w_292_309, w_003_059, w_084_038);
  and2 I292_433(w_292_433, w_189_175, w_274_238);
  and2 I292_494(w_292_494, w_276_349, w_166_123);
  or2  I292_533(w_292_533, w_203_016, w_019_020);
  not1 I292_554(w_292_554, w_226_190);
  and2 I293_021(w_293_021, w_037_101, w_131_007);
  or2  I293_033(w_293_033, w_191_232, w_061_147);
  or2  I293_036(w_293_036, w_202_153, w_077_552);
  or2  I293_038(w_293_038, w_015_091, w_165_056);
  nand2 I293_067(w_293_067, w_283_038, w_253_221);
  not1 I293_084(w_293_084, w_214_010);
  or2  I293_101(w_293_101, w_181_132, w_269_122);
  not1 I293_149(w_293_149, w_052_021);
  not1 I293_208(w_293_208, w_052_021);
  and2 I293_225(w_293_225, w_146_324, w_055_161);
  not1 I293_226(w_293_226, w_263_062);
  nand2 I293_325(w_293_325, w_150_334, w_160_611);
  not1 I293_359(w_293_359, w_242_162);
  not1 I293_386(w_293_386, w_182_010);
  or2  I294_000(w_294_000, w_109_240, w_149_159);
  nand2 I294_009(w_294_009, w_202_064, w_207_202);
  and2 I294_017(w_294_017, w_101_056, w_066_234);
  not1 I294_019(w_294_019, w_143_044);
  and2 I294_031(w_294_031, w_196_016, w_226_222);
  and2 I294_037(w_294_037, w_173_026, w_174_104);
  nand2 I294_046(w_294_046, w_051_372, w_146_142);
  not1 I294_055(w_294_055, w_117_040);
  and2 I294_064(w_294_064, w_240_125, w_122_093);
  nand2 I294_070(w_294_070, w_229_035, w_249_340);
  nand2 I294_074(w_294_074, w_086_091, w_233_012);
  nand2 I294_083(w_294_083, w_062_704, w_269_382);
  nand2 I294_110(w_294_110, w_176_049, w_121_192);
  not1 I294_111(w_294_111, w_210_139);
  nand2 I294_118(w_294_118, w_098_031, w_223_151);
  not1 I294_145(w_294_145, w_132_262);
  and2 I294_148(w_294_148, w_126_164, w_167_057);
  nand2 I295_020(w_295_020, w_274_055, w_125_439);
  nand2 I295_092(w_295_092, w_217_049, w_076_327);
  not1 I295_112(w_295_112, w_184_038);
  or2  I295_122(w_295_122, w_120_648, w_023_128);
  and2 I295_173(w_295_173, w_009_316, w_091_008);
  not1 I295_188(w_295_188, w_021_122);
  and2 I295_227(w_295_227, w_121_057, w_096_003);
  or2  I295_247(w_295_247, w_215_286, w_077_431);
  and2 I295_275(w_295_275, w_266_307, w_216_234);
  or2  I295_280(w_295_280, w_198_006, w_031_043);
  nand2 I295_308(w_295_308, w_086_049, w_064_014);
  or2  I295_312(w_295_312, w_290_048, w_122_113);
  or2  I295_400(w_295_400, w_101_280, w_031_120);
  or2  I296_032(w_296_032, w_227_036, w_031_015);
  nand2 I296_041(w_296_041, w_214_577, w_124_256);
  nand2 I296_129(w_296_129, w_042_220, w_065_411);
  not1 I296_132(w_296_132, w_064_315);
  or2  I296_200(w_296_200, w_123_104, w_273_112);
  nand2 I296_302(w_296_302, w_140_068, w_030_041);
  nand2 I296_316(w_296_316, w_196_217, w_120_626);
  or2  I296_354(w_296_354, w_037_234, w_194_262);
  nand2 I297_054(w_297_054, w_095_034, w_191_229);
  and2 I297_116(w_297_116, w_053_025, w_275_598);
  and2 I298_000(w_298_000, w_069_145, w_048_004);
  or2  I298_003(w_298_003, w_097_393, w_274_170);
  or2  I298_019(w_298_019, w_125_036, w_202_252);
  not1 I298_031(w_298_031, w_130_294);
  and2 I298_035(w_298_035, w_122_091, w_001_030);
  nand2 I298_038(w_298_038, w_044_496, w_260_030);
  nand2 I298_057(w_298_057, w_060_012, w_230_266);
  not1 I298_073(w_298_073, w_086_253);
  or2  I298_087(w_298_087, w_033_062, w_165_094);
  not1 I298_090(w_298_090, w_113_347);
  not1 I298_091(w_298_091, w_160_056);
  not1 I298_099(w_298_099, w_185_104);
  or2  I298_100(w_298_100, w_278_060, w_073_196);
  and2 I299_015(w_299_015, w_278_057, w_161_035);
  and2 I299_020(w_299_020, w_224_405, w_109_209);
  not1 I299_050(w_299_050, w_150_241);
  nand2 I299_053(w_299_053, w_116_004, w_084_043);
  not1 I299_097(w_299_097, w_079_000);
  or2  I299_149(w_299_149, w_171_013, w_109_204);
  or2  I299_164(w_299_164, w_163_099, w_120_176);
  and2 I299_245(w_299_245, w_203_083, w_113_136);
  or2  I299_261(w_299_261, w_005_184, w_210_107);
  not1 I299_270(w_299_270, w_128_070);
  not1 I299_288(w_299_288, w_116_042);
  not1 I299_315(w_299_315, w_047_032);
  not1 I299_316(w_299_316, w_040_090);
  and2 I299_475(w_299_477, w_299_476, w_091_024);
  or2  I299_476(w_299_478, w_299_477, w_284_049);
  and2 I299_477(w_299_479, w_299_478, w_154_095);
  not1 I299_478(w_299_480, w_299_479);
  nand2 I299_479(w_299_481, w_299_494, w_299_480);
  not1 I299_480(w_299_482, w_299_481);
  not1 I299_481(w_299_483, w_299_482);
  not1 I299_482(w_299_484, w_299_483);
  not1 I299_483(w_299_485, w_299_484);
  and2 I299_484(w_299_486, w_159_008, w_299_485);
  and2 I299_485(w_299_476, w_258_449, w_299_486);
  or2  I299_486(w_299_491, w_299_490, w_109_177);
  and2 I299_487(w_299_492, w_299_491, w_105_091);
  not1 I299_488(w_299_490, w_299_481);
  and2 I299_489(w_299_494, w_153_026, w_299_492);
  and2 I300_010(w_300_010, w_174_024, w_039_602);
  and2 I300_046(w_300_046, w_003_078, w_213_179);
  and2 I300_064(w_300_064, w_188_003, w_154_131);
  or2  I300_085(w_300_085, w_158_000, w_235_056);
  and2 I300_111(w_300_111, w_142_607, w_005_208);
  and2 I300_139(w_300_139, w_134_140, w_055_091);
  not1 I300_176(w_300_176, w_243_143);
  not1 I300_261(w_300_261, w_143_082);
  and2 I300_425(w_300_425, w_179_579, w_156_261);
  not1 I300_610(w_300_610, w_008_020);
  nand2 I301_002(w_301_002, w_118_017, w_203_143);
  nand2 I301_014(w_301_014, w_045_331, w_233_386);
  or2  I301_027(w_301_027, w_162_001, w_133_000);
  or2  I301_046(w_301_046, w_047_140, w_216_105);
  or2  I301_062(w_301_062, w_033_638, w_196_072);
  and2 I301_066(w_301_066, w_195_003, w_224_256);
  nand2 I301_091(w_301_091, w_194_173, w_217_061);
  and2 I301_121(w_301_121, w_179_583, w_291_085);
  or2  I301_153(w_301_153, w_097_373, w_299_245);
  or2  I301_182(w_301_182, w_034_035, w_284_039);
  nand2 I301_197(w_301_197, w_150_274, w_208_035);
  or2  I301_210(w_301_210, w_294_111, w_298_035);
  or2  I301_220(w_301_220, w_009_110, w_187_039);
  and2 I302_049(w_302_049, w_165_150, w_238_021);
  and2 I302_076(w_302_076, w_269_070, w_181_147);
  or2  I302_117(w_302_117, w_238_010, w_061_305);
  not1 I302_261(w_302_261, w_213_600);
  or2  I302_338(w_302_338, w_124_295, w_173_003);
  nand2 I302_495(w_302_495, w_044_373, w_074_370);
  not1 I302_529(w_302_529, w_271_602);
  nand2 I302_629(w_302_629, w_263_133, w_018_010);
  nand2 I303_059(w_303_059, w_148_286, w_248_142);
  and2 I303_070(w_303_070, w_268_079, w_299_149);
  or2  I303_078(w_303_078, w_213_005, w_230_095);
  and2 I303_080(w_303_080, w_164_374, w_225_086);
  nand2 I303_095(w_303_095, w_289_121, w_250_288);
  or2  I303_100(w_303_100, w_296_316, w_212_170);
  and2 I303_106(w_303_106, w_288_422, w_293_038);
  not1 I303_119(w_303_119, w_272_026);
  or2  I303_121(w_303_121, w_165_054, w_260_161);
  not1 I303_128(w_303_128, w_288_288);
  or2  I304_003(w_304_003, w_204_386, w_283_138);
  nand2 I304_022(w_304_022, w_144_105, w_279_068);
  not1 I304_079(w_304_079, w_057_257);
  or2  I304_083(w_304_083, w_016_006, w_237_063);
  and2 I304_100(w_304_100, w_109_358, w_140_052);
  nand2 I304_178(w_304_178, w_043_023, w_287_180);
  and2 I304_192(w_304_192, w_089_118, w_047_118);
  not1 I304_223(w_304_223, w_036_096);
  not1 I304_258(w_304_258, w_071_084);
  nand2 I304_315(w_304_315, w_036_242, w_027_191);
  nand2 I304_331(w_304_331, w_117_045, w_112_127);
  nand2 I304_414(w_304_414, w_044_689, w_116_500);
  nand2 I304_437(w_304_437, w_112_079, w_200_498);
  or2  I304_443(w_304_443, w_078_251, w_236_046);
  nand2 I304_468(w_304_468, w_003_001, w_058_420);
  or2  I304_500(w_304_500, w_161_365, w_213_541);
  nand2 I305_057(w_305_057, w_081_012, w_023_064);
  nand2 I305_077(w_305_077, w_282_110, w_076_091);
  or2  I305_083(w_305_083, w_242_132, w_132_390);
  not1 I305_103(w_305_103, w_109_358);
  or2  I305_157(w_305_157, w_218_698, w_071_304);
  not1 I305_178(w_305_178, w_069_159);
  or2  I305_188(w_305_188, w_055_006, w_084_047);
  not1 I305_239(w_305_239, w_166_199);
  not1 I305_270(w_305_270, w_257_293);
  and2 I305_471(w_305_471, w_145_068, w_116_387);
  not1 I305_536(w_305_536, w_125_065);
  not1 I306_018(w_306_018, w_039_510);
  nand2 I306_041(w_306_041, w_074_294, w_149_080);
  not1 I306_087(w_306_087, w_020_153);
  not1 I306_106(w_306_106, w_198_057);
  or2  I306_112(w_306_112, w_147_027, w_050_367);
  and2 I306_146(w_306_146, w_271_354, w_003_067);
  or2  I306_151(w_306_151, w_144_043, w_210_014);
  nand2 I306_165(w_306_165, w_272_021, w_010_162);
  and2 I306_177(w_306_177, w_130_463, w_088_016);
  not1 I306_207(w_306_207, w_104_073);
  and2 I306_236(w_306_236, w_099_131, w_158_000);
  or2  I306_272(w_306_272, w_227_647, w_226_171);
  and2 I306_281(w_306_281, w_180_023, w_065_026);
  not1 I307_036(w_307_036, w_008_036);
  and2 I307_040(w_307_040, w_247_162, w_164_119);
  not1 I307_043(w_307_043, w_159_032);
  or2  I307_075(w_307_075, w_220_322, w_245_153);
  not1 I307_081(w_307_081, w_224_494);
  or2  I307_093(w_307_093, w_156_130, w_023_016);
  and2 I307_095(w_307_095, w_000_663, w_173_012);
  not1 I307_123(w_307_123, w_247_154);
  and2 I307_166(w_307_166, w_137_223, w_259_224);
  nand2 I307_305(w_307_305, w_214_181, w_271_637);
  not1 I307_343(w_307_343, w_112_019);
  or2  I307_350(w_307_350, w_279_127, w_069_023);
  nand2 I307_391(w_307_391, w_035_036, w_060_119);
  nand2 I307_415(w_307_415, w_260_151, w_021_184);
  and2 I308_008(w_308_008, w_258_247, w_164_127);
  and2 I308_022(w_308_022, w_278_174, w_068_083);
  not1 I308_026(w_308_026, w_289_417);
  or2  I308_034(w_308_034, w_288_278, w_174_075);
  or2  I308_064(w_308_064, w_095_040, w_044_454);
  not1 I308_067(w_308_067, w_138_134);
  not1 I308_095(w_308_095, w_070_007);
  not1 I308_107(w_308_107, w_019_020);
  or2  I308_115(w_308_115, w_090_528, w_231_064);
  and2 I308_123(w_308_123, w_131_109, w_065_474);
  not1 I308_126(w_308_126, w_210_028);
  not1 I308_146(w_308_146, w_234_182);
  or2  I308_147(w_308_147, w_246_573, w_025_231);
  nand2 I308_155(w_308_155, w_194_117, w_012_106);
  nand2 I309_034(w_309_034, w_078_121, w_250_513);
  nand2 I309_187(w_309_187, w_222_521, w_061_388);
  nand2 I309_193(w_309_193, w_034_003, w_281_212);
  not1 I309_215(w_309_215, w_127_011);
  or2  I309_264(w_309_264, w_136_037, w_075_147);
  nand2 I309_270(w_309_270, w_118_080, w_044_054);
  not1 I309_301(w_309_301, w_132_179);
  not1 I309_352(w_309_352, w_225_240);
  not1 I309_380(w_309_380, w_241_032);
  and2 I309_381(w_309_383, w_309_382, w_069_144);
  and2 I309_382(w_309_384, w_242_133, w_309_383);
  nand2 I309_383(w_309_385, w_081_012, w_309_384);
  and2 I309_384(w_309_386, w_309_385, w_048_010);
  not1 I309_385(w_309_387, w_309_386);
  nand2 I309_386(w_309_388, w_309_387, w_222_226);
  and2 I309_387(w_309_389, w_309_388, w_200_436);
  or2  I309_388(w_309_390, w_309_389, w_217_034);
  and2 I309_389(w_309_391, w_309_390, w_046_299);
  or2  I309_390(w_309_382, w_226_077, w_309_391);
  nand2 I310_061(w_310_061, w_248_142, w_219_413);
  not1 I310_071(w_310_071, w_309_301);
  or2  I310_093(w_310_093, w_144_173, w_153_037);
  and2 I310_145(w_310_145, w_128_195, w_007_197);
  and2 I310_165(w_310_165, w_277_137, w_055_137);
  and2 I310_188(w_310_188, w_075_002, w_300_111);
  not1 I310_244(w_310_244, w_192_164);
  and2 I310_251(w_310_251, w_025_056, w_294_055);
  nand2 I310_258(w_310_258, w_052_025, w_071_247);
  and2 I310_365(w_310_365, w_228_374, w_254_084);
  and2 I310_412(w_310_412, w_202_085, w_248_042);
  not1 I310_447(w_310_447, w_251_017);
  not1 I310_496(w_310_496, w_072_187);
  or2  I310_557(w_310_557, w_040_594, w_272_043);
  and2 I310_582(w_310_582, w_123_592, w_171_265);
  not1 I311_003(w_311_003, w_057_084);
  not1 I311_080(w_311_080, w_063_004);
  or2  I311_123(w_311_123, w_230_077, w_070_084);
  and2 I311_131(w_311_131, w_192_113, w_307_075);
  and2 I311_134(w_311_134, w_229_285, w_172_033);
  nand2 I311_180(w_311_180, w_233_088, w_126_128);
  or2  I311_245(w_311_245, w_179_159, w_158_002);
  or2  I311_256(w_311_256, w_237_012, w_291_063);
  or2  I311_263(w_311_263, w_204_323, w_234_403);
  or2  I311_288(w_311_288, w_167_152, w_189_484);
  and2 I311_325(w_311_325, w_119_139, w_118_040);
  or2  I311_369(w_311_369, w_304_003, w_215_346);
  or2  I311_439(w_311_439, w_195_177, w_248_028);
  or2  I312_023(w_312_023, w_211_027, w_170_277);
  nand2 I312_040(w_312_040, w_293_208, w_196_095);
  nand2 I312_042(w_312_042, w_097_056, w_100_037);
  nand2 I312_056(w_312_056, w_241_021, w_193_137);
  nand2 I312_060(w_312_060, w_115_008, w_247_161);
  not1 I312_133(w_312_133, w_133_057);
  and2 I312_146(w_312_146, w_271_011, w_100_130);
  nand2 I312_238(w_312_238, w_245_730, w_273_105);
  or2  I312_355(w_312_355, w_003_025, w_049_288);
  and2 I312_363(w_312_363, w_156_029, w_074_153);
  nand2 I312_432(w_312_432, w_127_034, w_018_020);
  and2 I313_008(w_313_008, w_114_009, w_200_021);
  nand2 I313_030(w_313_030, w_059_423, w_143_090);
  and2 I313_080(w_313_080, w_218_178, w_199_076);
  and2 I313_083(w_313_083, w_066_134, w_301_062);
  not1 I313_090(w_313_090, w_192_134);
  and2 I313_118(w_313_118, w_033_241, w_202_196);
  not1 I313_128(w_313_128, w_174_092);
  or2  I313_149(w_313_149, w_264_666, w_046_068);
  nand2 I313_192(w_313_192, w_276_331, w_081_016);
  nand2 I313_231(w_313_231, w_200_045, w_041_453);
  nand2 I313_240(w_313_240, w_186_099, w_267_041);
  or2  I313_254(w_313_254, w_081_011, w_059_003);
  and2 I313_258(w_313_258, w_305_157, w_118_067);
  or2  I313_397(w_313_397, w_052_037, w_287_064);
  not1 I313_403(w_313_403, w_169_279);
  and2 I314_014(w_314_014, w_139_005, w_070_476);
  not1 I314_032(w_314_032, w_082_505);
  or2  I314_077(w_314_077, w_230_080, w_164_294);
  and2 I314_092(w_314_092, w_063_527, w_022_268);
  not1 I314_134(w_314_134, w_304_022);
  or2  I314_159(w_314_159, w_128_559, w_213_052);
  and2 I314_174(w_314_174, w_085_176, w_191_062);
  nand2 I314_191(w_314_191, w_268_268, w_059_055);
  or2  I314_204(w_314_204, w_076_311, w_072_116);
  and2 I314_218(w_314_220, w_314_219, w_086_059);
  and2 I314_219(w_314_221, w_314_220, w_314_234);
  nand2 I314_220(w_314_219, w_314_221, w_073_404);
  and2 I314_221(w_314_226, w_098_057, w_314_225);
  nand2 I314_222(w_314_227, w_314_226, w_246_307);
  nand2 I314_223(w_314_228, w_314_227, w_157_074);
  not1 I314_224(w_314_229, w_314_228);
  not1 I314_225(w_314_230, w_314_229);
  not1 I314_226(w_314_231, w_314_230);
  and2 I314_227(w_314_232, w_035_043, w_314_231);
  not1 I314_228(w_314_225, w_314_221);
  and2 I314_229(w_314_234, w_252_363, w_314_232);
  or2  I315_111(w_315_111, w_256_689, w_198_021);
  or2  I315_140(w_315_140, w_077_102, w_300_425);
  not1 I315_171(w_315_171, w_042_124);
  not1 I315_238(w_315_238, w_211_017);
  not1 I315_269(w_315_269, w_285_774);
  not1 I315_362(w_315_362, w_284_024);
  not1 I315_523(w_315_523, w_239_000);
  or2  I315_524(w_315_524, w_287_369, w_277_123);
  and2 I315_530(w_315_530, w_208_225, w_191_245);
  and2 I315_634(w_315_634, w_070_014, w_104_067);
  nand2 I315_665(w_315_665, w_220_350, w_116_343);
  nand2 I315_724(w_315_724, w_104_157, w_022_210);
  not1 I316_066(w_316_066, w_143_535);
  or2  I316_072(w_316_072, w_032_108, w_115_066);
  not1 I316_149(w_316_149, w_076_183);
  not1 I316_219(w_316_219, w_148_375);
  not1 I316_246(w_316_246, w_021_071);
  or2  I316_257(w_316_257, w_121_202, w_247_135);
  or2  I316_410(w_316_410, w_266_247, w_028_053);
  and2 I316_450(w_316_450, w_308_126, w_163_343);
  nand2 I316_453(w_316_453, w_005_065, w_276_170);
  nand2 I317_014(w_317_014, w_177_108, w_268_021);
  and2 I317_090(w_317_090, w_074_030, w_052_036);
  and2 I317_148(w_317_148, w_183_011, w_194_221);
  or2  I317_162(w_317_162, w_038_225, w_228_005);
  nand2 I317_249(w_317_249, w_113_237, w_204_135);
  and2 I317_261(w_317_261, w_152_513, w_233_239);
  and2 I317_264(w_317_264, w_272_018, w_107_219);
  nand2 I317_298(w_317_298, w_160_394, w_250_252);
  or2  I318_000(w_318_000, w_195_107, w_100_008);
  not1 I318_003(w_318_003, w_151_352);
  or2  I318_004(w_318_004, w_276_200, w_015_115);
  nand2 I318_011(w_318_011, w_279_069, w_187_002);
  nand2 I318_012(w_318_012, w_170_331, w_210_107);
  not1 I318_013(w_318_013, w_140_071);
  nand2 I318_014(w_318_014, w_192_009, w_184_130);
  nand2 I318_015(w_318_015, w_014_075, w_033_161);
  not1 I319_077(w_319_077, w_227_231);
  or2  I319_129(w_319_129, w_169_170, w_156_289);
  not1 I319_200(w_319_200, w_014_054);
  nand2 I319_210(w_319_210, w_032_168, w_181_195);
  nand2 I319_218(w_319_218, w_191_011, w_220_231);
  not1 I319_278(w_319_278, w_246_286);
  or2  I319_289(w_319_289, w_194_057, w_113_032);
  or2  I319_347(w_319_347, w_018_030, w_102_337);
  nand2 I320_004(w_320_004, w_008_490, w_053_055);
  and2 I320_019(w_320_019, w_273_042, w_062_377);
  not1 I320_123(w_320_123, w_118_090);
  not1 I320_178(w_320_178, w_121_055);
  or2  I320_218(w_320_218, w_053_051, w_054_009);
  nand2 I320_224(w_320_224, w_107_056, w_293_386);
  or2  I320_285(w_320_285, w_033_309, w_282_137);
  and2 I320_297(w_320_297, w_146_321, w_037_048);
  not1 I320_309(w_320_309, w_184_049);
  or2  I320_318(w_320_318, w_145_016, w_117_051);
  not1 I320_369(w_320_369, w_170_139);
  nand2 I320_389(w_320_389, w_003_063, w_206_047);
  and2 I320_411(w_320_411, w_289_103, w_128_181);
  nand2 I321_001(w_321_001, w_042_133, w_155_109);
  nand2 I321_005(w_321_005, w_156_472, w_315_530);
  nand2 I321_063(w_321_063, w_243_109, w_103_301);
  and2 I321_141(w_321_141, w_239_000, w_058_559);
  and2 I321_176(w_321_176, w_181_265, w_272_028);
  nand2 I321_282(w_321_282, w_092_481, w_125_128);
  nand2 I321_303(w_321_303, w_026_294, w_284_102);
  nand2 I321_536(w_321_536, w_241_055, w_293_225);
  not1 I322_001(w_322_001, w_244_238);
  or2  I322_002(w_322_002, w_103_220, w_098_034);
  not1 I322_005(w_322_005, w_216_376);
  nand2 I322_008(w_322_008, w_162_015, w_009_337);
  or2  I322_013(w_322_013, w_126_104, w_208_072);
  nand2 I322_014(w_322_014, w_184_025, w_040_053);
  or2  I322_015(w_322_015, w_089_134, w_106_037);
  or2  I322_017(w_322_017, w_161_533, w_082_431);
  or2  I322_022(w_322_022, w_025_035, w_247_076);
  nand2 I323_061(w_323_061, w_223_241, w_252_012);
  nand2 I323_089(w_323_089, w_305_536, w_137_116);
  nand2 I323_123(w_323_123, w_133_120, w_199_373);
  not1 I323_139(w_323_139, w_223_218);
  not1 I323_230(w_323_230, w_035_124);
  not1 I323_269(w_323_269, w_264_157);
  and2 I323_284(w_323_284, w_296_354, w_023_091);
  nand2 I324_008(w_324_008, w_292_533, w_228_050);
  and2 I324_011(w_324_011, w_257_054, w_196_075);
  not1 I324_012(w_324_012, w_097_430);
  or2  I324_029(w_324_029, w_209_145, w_022_173);
  and2 I324_031(w_324_031, w_220_346, w_212_048);
  not1 I324_035(w_324_035, w_284_080);
  or2  I324_045(w_324_045, w_246_014, w_053_000);
  and2 I324_052(w_324_052, w_158_003, w_025_063);
  or2  I325_000(w_325_000, w_072_157, w_293_036);
  nand2 I325_005(w_325_005, w_295_400, w_058_174);
  and2 I325_035(w_325_035, w_081_010, w_195_084);
  not1 I325_046(w_325_046, w_315_665);
  nand2 I325_139(w_325_139, w_244_117, w_153_019);
  or2  I325_238(w_325_238, w_176_097, w_324_052);
  not1 I325_272(w_325_272, w_043_047);
  and2 I325_310(w_325_310, w_241_031, w_066_095);
  and2 I326_031(w_326_031, w_034_008, w_157_160);
  nand2 I326_035(w_326_035, w_305_239, w_321_001);
  and2 I326_042(w_326_042, w_142_321, w_098_059);
  and2 I326_043(w_326_043, w_275_133, w_013_224);
  not1 I326_077(w_326_077, w_110_294);
  nand2 I326_104(w_326_104, w_227_026, w_139_014);
  nand2 I326_111(w_326_111, w_233_168, w_236_097);
  not1 I326_113(w_326_113, w_038_606);
  nand2 I326_114(w_326_114, w_002_645, w_241_085);
  or2  I326_179(w_326_179, w_046_447, w_277_013);
  nand2 I327_097(w_327_097, w_057_047, w_200_234);
  or2  I327_155(w_327_155, w_087_228, w_160_479);
  and2 I327_344(w_327_344, w_184_011, w_285_393);
  nand2 I327_363(w_327_363, w_212_019, w_081_010);
  and2 I327_364(w_327_364, w_047_443, w_199_240);
  nand2 I327_438(w_327_438, w_305_188, w_042_171);
  and2 I327_440(w_327_440, w_141_117, w_253_023);
  and2 I327_444(w_327_444, w_193_345, w_120_684);
  nand2 I328_004(w_328_004, w_138_205, w_063_110);
  and2 I328_010(w_328_010, w_320_123, w_195_023);
  nand2 I328_026(w_328_026, w_119_106, w_087_168);
  and2 I328_037(w_328_037, w_058_423, w_099_059);
  nand2 I328_053(w_328_053, w_288_087, w_188_091);
  and2 I328_110(w_328_110, w_245_188, w_147_037);
  or2  I328_120(w_328_120, w_110_262, w_132_249);
  not1 I328_153(w_328_153, w_243_111);
  or2  I329_037(w_329_037, w_014_229, w_262_068);
  nand2 I329_039(w_329_039, w_298_091, w_196_007);
  not1 I329_094(w_329_094, w_083_113);
  not1 I329_306(w_329_306, w_121_051);
  and2 I329_384(w_329_384, w_001_017, w_279_068);
  nand2 I330_016(w_330_016, w_160_039, w_249_152);
  nand2 I330_035(w_330_035, w_151_160, w_328_010);
  or2  I330_042(w_330_042, w_216_357, w_235_114);
  and2 I330_059(w_330_059, w_195_035, w_269_414);
  not1 I330_116(w_330_116, w_291_082);
  not1 I330_201(w_330_201, w_035_056);
  nand2 I330_247(w_330_247, w_138_238, w_111_106);
  nand2 I330_279(w_330_279, w_215_438, w_088_032);
  not1 I331_025(w_331_025, w_260_035);
  and2 I331_052(w_331_052, w_252_065, w_173_008);
  nand2 I331_072(w_331_072, w_186_537, w_023_019);
  nand2 I331_111(w_331_111, w_300_176, w_259_506);
  or2  I331_153(w_331_153, w_062_544, w_057_087);
  or2  I331_247(w_331_247, w_218_261, w_231_160);
  nand2 I331_255(w_331_255, w_284_081, w_125_354);
  and2 I331_315(w_331_315, w_274_232, w_243_015);
  or2  I331_330(w_331_330, w_090_272, w_244_053);
  or2  I331_439(w_331_439, w_125_282, w_245_339);
  nand2 I331_506(w_331_508, w_170_053, w_331_507);
  or2  I331_507(w_331_509, w_331_508, w_331_527);
  nand2 I331_508(w_331_510, w_128_353, w_331_509);
  nand2 I331_509(w_331_511, w_089_198, w_331_510);
  not1 I331_510(w_331_512, w_331_511);
  not1 I331_511(w_331_513, w_331_512);
  not1 I331_512(w_331_514, w_331_513);
  and2 I331_513(w_331_515, w_331_514, w_026_579);
  not1 I331_514(w_331_507, w_331_515);
  nand2 I331_515(w_331_520, w_331_519, w_039_616);
  or2  I331_516(w_331_521, w_331_520, w_102_561);
  or2  I331_517(w_331_522, w_149_430, w_331_521);
  and2 I331_518(w_331_523, w_030_056, w_331_522);
  or2  I331_519(w_331_524, w_331_523, w_189_119);
  and2 I331_520(w_331_525, w_331_524, w_175_477);
  not1 I331_521(w_331_519, w_331_509);
  and2 I331_522(w_331_527, w_147_166, w_331_525);
  not1 I332_004(w_332_004, w_054_074);
  and2 I332_142(w_332_142, w_102_035, w_329_037);
  and2 I332_224(w_332_224, w_190_095, w_096_000);
  nand2 I332_261(w_332_261, w_204_651, w_048_001);
  or2  I332_363(w_332_363, w_147_173, w_184_056);
  or2  I332_409(w_332_409, w_142_777, w_304_443);
  not1 I332_451(w_332_451, w_020_027);
  and2 I332_667(w_332_669, w_332_668, w_069_068);
  or2  I332_668(w_332_670, w_332_669, w_113_019);
  or2  I332_669(w_332_671, w_332_670, w_300_046);
  not1 I332_670(w_332_672, w_332_671);
  or2  I332_671(w_332_673, w_332_672, w_003_046);
  and2 I332_672(w_332_674, w_332_673, w_050_127);
  and2 I332_673(w_332_675, w_094_564, w_332_674);
  not1 I332_674(w_332_668, w_332_675);
  nand2 I333_011(w_333_011, w_019_017, w_316_072);
  not1 I333_115(w_333_115, w_311_131);
  or2  I333_137(w_333_137, w_094_057, w_138_168);
  nand2 I333_158(w_333_158, w_121_161, w_024_206);
  not1 I333_222(w_333_222, w_001_014);
  nand2 I333_223(w_333_223, w_320_369, w_087_379);
  nand2 I333_314(w_333_314, w_057_273, w_003_066);
  nand2 I334_098(w_334_098, w_250_609, w_075_027);
  nand2 I334_139(w_334_139, w_084_023, w_162_000);
  and2 I334_337(w_334_337, w_033_014, w_207_050);
  or2  I334_340(w_334_340, w_011_568, w_259_543);
  not1 I334_367(w_334_367, w_097_004);
  nand2 I334_368(w_334_368, w_144_186, w_007_234);
  not1 I334_486(w_334_486, w_302_117);
  and2 I334_640(w_334_640, w_205_173, w_240_114);
  not1 I335_033(w_335_033, w_290_103);
  and2 I335_041(w_335_041, w_167_014, w_182_015);
  or2  I335_098(w_335_098, w_207_233, w_177_402);
  nand2 I335_102(w_335_102, w_105_088, w_331_330);
  nand2 I335_116(w_335_116, w_083_170, w_205_330);
  or2  I335_134(w_335_134, w_128_291, w_077_540);
  or2  I335_151(w_335_151, w_043_003, w_260_101);
  and2 I335_162(w_335_162, w_145_070, w_240_019);
  nand2 I336_002(w_336_002, w_191_026, w_095_031);
  or2  I336_016(w_336_016, w_153_085, w_292_309);
  or2  I336_025(w_336_025, w_104_323, w_032_510);
  and2 I336_029(w_336_029, w_248_025, w_197_160);
  or2  I336_057(w_336_057, w_060_168, w_009_600);
  and2 I336_074(w_336_074, w_216_253, w_029_099);
  not1 I336_083(w_336_083, w_287_335);
  not1 I336_110(w_336_110, w_001_023);
  nand2 I336_124(w_336_124, w_061_058, w_257_143);
  and2 I336_140(w_336_140, w_298_031, w_151_208);
  not1 I336_177(w_336_177, w_281_237);
  and2 I336_209(w_336_209, w_063_438, w_093_208);
  or2  I336_235(w_336_235, w_070_033, w_003_060);
  or2  I337_004(w_337_004, w_054_262, w_236_010);
  nand2 I337_020(w_337_020, w_299_020, w_156_150);
  or2  I337_028(w_337_028, w_062_116, w_273_092);
  not1 I337_036(w_337_036, w_290_086);
  or2  I337_072(w_337_072, w_155_415, w_264_266);
  or2  I337_101(w_337_101, w_229_000, w_157_126);
  and2 I337_188(w_337_188, w_228_011, w_212_182);
  or2  I337_225(w_337_225, w_243_181, w_104_326);
  or2  I337_356(w_337_356, w_123_013, w_160_382);
  not1 I337_384(w_337_384, w_231_199);
  and2 I337_412(w_337_412, w_244_216, w_093_186);
  nand2 I338_003(w_338_003, w_041_248, w_246_521);
  nand2 I338_010(w_338_010, w_064_061, w_306_018);
  or2  I338_022(w_338_022, w_016_000, w_330_035);
  and2 I338_028(w_338_028, w_118_018, w_311_180);
  and2 I338_044(w_338_044, w_122_102, w_067_169);
  or2  I338_049(w_338_049, w_032_068, w_099_055);
  and2 I338_094(w_338_094, w_230_298, w_313_149);
  and2 I338_158(w_338_158, w_006_163, w_146_079);
  nand2 I338_239(w_338_239, w_267_083, w_125_081);
  and2 I338_264(w_338_264, w_314_134, w_123_029);
  or2  I338_312(w_338_312, w_105_226, w_037_050);
  and2 I339_003(w_339_003, w_192_146, w_090_042);
  and2 I339_008(w_339_008, w_062_349, w_032_520);
  not1 I339_012(w_339_012, w_267_114);
  nand2 I339_019(w_339_019, w_077_315, w_258_032);
  or2  I339_020(w_339_020, w_055_241, w_246_485);
  nand2 I339_022(w_339_022, w_063_252, w_153_055);
  not1 I339_028(w_339_028, w_044_109);
  or2  I339_029(w_339_029, w_107_288, w_269_405);
  not1 I339_039(w_339_039, w_072_111);
  or2  I339_041(w_339_041, w_284_129, w_206_145);
  and2 I340_000(w_340_000, w_092_272, w_154_031);
  or2  I340_004(w_340_004, w_331_439, w_234_254);
  not1 I340_010(w_340_010, w_215_344);
  and2 I340_011(w_340_011, w_079_015, w_294_055);
  and2 I340_013(w_340_013, w_194_178, w_070_220);
  not1 I340_026(w_340_026, w_158_004);
  nand2 I340_030(w_340_030, w_245_624, w_024_016);
  nand2 I340_038(w_340_038, w_164_588, w_004_151);
  or2  I340_046(w_340_046, w_266_124, w_295_280);
  not1 I340_048(w_340_050, w_340_049);
  not1 I340_049(w_340_051, w_340_050);
  and2 I340_050(w_340_052, w_089_197, w_340_051);
  and2 I340_051(w_340_053, w_051_037, w_340_052);
  or2  I340_052(w_340_054, w_216_002, w_340_053);
  nand2 I340_053(w_340_055, w_340_054, w_097_118);
  or2  I340_054(w_340_056, w_107_310, w_340_055);
  not1 I340_055(w_340_057, w_340_056);
  and2 I340_056(w_340_058, w_340_057, w_305_471);
  not1 I340_057(w_340_049, w_340_058);
  not1 I341_035(w_341_035, w_045_277);
  nand2 I341_245(w_341_245, w_216_308, w_320_285);
  and2 I341_351(w_341_351, w_016_005, w_187_019);
  not1 I341_408(w_341_408, w_163_327);
  and2 I341_418(w_341_418, w_235_121, w_222_469);
  and2 I341_458(w_341_458, w_338_094, w_256_021);
  not1 I341_487(w_341_487, w_047_232);
  not1 I341_599(w_341_599, w_306_165);
  or2  I341_704(w_341_704, w_326_104, w_234_309);
  and2 I341_774(w_341_774, w_251_048, w_182_009);
  not1 I342_047(w_342_047, w_307_081);
  nand2 I342_103(w_342_103, w_167_140, w_092_307);
  not1 I342_111(w_342_111, w_285_353);
  or2  I342_194(w_342_194, w_184_056, w_050_437);
  nand2 I342_213(w_342_213, w_257_112, w_156_013);
  nand2 I342_217(w_342_217, w_078_024, w_112_140);
  nand2 I342_311(w_342_311, w_070_496, w_134_156);
  not1 I342_344(w_342_344, w_008_595);
  and2 I342_358(w_342_358, w_139_007, w_295_112);
  nand2 I342_477(w_342_477, w_212_190, w_027_011);
  nand2 I343_138(w_343_138, w_209_182, w_306_151);
  and2 I343_246(w_343_246, w_195_194, w_253_415);
  or2  I343_251(w_343_251, w_104_221, w_335_116);
  or2  I343_335(w_343_335, w_039_016, w_298_087);
  or2  I343_360(w_343_360, w_181_064, w_002_062);
  or2  I343_425(w_343_425, w_267_085, w_280_259);
  not1 I343_478(w_343_478, w_248_136);
  not1 I343_479(w_343_479, w_160_223);
  nand2 I343_580(w_343_580, w_018_000, w_083_009);
  and2 I343_605(w_343_605, w_242_000, w_129_186);
  or2  I343_697(w_343_697, w_122_032, w_131_430);
  and2 I344_001(w_344_001, w_104_362, w_022_319);
  and2 I344_026(w_344_026, w_320_224, w_262_202);
  nand2 I344_042(w_344_042, w_062_164, w_008_566);
  or2  I344_061(w_344_061, w_233_038, w_182_010);
  and2 I344_063(w_344_063, w_098_046, w_306_112);
  not1 I344_077(w_344_077, w_078_345);
  not1 I344_088(w_344_088, w_321_176);
  not1 I344_116(w_344_116, w_194_187);
  not1 I344_148(w_344_148, w_099_180);
  not1 I344_263(w_344_263, w_303_119);
  and2 I344_455(w_344_455, w_003_056, w_007_304);
  and2 I345_013(w_345_013, w_025_210, w_191_076);
  or2  I345_017(w_345_017, w_326_031, w_312_060);
  not1 I345_053(w_345_053, w_245_660);
  nand2 I345_098(w_345_098, w_267_183, w_088_132);
  not1 I345_129(w_345_129, w_080_279);
  nand2 I345_216(w_345_216, w_118_079, w_037_082);
  or2  I345_250(w_345_250, w_210_014, w_147_007);
  not1 I346_076(w_346_076, w_046_298);
  nand2 I346_104(w_346_104, w_020_453, w_007_126);
  and2 I346_139(w_346_139, w_119_016, w_254_031);
  nand2 I346_565(w_346_565, w_069_028, w_037_268);
  or2  I347_016(w_347_016, w_008_329, w_333_223);
  or2  I347_021(w_347_021, w_129_113, w_053_067);
  not1 I347_036(w_347_036, w_066_025);
  or2  I347_053(w_347_053, w_304_315, w_006_064);
  and2 I347_098(w_347_098, w_248_045, w_310_496);
  nand2 I347_109(w_347_109, w_087_425, w_217_014);
  nand2 I347_117(w_347_117, w_142_147, w_186_205);
  nand2 I347_167(w_347_167, w_335_041, w_343_360);
  and2 I347_252(w_347_252, w_012_095, w_034_064);
  and2 I347_257(w_347_257, w_103_064, w_260_166);
  nand2 I347_268(w_347_268, w_192_063, w_032_180);
  not1 I347_328(w_347_328, w_058_472);
  and2 I347_331(w_347_331, w_313_083, w_056_501);
  not1 I348_101(w_348_101, w_049_025);
  or2  I348_114(w_348_114, w_210_093, w_000_506);
  nand2 I348_137(w_348_137, w_154_097, w_102_144);
  not1 I348_213(w_348_213, w_328_026);
  and2 I348_243(w_348_243, w_225_168, w_306_272);
  not1 I349_027(w_349_027, w_311_245);
  not1 I349_028(w_349_028, w_284_014);
  or2  I349_036(w_349_036, w_003_002, w_183_041);
  nand2 I349_060(w_349_060, w_222_163, w_233_249);
  not1 I349_089(w_349_089, w_094_051);
  not1 I349_177(w_349_177, w_114_181);
  and2 I349_214(w_349_214, w_175_373, w_139_015);
  or2  I349_230(w_349_230, w_138_104, w_042_312);
  nand2 I349_289(w_349_289, w_195_241, w_247_131);
  and2 I349_305(w_349_305, w_282_206, w_199_159);
  not1 I350_022(w_350_022, w_190_116);
  not1 I350_049(w_350_049, w_290_004);
  not1 I350_071(w_350_071, w_002_067);
  not1 I350_094(w_350_094, w_116_424);
  and2 I350_123(w_350_123, w_016_002, w_019_007);
  and2 I351_044(w_351_044, w_153_025, w_117_022);
  and2 I351_049(w_351_049, w_212_009, w_116_140);
  not1 I351_051(w_351_051, w_281_643);
  and2 I351_070(w_351_070, w_038_074, w_255_081);
  or2  I351_075(w_351_075, w_260_199, w_223_166);
  and2 I351_095(w_351_095, w_116_136, w_344_263);
  and2 I351_106(w_351_106, w_328_004, w_308_026);
  not1 I351_228(w_351_228, w_209_209);
  nand2 I351_235(w_351_235, w_280_559, w_063_504);
  or2  I351_240(w_351_240, w_101_050, w_007_436);
  not1 I351_336(w_351_336, w_197_248);
  not1 I352_047(w_352_047, w_313_030);
  and2 I352_296(w_352_296, w_202_055, w_193_033);
  or2  I352_314(w_352_314, w_225_053, w_335_102);
  nand2 I352_411(w_352_411, w_279_153, w_052_020);
  and2 I353_047(w_353_047, w_026_237, w_276_142);
  nand2 I353_106(w_353_106, w_251_097, w_337_188);
  nand2 I353_137(w_353_137, w_251_075, w_167_152);
  or2  I353_189(w_353_189, w_245_696, w_141_171);
  or2  I353_244(w_353_244, w_331_255, w_285_689);
  and2 I353_311(w_353_311, w_202_095, w_166_110);
  or2  I353_443(w_353_443, w_300_064, w_346_139);
  or2  I353_535(w_353_535, w_221_044, w_223_040);
  nand2 I353_570(w_353_570, w_016_005, w_251_131);
  nand2 I354_003(w_354_003, w_148_241, w_254_020);
  or2  I354_004(w_354_004, w_245_448, w_001_019);
  or2  I354_010(w_354_010, w_094_574, w_086_164);
  not1 I354_039(w_354_039, w_085_158);
  and2 I354_048(w_354_048, w_209_012, w_128_306);
  not1 I354_082(w_354_082, w_252_272);
  nand2 I354_112(w_354_112, w_347_098, w_023_088);
  nand2 I354_113(w_354_113, w_150_345, w_283_329);
  and2 I354_207(w_354_207, w_100_100, w_349_036);
  and2 I355_038(w_355_038, w_276_030, w_147_162);
  and2 I355_051(w_355_051, w_259_469, w_190_100);
  or2  I355_071(w_355_071, w_310_188, w_213_241);
  not1 I355_072(w_355_072, w_299_050);
  or2  I355_079(w_355_079, w_026_250, w_196_149);
  or2  I355_100(w_355_100, w_209_062, w_056_463);
  or2  I355_113(w_355_113, w_107_400, w_152_573);
  nand2 I355_192(w_355_192, w_144_202, w_207_144);
  nand2 I355_295(w_355_295, w_282_291, w_107_021);
  not1 I355_297(w_355_297, w_180_024);
  and2 I355_405(w_355_405, w_107_293, w_277_067);
  and2 I356_001(w_356_001, w_340_046, w_001_028);
  and2 I356_003(w_356_003, w_062_384, w_291_073);
  or2  I356_039(w_356_039, w_209_345, w_316_453);
  or2  I356_043(w_356_043, w_087_058, w_098_014);
  and2 I356_044(w_356_044, w_086_029, w_078_511);
  nand2 I356_048(w_356_048, w_224_069, w_141_176);
  not1 I356_061(w_356_061, w_200_089);
  not1 I356_078(w_356_078, w_009_317);
  or2  I356_108(w_356_108, w_216_048, w_267_103);
  not1 I357_005(w_357_005, w_262_002);
  not1 I357_096(w_357_096, w_307_123);
  and2 I357_296(w_357_296, w_339_003, w_137_345);
  nand2 I357_302(w_357_302, w_002_349, w_109_251);
  nand2 I357_304(w_357_304, w_021_149, w_041_515);
  and2 I357_318(w_357_318, w_212_052, w_130_283);
  or2  I357_319(w_357_319, w_279_139, w_007_330);
  nand2 I357_381(w_357_381, w_278_100, w_202_014);
  or2  I357_408(w_357_408, w_311_134, w_004_275);
  and2 I357_460(w_357_460, w_214_148, w_131_431);
  and2 I357_588(w_357_588, w_112_120, w_033_783);
  or2  I357_658(w_357_658, w_063_084, w_197_017);
  nand2 I358_066(w_358_066, w_317_261, w_357_318);
  nand2 I358_227(w_358_227, w_283_216, w_055_155);
  nand2 I358_284(w_358_284, w_247_147, w_110_295);
  or2  I358_295(w_358_295, w_325_310, w_085_056);
  and2 I359_015(w_359_015, w_352_296, w_190_036);
  and2 I359_021(w_359_021, w_324_011, w_305_270);
  nand2 I359_041(w_359_041, w_233_101, w_164_302);
  and2 I359_047(w_359_047, w_254_058, w_214_021);
  nand2 I359_051(w_359_051, w_034_034, w_058_522);
  not1 I359_074(w_359_074, w_081_009);
  or2  I359_075(w_359_075, w_345_013, w_045_335);
  and2 I359_089(w_359_089, w_111_078, w_241_008);
  nand2 I359_090(w_359_090, w_304_331, w_243_297);
  nand2 I359_154(w_359_154, w_323_284, w_099_053);
  nand2 I359_170(w_359_170, w_204_493, w_016_002);
  and2 I359_176(w_359_176, w_116_426, w_027_140);
  not1 I359_198(w_359_198, w_071_056);
  and2 I359_208(w_359_210, w_359_209, w_009_146);
  or2  I359_209(w_359_211, w_359_210, w_229_046);
  not1 I359_210(w_359_212, w_359_211);
  not1 I359_211(w_359_213, w_359_212);
  not1 I359_212(w_359_214, w_359_213);
  not1 I359_213(w_359_215, w_359_214);
  nand2 I359_214(w_359_216, w_359_215, w_173_023);
  and2 I359_215(w_359_217, w_359_216, w_359_227);
  not1 I359_216(w_359_209, w_359_217);
  nand2 I359_217(w_359_222, w_349_089, w_359_221);
  nand2 I359_218(w_359_223, w_121_136, w_359_222);
  and2 I359_219(w_359_224, w_006_059, w_359_223);
  and2 I359_220(w_359_225, w_359_224, w_350_123);
  not1 I359_221(w_359_221, w_359_217);
  and2 I359_222(w_359_227, w_120_262, w_359_225);
  not1 I360_021(w_360_021, w_075_045);
  and2 I360_150(w_360_150, w_325_046, w_128_048);
  nand2 I360_266(w_360_266, w_159_029, w_302_076);
  and2 I360_269(w_360_269, w_200_128, w_109_219);
  nand2 I360_288(w_360_288, w_302_261, w_358_227);
  nand2 I360_315(w_360_315, w_186_361, w_121_004);
  nand2 I360_353(w_360_353, w_320_004, w_156_032);
  not1 I360_373(w_360_373, w_144_077);
  nand2 I360_383(w_360_383, w_212_034, w_320_318);
  or2  I360_414(w_360_414, w_253_074, w_075_007);
  and2 I360_419(w_360_419, w_091_039, w_239_000);
  nand2 I360_429(w_360_429, w_253_143, w_291_071);
  or2  I360_482(w_360_482, w_037_195, w_083_149);
  or2  I360_520(w_360_521, w_360_520, w_195_140);
  not1 I360_521(w_360_522, w_360_521);
  or2  I360_522(w_360_523, w_360_522, w_304_414);
  and2 I360_523(w_360_524, w_247_035, w_360_523);
  not1 I360_524(w_360_520, w_360_524);
  nand2 I361_031(w_361_031, w_127_047, w_343_251);
  or2  I361_070(w_361_070, w_203_433, w_292_298);
  or2  I361_097(w_361_097, w_359_074, w_214_457);
  or2  I361_104(w_361_104, w_089_144, w_249_202);
  or2  I361_200(w_361_200, w_076_157, w_232_190);
  and2 I361_221(w_361_221, w_307_095, w_182_015);
  not1 I361_249(w_361_249, w_282_166);
  and2 I361_354(w_361_354, w_203_259, w_256_550);
  nand2 I361_369(w_361_369, w_202_295, w_150_191);
  and2 I362_013(w_362_013, w_253_198, w_028_547);
  or2  I362_019(w_362_019, w_294_148, w_162_002);
  or2  I362_031(w_362_031, w_298_019, w_072_167);
  and2 I362_104(w_362_104, w_009_087, w_332_142);
  and2 I362_193(w_362_193, w_103_072, w_195_140);
  and2 I362_283(w_362_283, w_144_173, w_334_486);
  not1 I362_337(w_362_337, w_064_111);
  not1 I362_420(w_362_420, w_083_127);
  nand2 I363_009(w_363_009, w_266_160, w_146_311);
  not1 I363_056(w_363_056, w_107_151);
  not1 I363_057(w_363_057, w_198_030);
  nand2 I363_123(w_363_123, w_038_182, w_172_046);
  or2  I363_359(w_363_359, w_194_136, w_242_077);
  nand2 I363_372(w_363_372, w_085_176, w_228_123);
  not1 I364_009(w_364_009, w_194_021);
  nand2 I364_013(w_364_013, w_276_350, w_272_024);
  or2  I364_027(w_364_027, w_147_089, w_244_026);
  nand2 I365_045(w_365_045, w_208_175, w_307_040);
  and2 I365_106(w_365_106, w_165_003, w_009_601);
  or2  I365_128(w_365_128, w_148_650, w_145_035);
  not1 I365_196(w_365_196, w_081_009);
  and2 I365_199(w_365_199, w_287_354, w_032_021);
  not1 I365_252(w_365_252, w_182_021);
  or2  I365_390(w_365_390, w_280_448, w_112_063);
  or2  I366_013(w_366_013, w_047_251, w_241_081);
  or2  I366_072(w_366_072, w_085_024, w_083_073);
  not1 I366_144(w_366_144, w_347_021);
  and2 I366_174(w_366_174, w_051_033, w_069_078);
  or2  I366_238(w_366_238, w_365_252, w_322_001);
  nand2 I366_313(w_366_313, w_272_030, w_202_184);
  or2  I366_358(w_366_358, w_068_131, w_004_126);
  nand2 I367_035(w_367_035, w_010_209, w_341_245);
  not1 I367_075(w_367_075, w_064_034);
  or2  I367_123(w_367_123, w_359_051, w_197_098);
  nand2 I367_125(w_367_125, w_170_194, w_149_060);
  nand2 I367_160(w_367_160, w_242_163, w_209_033);
  nand2 I367_221(w_367_221, w_228_214, w_150_182);
  not1 I367_295(w_367_295, w_003_059);
  and2 I367_491(w_367_491, w_307_415, w_193_021);
  not1 I367_654(w_367_654, w_117_004);
  nand2 I367_755(w_367_755, w_269_564, w_227_339);
  nand2 I368_015(w_368_015, w_275_605, w_207_026);
  not1 I368_022(w_368_022, w_006_110);
  not1 I368_024(w_368_024, w_118_081);
  not1 I368_029(w_368_029, w_032_379);
  and2 I368_066(w_368_066, w_345_017, w_025_029);
  and2 I368_067(w_368_067, w_076_043, w_232_456);
  not1 I368_081(w_368_081, w_144_142);
  not1 I368_084(w_368_084, w_050_417);
  not1 I368_111(w_368_111, w_046_625);
  nand2 I369_115(w_369_115, w_331_025, w_137_013);
  and2 I369_133(w_369_133, w_100_014, w_223_073);
  not1 I369_282(w_369_282, w_137_146);
  and2 I369_524(w_369_524, w_037_042, w_367_755);
  nand2 I369_666(w_369_666, w_263_022, w_124_108);
  not1 I369_722(w_369_722, w_290_118);
  nand2 I369_739(w_369_741, w_028_028, w_369_740);
  and2 I369_740(w_369_742, w_355_295, w_369_741);
  not1 I369_741(w_369_743, w_369_742);
  not1 I369_742(w_369_744, w_369_743);
  and2 I369_743(w_369_745, w_217_023, w_369_744);
  and2 I369_744(w_369_740, w_369_745, w_369_757);
  and2 I369_745(w_369_750, w_238_449, w_369_749);
  or2  I369_746(w_369_751, w_336_124, w_369_750);
  and2 I369_747(w_369_752, w_079_056, w_369_751);
  not1 I369_748(w_369_753, w_369_752);
  and2 I369_749(w_369_754, w_284_022, w_369_753);
  and2 I369_750(w_369_755, w_158_002, w_369_754);
  not1 I369_751(w_369_749, w_369_740);
  and2 I369_752(w_369_757, w_022_390, w_369_755);
  and2 I369_753(w_369_760, w_369_759, w_265_450);
  or2  I369_754(w_369_761, w_369_760, w_165_026);
  and2 I369_755(w_369_762, w_369_761, w_101_194);
  and2 I369_756(w_369_763, w_369_762, w_369_775);
  not1 I369_757(w_369_759, w_369_763);
  or2  I369_758(w_369_768, w_180_013, w_369_767);
  or2  I369_759(w_369_769, w_207_049, w_369_768);
  not1 I369_760(w_369_770, w_369_769);
  or2  I369_761(w_369_771, w_369_770, w_023_044);
  and2 I369_762(w_369_772, w_107_005, w_369_771);
  and2 I369_763(w_369_773, w_156_386, w_369_772);
  not1 I369_764(w_369_767, w_369_763);
  and2 I369_765(w_369_775, w_299_053, w_369_773);
  or2  I370_020(w_370_020, w_100_106, w_038_471);
  or2  I370_031(w_370_031, w_283_003, w_293_021);
  not1 I370_051(w_370_051, w_355_100);
  not1 I370_056(w_370_056, w_368_066);
  not1 I370_065(w_370_065, w_329_094);
  nand2 I370_084(w_370_084, w_016_006, w_041_476);
  and2 I370_095(w_370_095, w_037_223, w_176_151);
  nand2 I370_099(w_370_099, w_314_159, w_129_275);
  and2 I370_104(w_369_747, w_352_411, w_369_740);
  and2 I370_105(w_369_765, w_369_747, w_369_759);
  or2  I371_000(w_371_000, w_369_765, w_072_163);
  and2 I372_000(w_372_000, w_147_031, w_255_062);
  not1 I372_003(w_372_003, w_340_010);
  or2  I372_008(w_372_008, w_090_242, w_127_048);
  and2 I372_031(w_372_031, w_238_412, w_242_002);
  not1 I372_033(w_372_033, w_183_243);
  not1 I372_038(w_372_038, w_011_118);
  or2  I373_001(w_373_001, w_277_038, w_169_283);
  or2  I373_013(w_373_013, w_271_188, w_327_097);
  nand2 I373_057(w_373_057, w_030_308, w_255_035);
  not1 I373_092(w_373_092, w_223_267);
  and2 I373_241(w_373_241, w_341_418, w_028_463);
  not1 I373_268(w_373_268, w_254_061);
  nand2 I373_327(w_373_327, w_050_388, w_096_005);
  or2  I374_056(w_374_056, w_270_284, w_141_050);
  nand2 I374_076(w_374_076, w_061_200, w_288_198);
  nand2 I374_091(w_374_091, w_061_257, w_186_093);
  and2 I374_141(w_374_141, w_172_035, w_238_429);
  nand2 I375_032(w_375_032, w_261_044, w_340_000);
  nand2 I375_071(w_375_071, w_315_634, w_190_066);
  not1 I375_142(w_375_142, w_004_026);
  not1 I375_171(w_375_171, w_349_036);
  and2 I375_178(w_375_178, w_180_007, w_042_443);
  or2  I375_189(w_375_191, w_006_111, w_375_190);
  nand2 I375_190(w_375_192, w_101_003, w_375_191);
  nand2 I375_191(w_375_193, w_070_292, w_375_192);
  and2 I375_192(w_375_194, w_375_193, w_375_214);
  and2 I375_193(w_375_195, w_375_194, w_254_065);
  nand2 I375_194(w_375_196, w_339_019, w_375_195);
  nand2 I375_195(w_375_197, w_375_196, w_049_259);
  not1 I375_196(w_375_198, w_375_197);
  or2  I375_197(w_375_199, w_037_023, w_375_198);
  and2 I375_198(w_375_200, w_375_199, w_341_704);
  and2 I375_199(w_375_190, w_288_068, w_375_200);
  not1 I375_200(w_375_205, w_375_204);
  or2  I375_201(w_375_206, w_375_205, w_006_223);
  not1 I375_202(w_375_207, w_375_206);
  or2  I375_203(w_375_208, w_375_207, w_122_031);
  and2 I375_204(w_375_209, w_113_258, w_375_208);
  not1 I375_205(w_375_210, w_375_209);
  nand2 I375_206(w_375_211, w_375_210, w_310_251);
  and2 I375_207(w_375_212, w_375_211, w_011_181);
  not1 I375_208(w_375_204, w_375_194);
  and2 I375_209(w_375_214, w_012_070, w_375_212);
  and2 I376_055(w_376_055, w_200_002, w_265_507);
  or2  I376_070(w_376_070, w_055_266, w_120_693);
  and2 I376_138(w_376_138, w_279_228, w_260_108);
  and2 I376_176(w_376_176, w_324_045, w_164_593);
  or2  I376_251(w_376_251, w_244_185, w_047_042);
  not1 I376_275(w_376_275, w_060_204);
  nand2 I376_276(w_376_278, w_376_277, w_105_282);
  nand2 I376_277(w_376_279, w_376_278, w_182_007);
  and2 I376_278(w_376_280, w_376_279, w_376_295);
  nand2 I376_279(w_376_281, w_376_280, w_263_120);
  nand2 I376_280(w_376_282, w_376_281, w_240_024);
  nand2 I376_281(w_376_283, w_376_282, w_020_410);
  not1 I376_282(w_376_284, w_376_283);
  or2  I376_283(w_376_285, w_291_022, w_376_284);
  and2 I376_284(w_376_286, w_075_058, w_376_285);
  or2  I376_285(w_376_277, w_171_711, w_376_286);
  or2  I376_286(w_376_291, w_247_184, w_376_290);
  or2  I376_287(w_376_292, w_376_291, w_022_241);
  and2 I376_288(w_376_293, w_376_292, w_261_041);
  not1 I376_289(w_376_290, w_376_280);
  and2 I376_290(w_376_295, w_267_065, w_376_293);
  nand2 I377_013(w_377_013, w_022_117, w_240_147);
  nand2 I377_040(w_377_040, w_037_153, w_279_026);
  not1 I377_065(w_377_065, w_240_104);
  and2 I377_066(w_377_066, w_160_080, w_158_000);
  nand2 I377_087(w_377_087, w_327_438, w_233_001);
  not1 I378_022(w_378_022, w_155_180);
  and2 I378_046(w_378_046, w_231_003, w_149_631);
  and2 I378_107(w_378_107, w_125_224, w_050_047);
  or2  I378_111(w_378_111, w_213_605, w_356_048);
  and2 I378_112(w_378_112, w_299_015, w_092_494);
  not1 I378_119(w_378_119, w_356_108);
  not1 I379_071(w_379_071, w_298_003);
  or2  I379_085(w_379_085, w_348_243, w_053_067);
  not1 I379_099(w_379_099, w_342_194);
  nand2 I379_103(w_379_103, w_078_597, w_310_447);
  or2  I379_182(w_379_182, w_022_154, w_220_248);
  not1 I379_186(w_379_186, w_110_242);
  or2  I380_035(w_380_035, w_176_008, w_338_028);
  or2  I380_162(w_380_162, w_091_105, w_084_046);
  or2  I380_284(w_380_284, w_040_599, w_143_408);
  not1 I380_296(w_380_296, w_214_381);
  and2 I380_317(w_380_317, w_103_063, w_076_134);
  not1 I380_615(w_380_615, w_175_549);
  nand2 I380_731(w_380_731, w_068_304, w_353_189);
  not1 I381_038(w_381_038, w_128_380);
  not1 I381_104(w_381_104, w_346_104);
  or2  I381_163(w_381_163, w_163_188, w_139_010);
  and2 I381_284(w_381_284, w_250_548, w_223_047);
  or2  I381_319(w_381_319, w_343_425, w_021_199);
  or2  I381_653(w_381_653, w_124_105, w_280_019);
  and2 I381_670(w_381_670, w_125_204, w_148_209);
  and2 I382_033(w_382_033, w_130_230, w_280_503);
  or2  I382_046(w_382_046, w_164_023, w_322_014);
  and2 I382_341(w_382_341, w_145_011, w_227_209);
  or2  I382_477(w_382_477, w_301_197, w_182_011);
  and2 I382_563(w_382_563, w_354_207, w_160_092);
  and2 I382_615(w_382_615, w_245_735, w_340_038);
  nand2 I383_018(w_383_018, w_138_221, w_053_140);
  and2 I383_031(w_383_031, w_085_226, w_382_477);
  nand2 I383_092(w_383_092, w_044_050, w_311_439);
  and2 I383_112(w_383_112, w_212_218, w_377_040);
  and2 I383_240(w_383_240, w_192_010, w_198_044);
  not1 I383_350(w_383_350, w_214_016);
  not1 I383_394(w_383_394, w_367_075);
  nand2 I383_450(w_383_450, w_332_363, w_024_071);
  or2  I383_455(w_383_455, w_048_008, w_142_303);
  or2  I383_591(w_383_591, w_073_621, w_343_246);
  not1 I383_618(w_383_618, w_001_004);
  or2  I383_732(w_383_734, w_138_067, w_383_733);
  not1 I383_733(w_383_735, w_383_734);
  or2  I383_734(w_383_736, w_383_735, w_044_407);
  nand2 I383_735(w_383_737, w_034_055, w_383_736);
  nand2 I383_736(w_383_738, w_383_737, w_148_528);
  and2 I383_737(w_383_739, w_383_738, w_156_231);
  and2 I383_738(w_383_733, w_051_246, w_383_739);
  nand2 I383_739(w_383_744, w_383_743, w_204_218);
  nand2 I383_740(w_383_745, w_383_744, w_268_237);
  nand2 I383_741(w_383_746, w_357_005, w_383_745);
  or2  I383_742(w_383_747, w_212_226, w_383_746);
  not1 I383_743(w_383_748, w_383_747);
  and2 I383_744(w_383_749, w_383_758, w_383_748);
  nand2 I383_745(w_383_743, w_383_749, w_033_539);
  not1 I383_746(w_383_754, w_383_753);
  and2 I383_747(w_383_755, w_254_053, w_383_754);
  and2 I383_748(w_383_756, w_383_755, w_054_186);
  not1 I383_749(w_383_753, w_383_749);
  and2 I383_750(w_383_758, w_334_368, w_383_756);
  not1 I383_751(w_383_761, w_383_760);
  and2 I383_752(w_383_762, w_087_165, w_383_761);
  not1 I383_753(w_383_763, w_383_762);
  nand2 I383_754(w_383_764, w_383_763, w_383_782);
  not1 I383_755(w_383_765, w_383_764);
  or2  I383_756(w_383_766, w_364_009, w_383_765);
  nand2 I383_757(w_383_767, w_154_010, w_383_766);
  or2  I383_758(w_383_768, w_383_767, w_359_041);
  nand2 I383_759(w_383_769, w_183_194, w_383_768);
  and2 I383_760(w_383_770, w_321_536, w_383_769);
  and2 I383_761(w_383_771, w_249_268, w_383_770);
  or2  I383_762(w_383_760, w_310_365, w_383_771);
  nand2 I383_763(w_383_776, w_383_775, w_373_268);
  and2 I383_764(w_383_777, w_095_022, w_383_776);
  or2  I383_765(w_383_778, w_383_777, w_149_364);
  nand2 I383_766(w_383_779, w_383_778, w_001_030);
  and2 I383_767(w_383_780, w_383_779, w_205_186);
  not1 I383_768(w_383_775, w_383_764);
  and2 I383_769(w_383_782, w_016_000, w_383_780);
  not1 I384_042(w_384_042, w_240_005);
  and2 I384_046(w_384_046, w_045_315, w_009_497);
  nand2 I384_121(w_384_121, w_160_398, w_105_198);
  nand2 I384_149(w_384_149, w_092_001, w_362_013);
  nand2 I384_162(w_384_162, w_191_052, w_103_113);
  and2 I384_197(w_383_741, w_220_142, w_383_733);
  and2 I384_199(w_383_773, w_172_035, w_383_760);
  nand2 I385_007(w_385_007, w_383_741, w_204_056);
  nand2 I385_089(w_385_089, w_383_773, w_084_003);
  and2 I385_106(w_385_106, w_281_551, w_355_192);
  or2  I385_124(w_385_124, w_186_262, w_199_253);
  or2  I385_213(w_385_213, w_292_494, w_225_220);
  not1 I385_227(w_385_227, w_318_012);
  nand2 I385_427(w_385_427, w_255_042, w_275_603);
  or2  I385_429(w_385_429, w_072_288, w_239_000);
  and2 I386_015(w_386_015, w_324_012, w_288_158);
  nand2 I386_041(w_386_041, w_191_069, w_384_162);
  not1 I386_080(w_386_080, w_161_294);
  or2  I386_115(w_386_115, w_200_061, w_036_110);
  and2 I386_146(w_386_146, w_240_171, w_159_101);
  nand2 I386_152(w_386_152, w_212_202, w_144_228);
  and2 I386_161(w_386_161, w_257_110, w_344_001);
  not1 I386_188(w_386_188, w_051_166);
  and2 I386_226(w_386_226, w_091_034, w_344_088);
  nand2 I386_473(w_386_473, w_277_143, w_042_002);
  nand2 I387_012(w_387_012, w_261_015, w_024_354);
  or2  I387_219(w_387_219, w_336_074, w_171_263);
  nand2 I387_252(w_387_252, w_264_273, w_242_153);
  not1 I388_012(w_388_012, w_123_067);
  and2 I388_025(w_388_025, w_003_010, w_173_013);
  not1 I388_057(w_388_057, w_311_325);
  not1 I388_076(w_388_076, w_312_432);
  and2 I388_090(w_388_090, w_267_054, w_261_029);
  nand2 I388_100(w_388_100, w_122_001, w_122_032);
  and2 I388_159(w_388_159, w_373_241, w_300_610);
  and2 I389_066(w_389_066, w_301_220, w_226_152);
  or2  I389_087(w_389_087, w_119_106, w_177_375);
  and2 I389_150(w_389_150, w_313_118, w_311_256);
  and2 I389_234(w_389_234, w_213_479, w_154_099);
  not1 I389_279(w_389_279, w_154_046);
  nand2 I389_308(w_389_308, w_098_033, w_115_122);
  or2  I389_437(w_389_437, w_260_027, w_165_111);
  and2 I390_031(w_390_031, w_386_226, w_105_001);
  and2 I390_054(w_390_054, w_319_077, w_344_116);
  or2  I390_138(w_390_138, w_313_254, w_230_037);
  not1 I390_148(w_390_148, w_069_176);
  not1 I390_173(w_390_173, w_102_070);
  nand2 I390_187(w_390_187, w_021_028, w_029_073);
  or2  I390_252(w_390_252, w_342_111, w_065_000);
  or2  I391_100(w_391_100, w_212_006, w_312_056);
  and2 I391_105(w_391_105, w_160_601, w_065_522);
  nand2 I391_249(w_391_249, w_280_306, w_123_195);
  nand2 I391_463(w_391_463, w_284_113, w_326_043);
  not1 I391_491(w_391_491, w_311_080);
  or2  I391_610(w_391_610, w_214_550, w_364_013);
  or2  I391_670(w_391_670, w_131_263, w_104_053);
  or2  I391_738(w_391_738, w_303_070, w_097_175);
  or2  I392_081(w_392_081, w_060_344, w_073_068);
  not1 I392_083(w_392_083, w_264_743);
  and2 I392_185(w_392_185, w_051_381, w_056_627);
  nand2 I392_244(w_392_244, w_340_026, w_203_444);
  and2 I392_245(w_392_245, w_281_089, w_239_000);
  and2 I392_262(w_392_262, w_266_533, w_281_283);
  and2 I392_551(w_392_553, w_392_572, w_392_552);
  not1 I392_552(w_392_554, w_392_553);
  not1 I392_553(w_392_555, w_392_554);
  and2 I392_554(w_392_556, w_392_555, w_190_074);
  or2  I392_555(w_392_552, w_392_556, w_165_110);
  or2  I392_556(w_392_561, w_392_560, w_351_228);
  or2  I392_557(w_392_562, w_392_561, w_182_018);
  and2 I392_558(w_392_563, w_182_023, w_392_562);
  not1 I392_559(w_392_564, w_392_563);
  and2 I392_560(w_392_565, w_077_626, w_392_564);
  and2 I392_561(w_392_566, w_164_502, w_392_565);
  nand2 I392_562(w_392_567, w_011_217, w_392_566);
  nand2 I392_563(w_392_568, w_306_236, w_392_567);
  nand2 I392_564(w_392_569, w_336_140, w_392_568);
  and2 I392_565(w_392_570, w_392_569, w_221_033);
  not1 I392_566(w_392_560, w_392_553);
  and2 I392_567(w_392_572, w_338_049, w_392_570);
  not1 I393_003(w_393_003, w_340_013);
  nand2 I393_016(w_393_016, w_033_419, w_387_219);
  nand2 I393_020(w_393_020, w_130_191, w_331_315);
  or2  I393_050(w_393_050, w_379_085, w_360_419);
  nand2 I393_084(w_393_084, w_197_247, w_313_128);
  or2  I393_102(w_393_102, w_007_452, w_256_028);
  not1 I393_109(w_393_109, w_343_580);
  and2 I393_113(w_393_113, w_146_133, w_042_222);
  nand2 I393_129(w_393_129, w_368_084, w_011_203);
  or2  I393_136(w_393_136, w_186_223, w_391_738);
  and2 I393_149(w_393_149, w_213_315, w_014_240);
  nand2 I393_194(w_393_194, w_000_444, w_192_175);
  nand2 I393_204(w_393_204, w_182_023, w_279_160);
  not1 I393_238(w_393_240, w_393_239);
  or2  I393_239(w_393_241, w_393_262, w_393_240);
  not1 I393_240(w_393_242, w_393_241);
  or2  I393_241(w_393_243, w_393_242, w_347_268);
  not1 I393_242(w_393_244, w_393_243);
  not1 I393_243(w_393_245, w_393_244);
  and2 I393_244(w_393_246, w_205_353, w_393_245);
  and2 I393_245(w_393_239, w_042_094, w_393_246);
  or2  I393_246(w_393_251, w_287_019, w_393_250);
  and2 I393_247(w_393_252, w_063_109, w_393_251);
  and2 I393_248(w_393_253, w_393_252, w_391_249);
  or2  I393_249(w_393_254, w_393_253, w_086_003);
  nand2 I393_250(w_393_255, w_393_254, w_254_054);
  not1 I393_251(w_393_256, w_393_255);
  nand2 I393_252(w_393_257, w_393_256, w_158_001);
  and2 I393_253(w_393_258, w_056_235, w_393_257);
  nand2 I393_254(w_393_259, w_247_170, w_393_258);
  and2 I393_255(w_393_260, w_043_033, w_393_259);
  not1 I393_256(w_393_250, w_393_241);
  and2 I393_257(w_393_262, w_029_058, w_393_260);
  nand2 I394_040(w_394_040, w_094_544, w_166_279);
  and2 I394_070(w_394_070, w_208_083, w_185_039);
  nand2 I394_080(w_394_080, w_194_241, w_091_080);
  nand2 I394_107(w_394_107, w_167_082, w_291_030);
  or2  I395_029(w_395_029, w_368_067, w_004_014);
  or2  I395_041(w_395_041, w_304_468, w_251_035);
  and2 I395_072(w_395_072, w_164_093, w_365_196);
  or2  I395_080(w_395_080, w_075_087, w_048_002);
  or2  I395_229(w_395_229, w_189_446, w_041_676);
  not1 I395_235(w_395_235, w_103_114);
  and2 I395_290(w_395_290, w_069_232, w_268_058);
  or2  I395_372(w_395_372, w_194_304, w_076_201);
  and2 I396_004(w_396_004, w_341_408, w_119_157);
  not1 I396_007(w_396_007, w_070_100);
  not1 I396_025(w_396_025, w_195_208);
  nand2 I396_045(w_396_045, w_113_267, w_384_121);
  and2 I396_065(w_396_065, w_033_656, w_183_139);
  nand2 I397_018(w_397_018, w_355_051, w_060_387);
  and2 I397_019(w_397_019, w_120_638, w_277_203);
  not1 I397_036(w_397_036, w_093_245);
  nand2 I397_046(w_397_046, w_136_011, w_180_021);
  and2 I397_048(w_397_048, w_015_259, w_285_091);
  and2 I397_050(w_397_050, w_224_104, w_335_134);
  not1 I397_060(w_397_060, w_231_198);
  or2  I397_064(w_397_064, w_295_092, w_391_491);
  and2 I397_081(w_397_081, w_014_117, w_240_098);
  not1 I397_092(w_397_092, w_281_710);
  not1 I397_137(w_397_137, w_103_059);
  nand2 I397_141(w_397_141, w_127_074, w_293_226);
  and2 I398_023(w_398_023, w_189_471, w_353_244);
  or2  I398_029(w_398_029, w_287_394, w_291_108);
  or2  I398_043(w_398_043, w_082_058, w_095_046);
  or2  I398_050(w_398_050, w_173_022, w_272_038);
  not1 I398_058(w_398_058, w_125_561);
  not1 I398_061(w_398_061, w_329_306);
  nand2 I398_067(w_398_067, w_232_478, w_172_001);
  or2  I398_074(w_398_074, w_383_031, w_291_043);
  or2  I399_023(w_399_023, w_122_081, w_285_104);
  and2 I399_035(w_399_035, w_203_271, w_163_178);
  and2 I399_098(w_399_098, w_012_007, w_030_236);
  nand2 I399_118(w_399_118, w_276_264, w_058_081);
  and2 I399_137(w_399_137, w_397_050, w_337_036);
  or2  I399_163(w_399_163, w_024_317, w_098_022);
  or2  I399_285(w_399_285, w_074_297, w_049_260);
  and2 I399_297(w_399_297, w_187_020, w_232_079);
  not1 I400_009(w_400_009, w_213_017);
  not1 I400_024(w_400_024, w_246_079);
  not1 I400_051(w_400_051, w_150_197);
  or2  I400_091(w_400_091, w_319_347, w_342_344);
  and2 I401_008(w_401_008, w_148_371, w_389_437);
  not1 I401_079(w_401_079, w_024_215);
  nand2 I401_158(w_401_158, w_018_019, w_155_024);
  not1 I401_170(w_401_170, w_224_401);
  and2 I401_178(w_401_178, w_320_309, w_277_373);
  nand2 I401_205(w_401_205, w_077_054, w_056_476);
  and2 I401_230(w_401_230, w_267_298, w_228_584);
  not1 I401_244(w_401_244, w_011_060);
  or2  I401_246(w_401_246, w_290_128, w_109_238);
  and2 I402_021(w_402_021, w_042_152, w_319_129);
  nand2 I402_027(w_402_027, w_329_039, w_391_670);
  not1 I402_028(w_402_028, w_154_075);
  not1 I402_032(w_402_032, w_225_062);
  or2  I402_068(w_402_068, w_080_313, w_015_426);
  and2 I402_080(w_402_080, w_009_115, w_147_061);
  not1 I402_087(w_402_087, w_135_013);
  and2 I402_114(w_402_114, w_350_071, w_179_737);
  not1 I402_135(w_402_135, w_091_135);
  not1 I403_120(w_403_120, w_291_044);
  or2  I403_216(w_403_216, w_087_235, w_058_280);
  or2  I403_289(w_403_289, w_168_216, w_281_740);
  or2  I403_315(w_403_315, w_099_263, w_382_615);
  nand2 I403_325(w_403_325, w_089_078, w_069_033);
  or2  I403_439(w_403_439, w_171_252, w_066_185);
  or2  I404_022(w_404_022, w_139_026, w_138_214);
  or2  I404_182(w_404_182, w_380_162, w_133_334);
  not1 I404_196(w_404_196, w_056_710);
  nand2 I404_339(w_404_339, w_357_096, w_305_057);
  not1 I404_361(w_404_361, w_136_059);
  and2 I404_588(w_404_588, w_147_077, w_337_028);
  not1 I404_606(w_404_606, w_018_037);
  nand2 I404_648(w_404_648, w_237_062, w_215_246);
  and2 I405_026(w_405_026, w_306_146, w_212_117);
  or2  I405_027(w_405_027, w_032_168, w_386_041);
  nand2 I405_071(w_405_071, w_397_060, w_262_371);
  not1 I405_073(w_405_073, w_352_047);
  or2  I405_132(w_405_132, w_029_105, w_370_065);
  or2  I405_137(w_405_137, w_252_386, w_130_204);
  not1 I405_166(w_405_166, w_007_035);
  and2 I405_182(w_405_182, w_190_009, w_237_128);
  nand2 I406_004(w_406_004, w_020_546, w_026_013);
  nand2 I406_022(w_406_022, w_013_078, w_097_007);
  and2 I406_050(w_406_050, w_105_274, w_180_010);
  or2  I406_116(w_406_116, w_356_039, w_127_022);
  and2 I406_221(w_406_221, w_134_185, w_283_126);
  and2 I406_280(w_406_280, w_163_162, w_091_162);
  or2  I406_282(w_406_282, w_313_240, w_244_220);
  or2  I407_063(w_407_063, w_358_295, w_032_189);
  and2 I407_070(w_407_070, w_348_137, w_368_111);
  and2 I407_133(w_407_133, w_038_311, w_084_048);
  nand2 I407_267(w_407_267, w_010_204, w_123_538);
  or2  I407_293(w_407_293, w_320_178, w_318_014);
  and2 I407_356(w_407_356, w_190_073, w_012_002);
  nand2 I407_572(w_407_572, w_119_156, w_211_003);
  nand2 I407_643(w_407_643, w_044_460, w_229_268);
  or2  I408_002(w_408_002, w_327_444, w_265_064);
  nand2 I408_003(w_408_003, w_244_111, w_148_279);
  nand2 I408_004(w_408_004, w_299_164, w_173_005);
  not1 I408_005(w_408_005, w_309_034);
  or2  I409_049(w_409_049, w_094_317, w_137_354);
  or2  I409_153(w_409_153, w_318_011, w_236_028);
  or2  I409_304(w_409_304, w_299_270, w_235_018);
  or2  I409_408(w_409_408, w_190_093, w_141_149);
  or2  I409_455(w_409_455, w_136_057, w_026_169);
  and2 I410_011(w_410_011, w_018_023, w_159_013);
  not1 I410_027(w_410_027, w_140_071);
  nand2 I410_048(w_410_048, w_313_258, w_114_116);
  not1 I410_064(w_410_064, w_314_014);
  nand2 I410_085(w_410_085, w_307_043, w_405_166);
  or2  I410_102(w_410_102, w_216_410, w_221_067);
  not1 I410_142(w_410_142, w_282_265);
  and2 I411_130(w_411_130, w_281_462, w_385_429);
  not1 I411_567(w_411_567, w_267_067);
  and2 I411_581(w_411_581, w_285_184, w_050_101);
  and2 I412_076(w_412_076, w_164_395, w_355_297);
  or2  I412_202(w_412_202, w_267_155, w_052_042);
  not1 I412_275(w_412_275, w_392_262);
  and2 I412_300(w_412_300, w_046_360, w_150_159);
  not1 I412_374(w_412_374, w_111_010);
  and2 I412_398(w_412_398, w_316_149, w_346_565);
  not1 I413_015(w_413_015, w_293_101);
  and2 I413_022(w_413_022, w_115_215, w_349_028);
  nand2 I413_029(w_413_029, w_145_027, w_217_068);
  nand2 I413_045(w_413_045, w_054_365, w_220_380);
  or2  I413_083(w_413_083, w_186_212, w_067_150);
  or2  I414_089(w_414_089, w_294_070, w_326_111);
  or2  I414_151(w_414_151, w_296_200, w_253_344);
  or2  I414_241(w_414_241, w_309_301, w_407_063);
  not1 I414_303(w_414_303, w_129_048);
  or2  I414_325(w_414_325, w_116_576, w_295_122);
  nand2 I415_046(w_415_046, w_082_020, w_318_013);
  and2 I415_050(w_415_050, w_156_172, w_078_200);
  nand2 I415_072(w_415_072, w_321_063, w_339_020);
  or2  I415_079(w_415_079, w_237_107, w_293_067);
  nand2 I415_283(w_415_283, w_298_038, w_085_026);
  or2  I416_134(w_416_134, w_367_221, w_184_033);
  or2  I416_168(w_416_168, w_323_230, w_132_188);
  and2 I416_325(w_416_325, w_253_059, w_103_108);
  nand2 I416_344(w_416_344, w_122_058, w_266_043);
  not1 I416_427(w_416_427, w_272_031);
  nand2 I417_050(w_417_050, w_162_019, w_313_403);
  not1 I417_057(w_417_057, w_365_106);
  nand2 I417_060(w_417_060, w_262_321, w_070_542);
  and2 I417_065(w_417_065, w_050_578, w_230_024);
  or2  I417_075(w_417_075, w_135_661, w_056_596);
  and2 I417_083(w_417_083, w_054_167, w_085_037);
  nand2 I417_100(w_417_100, w_215_049, w_027_141);
  nand2 I417_116(w_417_116, w_001_024, w_081_003);
  not1 I417_120(w_417_120, w_167_131);
  and2 I417_137(w_417_137, w_070_000, w_363_057);
  and2 I418_029(w_418_029, w_097_166, w_294_083);
  and2 I418_045(w_418_045, w_044_447, w_010_352);
  nand2 I418_048(w_418_048, w_173_026, w_143_353);
  or2  I418_052(w_418_052, w_269_441, w_157_098);
  nand2 I418_068(w_418_068, w_003_035, w_398_061);
  nand2 I418_091(w_418_091, w_279_302, w_175_141);
  or2  I418_105(w_418_105, w_026_315, w_225_033);
  not1 I419_044(w_419_044, w_272_028);
  not1 I419_139(w_419_139, w_224_386);
  nand2 I419_155(w_419_155, w_067_342, w_280_282);
  nand2 I419_240(w_419_240, w_048_005, w_268_035);
  or2  I419_308(w_419_308, w_075_117, w_063_524);
  not1 I419_323(w_419_325, w_419_324);
  nand2 I419_324(w_419_326, w_102_248, w_419_325);
  and2 I419_325(w_419_327, w_419_326, w_419_336);
  and2 I419_326(w_419_328, w_419_327, w_379_103);
  or2  I419_327(w_419_324, w_419_328, w_086_051);
  nand2 I419_328(w_419_333, w_419_332, w_374_076);
  and2 I419_329(w_419_334, w_419_333, w_014_114);
  not1 I419_330(w_419_332, w_419_327);
  and2 I419_331(w_419_336, w_243_150, w_419_334);
  nand2 I420_161(w_420_161, w_207_152, w_253_163);
  or2  I420_483(w_420_483, w_171_384, w_389_308);
  not1 I420_519(w_420_519, w_242_122);
  nand2 I420_574(w_420_574, w_155_242, w_241_058);
  and2 I420_587(w_420_587, w_009_108, w_202_231);
  not1 I420_607(w_420_607, w_362_104);
  and2 I420_673(w_420_673, w_301_066, w_044_243);
  or2  I421_047(w_421_047, w_316_410, w_151_268);
  nand2 I421_052(w_421_052, w_094_434, w_343_697);
  and2 I421_075(w_421_075, w_195_232, w_131_029);
  nand2 I421_126(w_421_126, w_277_315, w_284_054);
  or2  I421_243(w_421_243, w_083_192, w_408_003);
  nand2 I422_001(w_422_001, w_123_169, w_417_137);
  nand2 I422_002(w_422_002, w_333_115, w_043_036);
  and2 I422_005(w_422_005, w_110_304, w_154_054);
  nand2 I422_007(w_422_007, w_029_001, w_287_274);
  and2 I422_008(w_422_008, w_152_468, w_195_100);
  not1 I422_010(w_422_010, w_239_000);
  nand2 I422_013(w_422_013, w_401_170, w_271_142);
  nand2 I423_019(w_423_019, w_326_113, w_403_439);
  or2  I423_021(w_423_021, w_408_004, w_071_014);
  or2  I423_022(w_423_022, w_151_088, w_421_243);
  or2  I423_038(w_423_038, w_258_026, w_227_403);
  not1 I423_052(w_423_052, w_097_207);
  nand2 I423_057(w_423_057, w_367_654, w_294_118);
  not1 I423_073(w_423_073, w_021_199);
  not1 I423_075(w_423_075, w_163_445);
  and2 I423_092(w_423_092, w_217_031, w_007_212);
  nand2 I424_087(w_424_087, w_280_444, w_368_024);
  not1 I424_111(w_424_111, w_391_463);
  or2  I424_156(w_424_156, w_169_192, w_075_133);
  not1 I424_222(w_424_222, w_381_670);
  nand2 I424_228(w_424_228, w_256_515, w_341_487);
  or2  I425_000(w_425_000, w_347_252, w_170_185);
  and2 I425_102(w_425_102, w_392_244, w_158_003);
  not1 I425_214(w_425_214, w_133_378);
  not1 I425_247(w_425_247, w_101_170);
  and2 I425_358(w_425_358, w_062_157, w_330_042);
  nand2 I425_362(w_425_362, w_268_113, w_079_005);
  or2  I425_550(w_425_552, w_148_085, w_425_551);
  and2 I425_551(w_425_553, w_309_270, w_425_552);
  and2 I425_552(w_425_554, w_108_001, w_425_553);
  or2  I425_553(w_425_555, w_386_152, w_425_554);
  not1 I425_554(w_425_556, w_425_555);
  and2 I425_555(w_425_557, w_119_017, w_425_556);
  and2 I425_556(w_425_558, w_425_567, w_425_557);
  and2 I425_557(w_425_551, w_425_558, w_033_511);
  not1 I425_558(w_425_563, w_425_562);
  not1 I425_559(w_425_564, w_425_563);
  and2 I425_560(w_425_565, w_425_564, w_413_022);
  not1 I425_561(w_425_562, w_425_558);
  and2 I425_562(w_425_567, w_071_129, w_425_565);
  not1 I426_017(w_426_017, w_366_313);
  not1 I426_022(w_426_022, w_351_075);
  not1 I426_162(w_426_162, w_421_126);
  nand2 I427_050(w_427_050, w_161_013, w_341_458);
  nand2 I427_051(w_427_051, w_130_122, w_152_108);
  nand2 I427_053(w_427_053, w_276_326, w_213_013);
  nand2 I427_059(w_427_059, w_366_013, w_381_038);
  or2  I428_010(w_428_010, w_065_263, w_257_257);
  not1 I428_124(w_428_124, w_025_007);
  not1 I428_181(w_428_181, w_239_000);
  or2  I429_003(w_429_003, w_095_057, w_212_163);
  nand2 I429_085(w_429_085, w_069_207, w_321_141);
  nand2 I429_096(w_429_096, w_339_041, w_079_010);
  and2 I429_115(w_429_115, w_069_177, w_141_018);
  not1 I429_130(w_429_130, w_294_064);
  nand2 I429_137(w_429_137, w_113_187, w_163_081);
  or2  I429_218(w_429_218, w_374_141, w_426_022);
  nand2 I429_236(w_429_236, w_332_004, w_033_580);
  not1 I429_259(w_429_259, w_231_157);
  and2 I430_060(w_430_060, w_020_306, w_134_109);
  nand2 I430_092(w_430_092, w_085_022, w_238_105);
  not1 I430_114(w_430_114, w_315_362);
  nand2 I430_286(w_430_286, w_173_027, w_329_384);
  not1 I430_422(w_430_422, w_304_100);
  and2 I430_484(w_430_484, w_380_284, w_250_367);
  not1 I430_534(w_430_534, w_175_019);
  and2 I431_210(w_431_210, w_110_175, w_193_169);
  or2  I432_051(w_432_051, w_384_042, w_235_066);
  not1 I432_053(w_432_053, w_395_072);
  and2 I432_120(w_432_120, w_398_029, w_399_035);
  and2 I432_136(w_432_136, w_187_019, w_315_269);
  not1 I432_218(w_432_218, w_239_000);
  nand2 I432_288(w_432_288, w_383_455, w_312_042);
  not1 I432_300(w_432_300, w_245_465);
  and2 I432_307(w_432_307, w_041_160, w_103_292);
  not1 I432_313(w_432_313, w_282_031);
  and2 I433_054(w_433_054, w_178_075, w_277_317);
  not1 I433_120(w_433_120, w_088_031);
  not1 I433_180(w_433_180, w_227_658);
  not1 I433_213(w_433_213, w_387_012);
  not1 I433_268(w_433_268, w_253_318);
  not1 I433_398(w_433_398, w_068_340);
  not1 I433_409(w_433_409, w_222_255);
  and2 I433_444(w_433_444, w_361_104, w_072_051);
  or2  I434_061(w_434_061, w_125_072, w_331_052);
  not1 I434_098(w_434_098, w_111_049);
  and2 I434_335(w_434_335, w_023_028, w_176_002);
  not1 I434_382(w_434_382, w_151_222);
  nand2 I434_495(w_434_495, w_357_304, w_117_059);
  and2 I435_075(w_435_075, w_313_080, w_377_087);
  and2 I435_085(w_435_085, w_101_284, w_059_032);
  or2  I435_136(w_435_136, w_304_192, w_087_298);
  or2  I435_156(w_435_156, w_263_106, w_211_018);
  not1 I436_218(w_436_218, w_324_031);
  and2 I436_224(w_436_224, w_084_016, w_281_627);
  not1 I436_410(w_436_410, w_283_094);
  nand2 I436_562(w_436_562, w_388_090, w_015_562);
  and2 I436_564(w_436_564, w_183_202, w_351_106);
  nand2 I437_010(w_437_010, w_343_335, w_206_157);
  or2  I437_429(w_437_429, w_184_073, w_413_029);
  nand2 I438_084(w_438_084, w_224_156, w_177_006);
  or2  I438_253(w_438_253, w_294_037, w_359_090);
  not1 I438_273(w_438_273, w_282_150);
  and2 I439_038(w_439_038, w_054_089, w_304_083);
  nand2 I439_039(w_439_039, w_373_013, w_244_136);
  or2  I439_045(w_439_045, w_005_002, w_093_080);
  nand2 I439_116(w_439_116, w_333_137, w_225_059);
  not1 I439_295(w_439_295, w_046_189);
  and2 I439_313(w_439_313, w_341_599, w_330_059);
  not1 I440_032(w_440_032, w_131_101);
  or2  I440_037(w_440_037, w_275_291, w_319_218);
  nand2 I440_040(w_440_040, w_068_204, w_299_315);
  or2  I440_057(w_440_057, w_213_078, w_222_623);
  not1 I440_064(w_440_064, w_287_279);
  and2 I440_079(w_440_079, w_318_003, w_402_080);
  not1 I441_007(w_441_007, w_372_003);
  and2 I441_023(w_441_023, w_295_020, w_137_123);
  nand2 I441_144(w_441_144, w_372_000, w_032_115);
  and2 I441_407(w_441_407, w_069_063, w_331_153);
  and2 I441_505(w_441_505, w_145_032, w_395_235);
  or2  I442_045(w_442_045, w_090_203, w_397_064);
  and2 I442_104(w_442_104, w_166_313, w_366_358);
  or2  I442_123(w_442_123, w_057_105, w_213_392);
  nand2 I442_126(w_442_126, w_156_430, w_001_010);
  and2 I442_135(w_442_135, w_293_149, w_030_185);
  or2  I442_141(w_442_143, w_442_142, w_393_050);
  or2  I442_142(w_442_144, w_068_176, w_442_143);
  and2 I442_143(w_442_145, w_442_144, w_442_161);
  not1 I442_144(w_442_142, w_442_145);
  nand2 I442_145(w_442_150, w_442_149, w_378_119);
  and2 I442_146(w_442_151, w_277_258, w_442_150);
  and2 I442_147(w_442_152, w_442_151, w_183_073);
  or2  I442_148(w_442_153, w_442_152, w_167_068);
  and2 I442_149(w_442_154, w_231_056, w_442_153);
  and2 I442_150(w_442_155, w_143_061, w_442_154);
  nand2 I442_151(w_442_156, w_336_029, w_442_155);
  not1 I442_152(w_442_157, w_442_156);
  not1 I442_153(w_442_158, w_442_157);
  and2 I442_154(w_442_159, w_442_158, w_079_037);
  not1 I442_155(w_442_149, w_442_145);
  and2 I442_156(w_442_161, w_412_275, w_442_159);
  nand2 I443_130(w_443_130, w_092_572, w_215_335);
  nand2 I443_263(w_443_263, w_118_019, w_060_212);
  not1 I443_327(w_443_327, w_155_033);
  not1 I444_022(w_444_022, w_165_032);
  and2 I444_101(w_444_101, w_362_283, w_152_348);
  not1 I444_165(w_444_165, w_058_656);
  or2  I444_307(w_444_307, w_385_007, w_314_191);
  and2 I444_425(w_444_425, w_258_138, w_283_219);
  and2 I444_462(w_444_462, w_101_085, w_250_588);
  not1 I444_520(w_444_520, w_096_005);
  nand2 I444_585(w_444_585, w_163_491, w_318_004);
  not1 I444_709(w_444_709, w_122_093);
  and2 I445_012(w_445_012, w_100_058, w_380_035);
  nand2 I445_021(w_445_021, w_149_261, w_208_277);
  and2 I445_025(w_445_025, w_251_037, w_422_007);
  and2 I445_029(w_445_029, w_390_138, w_359_170);
  nand2 I445_069(w_445_069, w_232_084, w_184_132);
  and2 I445_135(w_445_135, w_360_266, w_391_610);
  or2  I445_181(w_445_183, w_445_182, w_163_249);
  nand2 I445_182(w_445_184, w_445_183, w_213_303);
  and2 I445_183(w_445_185, w_445_184, w_202_033);
  or2  I445_184(w_445_186, w_445_185, w_351_049);
  or2  I445_185(w_445_187, w_445_186, w_269_363);
  nand2 I445_186(w_445_188, w_445_187, w_417_100);
  or2  I445_187(w_445_189, w_166_202, w_445_188);
  not1 I445_188(w_445_190, w_445_189);
  not1 I445_189(w_445_191, w_445_190);
  and2 I445_190(w_445_192, w_445_191, w_041_403);
  nand2 I445_191(w_445_182, w_268_216, w_445_192);
  nand2 I445_192(w_445_197, w_317_148, w_445_196);
  not1 I445_193(w_445_198, w_445_197);
  and2 I445_194(w_445_199, w_235_062, w_445_198);
  or2  I445_195(w_445_200, w_445_199, w_314_092);
  not1 I445_196(w_445_201, w_445_200);
  or2  I445_197(w_445_202, w_445_201, w_130_321);
  and2 I445_198(w_445_203, w_445_202, w_159_024);
  not1 I445_199(w_445_204, w_445_203);
  nand2 I445_200(w_445_205, w_034_065, w_445_204);
  and2 I445_201(w_445_206, w_445_205, w_229_034);
  and2 I445_202(w_445_207, w_445_206, w_129_106);
  or2  I445_203(w_445_196, w_360_429, w_445_207);
  nand2 I445_204(w_445_212, w_445_211, w_029_004);
  not1 I445_205(w_445_213, w_445_212);
  or2  I445_206(w_445_214, w_445_213, w_268_214);
  and2 I445_207(w_445_215, w_445_214, w_430_286);
  nand2 I445_208(w_445_211, w_445_215, w_425_358);
  not1 I446_025(w_446_025, w_252_242);
  nand2 I446_151(w_446_151, w_093_360, w_091_044);
  or2  I446_152(w_446_152, w_347_036, w_298_000);
  not1 I446_242(w_446_242, w_285_057);
  and2 I446_298(w_446_298, w_310_093, w_131_483);
  and2 I446_406(w_446_406, w_125_025, w_412_374);
  nand2 I446_438(w_446_438, w_395_372, w_408_004);
  and2 I446_533(w_446_533, w_276_050, w_149_004);
  or2  I446_544(w_446_544, w_185_140, w_376_070);
  nand2 I446_577(w_446_577, w_061_175, w_347_257);
  and2 I447_093(w_447_093, w_080_389, w_210_020);
  nand2 I447_099(w_447_099, w_271_532, w_201_190);
  nand2 I447_125(w_447_125, w_165_155, w_345_053);
  or2  I447_160(w_447_160, w_355_405, w_340_030);
  or2  I447_173(w_447_173, w_119_101, w_258_390);
  not1 I447_336(w_447_336, w_221_225);
  or2  I447_338(w_447_338, w_180_007, w_110_405);
  nand2 I448_104(w_448_104, w_296_132, w_409_049);
  and2 I448_117(w_448_117, w_091_056, w_368_029);
  and2 I448_151(w_448_151, w_239_000, w_182_015);
  and2 I448_161(w_448_161, w_386_473, w_212_067);
  not1 I448_245(w_448_245, w_328_053);
  nand2 I448_260(w_448_260, w_272_009, w_165_012);
  or2  I448_264(w_448_264, w_164_079, w_107_082);
  nand2 I448_283(w_448_283, w_068_194, w_053_042);
  nand2 I449_138(w_449_138, w_058_025, w_183_025);
  nand2 I449_218(w_449_218, w_336_083, w_344_148);
  nand2 I449_261(w_449_261, w_407_070, w_303_078);
  not1 I450_029(w_450_029, w_137_122);
  and2 I450_052(w_450_052, w_004_450, w_395_041);
  nand2 I450_067(w_450_067, w_303_100, w_228_466);
  not1 I450_070(w_450_070, w_449_261);
  or2  I450_103(w_450_103, w_180_024, w_157_054);
  or2  I450_104(w_450_104, w_295_312, w_360_288);
  or2  I450_107(w_450_107, w_347_328, w_418_105);
  and2 I450_175(w_450_175, w_044_450, w_241_030);
  and2 I451_006(w_451_006, w_405_026, w_388_012);
  not1 I451_064(w_451_064, w_124_046);
  or2  I451_105(w_451_105, w_191_275, w_249_150);
  nand2 I451_133(w_451_133, w_251_064, w_319_210);
  or2  I451_217(w_451_217, w_299_261, w_330_279);
  not1 I451_240(w_451_240, w_063_155);
  and2 I452_045(w_452_045, w_097_153, w_288_070);
  and2 I452_112(w_452_112, w_285_460, w_069_259);
  not1 I452_125(w_452_125, w_212_189);
  not1 I452_300(w_452_300, w_313_192);
  and2 I452_341(w_452_341, w_082_191, w_020_118);
  or2  I453_090(w_453_090, w_284_029, w_240_047);
  not1 I453_552(w_453_552, w_270_217);
  nand2 I454_025(w_454_025, w_263_007, w_071_154);
  and2 I454_039(w_454_039, w_010_488, w_008_471);
  and2 I454_064(w_454_064, w_129_348, w_155_197);
  not1 I454_073(w_454_073, w_094_609);
  not1 I454_079(w_454_079, w_239_000);
  nand2 I454_085(w_454_085, w_019_019, w_127_052);
  nand2 I454_111(w_454_111, w_403_120, w_079_058);
  and2 I454_119(w_454_119, w_018_021, w_338_044);
  and2 I454_158(w_454_158, w_130_134, w_353_535);
  and2 I454_305(w_454_305, w_452_045, w_066_493);
  or2  I454_340(w_454_340, w_021_217, w_417_057);
  nand2 I455_026(w_455_026, w_143_018, w_454_064);
  not1 I455_112(w_455_112, w_070_515);
  not1 I455_144(w_455_144, w_191_134);
  not1 I455_172(w_455_172, w_069_033);
  and2 I455_205(w_455_205, w_083_144, w_100_057);
  nand2 I455_418(w_455_418, w_375_178, w_348_101);
  nand2 I456_039(w_456_039, w_269_276, w_157_097);
  or2  I456_127(w_456_127, w_051_023, w_444_101);
  nand2 I456_193(w_456_193, w_389_066, w_416_134);
  or2  I457_002(w_457_002, w_105_169, w_161_460);
  or2  I457_053(w_457_053, w_075_113, w_190_100);
  or2  I457_054(w_457_054, w_112_169, w_168_266);
  and2 I457_089(w_457_089, w_345_216, w_237_131);
  or2  I457_099(w_457_099, w_371_000, w_376_275);
  not1 I457_107(w_457_107, w_367_295);
  nand2 I457_132(w_457_132, w_135_549, w_298_057);
  or2  I457_139(w_457_139, w_439_045, w_247_163);
  and2 I457_154(w_457_154, w_143_068, w_324_035);
  not1 I457_164(w_457_164, w_221_125);
  or2  I458_038(w_458_038, w_450_029, w_400_091);
  or2  I458_060(w_458_060, w_082_079, w_334_340);
  and2 I458_072(w_458_072, w_227_062, w_271_030);
  not1 I459_035(w_459_035, w_455_205);
  not1 I459_109(w_459_109, w_359_047);
  not1 I459_216(w_459_216, w_154_103);
  and2 I460_003(w_460_003, w_019_003, w_397_036);
  nand2 I460_040(w_460_040, w_246_092, w_351_044);
  nand2 I460_089(w_460_089, w_360_383, w_107_220);
  nand2 I460_173(w_460_173, w_447_338, w_084_012);
  or2  I460_233(w_460_233, w_232_503, w_202_111);
  not1 I460_237(w_460_237, w_216_340);
  and2 I461_173(w_461_173, w_163_593, w_366_144);
  and2 I461_637(w_461_637, w_014_082, w_221_190);
  or2  I462_016(w_462_016, w_424_111, w_035_106);
  and2 I462_379(w_462_379, w_002_643, w_009_591);
  nand2 I462_400(w_462_400, w_280_652, w_232_166);
  nand2 I462_524(w_462_524, w_001_029, w_237_074);
  not1 I462_547(w_462_547, w_080_076);
  or2  I463_000(w_463_000, w_087_028, w_010_649);
  not1 I463_029(w_463_029, w_149_041);
  not1 I463_119(w_463_119, w_429_218);
  or2  I463_192(w_463_192, w_079_008, w_157_164);
  not1 I464_118(w_464_118, w_406_022);
  and2 I464_242(w_464_242, w_015_517, w_232_125);
  and2 I464_281(w_464_281, w_151_295, w_349_027);
  not1 I464_299(w_464_299, w_433_444);
  not1 I464_668(w_464_668, w_380_731);
  nand2 I464_676(w_464_676, w_104_310, w_335_033);
  not1 I465_014(w_465_014, w_435_136);
  or2  I465_019(w_465_019, w_212_061, w_100_120);
  not1 I465_165(w_465_165, w_222_032);
  not1 I465_192(w_465_192, w_187_030);
  nand2 I465_208(w_465_208, w_026_174, w_363_009);
  not1 I465_224(w_465_224, w_253_363);
  not1 I465_269(w_465_269, w_046_401);
  not1 I465_332(w_465_332, w_104_291);
  nand2 I466_053(w_466_053, w_197_064, w_255_076);
  not1 I466_066(w_466_066, w_058_379);
  or2  I466_103(w_466_103, w_117_035, w_045_029);
  nand2 I466_136(w_466_136, w_312_238, w_256_477);
  nand2 I466_214(w_466_214, w_033_172, w_116_023);
  or2  I466_296(w_466_296, w_355_072, w_239_000);
  or2  I467_167(w_467_167, w_046_061, w_416_344);
  and2 I467_177(w_467_177, w_411_130, w_363_359);
  or2  I467_181(w_467_181, w_196_040, w_069_254);
  and2 I467_251(w_467_251, w_439_295, w_395_080);
  and2 I467_284(w_467_284, w_170_240, w_234_429);
  or2  I467_367(w_467_367, w_094_286, w_146_305);
  not1 I468_021(w_468_021, w_124_145);
  or2  I468_025(w_468_025, w_315_238, w_448_161);
  not1 I468_035(w_468_035, w_342_477);
  or2  I468_062(w_468_062, w_321_005, w_465_332);
  nand2 I468_070(w_468_070, w_150_393, w_129_168);
  nand2 I468_079(w_468_079, w_185_072, w_157_094);
  or2  I468_090(w_468_090, w_444_022, w_307_036);
  or2  I468_105(w_468_105, w_336_110, w_284_142);
  nand2 I468_137(w_468_137, w_161_133, w_399_137);
  or2  I468_154(w_468_154, w_354_003, w_307_166);
  nand2 I469_024(w_469_024, w_436_564, w_295_188);
  or2  I469_062(w_469_062, w_048_011, w_198_059);
  nand2 I469_069(w_469_069, w_390_054, w_183_039);
  and2 I469_080(w_469_080, w_337_020, w_088_044);
  or2  I470_407(w_470_407, w_283_272, w_338_312);
  or2  I470_504(w_470_504, w_382_341, w_298_090);
  and2 I471_074(w_471_074, w_150_239, w_232_479);
  or2  I471_169(w_471_169, w_320_411, w_307_391);
  not1 I471_190(w_471_190, w_448_151);
  nand2 I472_163(w_472_163, w_029_063, w_013_021);
  not1 I473_502(w_473_502, w_013_137);
  or2  I474_160(w_474_160, w_194_098, w_318_000);
  and2 I474_202(w_474_202, w_219_636, w_126_061);
  and2 I474_307(w_474_307, w_192_031, w_162_003);
  nand2 I475_011(w_475_011, w_069_096, w_128_495);
  not1 I475_057(w_475_057, w_463_000);
  not1 I475_190(w_475_190, w_433_120);
  and2 I475_193(w_475_193, w_205_034, w_338_264);
  nand2 I475_293(w_475_293, w_093_270, w_146_297);
  not1 I475_296(w_475_296, w_441_144);
  nand2 I475_511(w_475_511, w_145_038, w_134_292);
  or2  I476_235(w_476_235, w_349_289, w_463_029);
  and2 I476_274(w_476_274, w_274_104, w_058_416);
  not1 I476_513(w_476_513, w_124_025);
  or2  I477_022(w_477_022, w_127_053, w_242_093);
  nand2 I477_030(w_477_030, w_018_027, w_110_154);
  or2  I477_032(w_477_032, w_143_088, w_347_109);
  not1 I477_034(w_477_034, w_420_574);
  and2 I477_041(w_477_041, w_237_000, w_326_042);
  and2 I477_057(w_477_057, w_048_006, w_210_098);
  not1 I477_070(w_477_070, w_141_151);
  not1 I478_078(w_478_078, w_173_030);
  and2 I478_177(w_478_177, w_157_031, w_315_111);
  and2 I478_275(w_478_275, w_454_085, w_055_061);
  and2 I478_335(w_478_335, w_180_010, w_317_090);
  or2  I478_381(w_478_381, w_156_242, w_056_629);
  and2 I479_034(w_479_034, w_055_316, w_347_167);
  and2 I479_072(w_479_072, w_083_023, w_022_076);
  and2 I479_088(w_479_088, w_337_101, w_136_017);
  not1 I479_107(w_479_107, w_074_233);
  not1 I479_169(w_479_169, w_080_192);
  not1 I479_185(w_479_185, w_166_322);
  or2  I479_281(w_479_281, w_045_305, w_191_336);
  and2 I479_314(w_479_314, w_061_306, w_379_182);
  nand2 I479_325(w_479_325, w_365_199, w_118_012);
  or2  I480_029(w_480_029, w_373_327, w_229_041);
  nand2 I480_046(w_480_046, w_383_394, w_132_012);
  and2 I480_057(w_480_057, w_308_095, w_265_641);
  or2  I480_075(w_480_075, w_479_169, w_100_060);
  or2  I480_078(w_480_078, w_219_067, w_385_227);
  not1 I480_102(w_480_102, w_074_182);
  nand2 I480_107(w_480_107, w_113_348, w_005_240);
  nand2 I481_039(w_481_039, w_144_044, w_261_061);
  and2 I481_042(w_481_042, w_313_008, w_001_012);
  not1 I481_050(w_481_050, w_255_078);
  nand2 I481_054(w_481_054, w_218_660, w_376_138);
  not1 I481_057(w_481_057, w_007_309);
  and2 I481_058(w_481_058, w_140_155, w_360_269);
  or2  I481_104(w_481_104, w_192_017, w_421_052);
  and2 I481_198(w_481_198, w_242_058, w_009_525);
  or2  I481_215(w_481_215, w_239_000, w_327_155);
  or2  I481_280(w_481_280, w_395_029, w_134_089);
  and2 I482_003(w_482_003, w_349_305, w_413_029);
  not1 I482_077(w_482_077, w_304_223);
  not1 I482_175(w_482_175, w_205_453);
  or2  I482_287(w_482_287, w_179_423, w_174_001);
  not1 I482_327(w_482_327, w_223_016);
  and2 I482_434(w_482_434, w_205_122, w_191_045);
  and2 I483_358(w_483_358, w_446_577, w_139_014);
  not1 I483_428(w_483_428, w_406_050);
  nand2 I483_777(w_483_777, w_390_173, w_165_017);
  not1 I484_008(w_484_008, w_316_246);
  or2  I484_249(w_484_249, w_481_058, w_085_173);
  not1 I484_277(w_484_277, w_452_341);
  and2 I484_296(w_484_296, w_096_001, w_060_085);
  not1 I484_326(w_484_326, w_205_309);
  nand2 I484_329(w_484_329, w_050_106, w_278_116);
  not1 I484_346(w_484_346, w_274_029);
  or2  I484_349(w_484_349, w_246_593, w_138_231);
  and2 I484_379(w_484_379, w_116_495, w_004_462);
  not1 I485_072(w_485_072, w_416_325);
  or2  I485_143(w_485_143, w_468_062, w_132_196);
  and2 I486_038(w_486_038, w_115_241, w_447_099);
  nand2 I486_111(w_486_111, w_179_721, w_294_074);
  or2  I487_002(w_487_002, w_175_038, w_183_111);
  not1 I487_101(w_487_101, w_119_018);
  or2  I487_127(w_487_127, w_326_035, w_164_241);
  and2 I487_141(w_487_141, w_432_307, w_131_071);
  or2  I487_319(w_487_319, w_378_046, w_399_297);
  and2 I487_510(w_487_510, w_124_096, w_308_008);
  not1 I488_017(w_488_017, w_155_045);
  not1 I488_018(w_488_018, w_191_240);
  and2 I488_021(w_488_021, w_016_007, w_110_139);
  and2 I488_037(w_488_037, w_285_011, w_176_129);
  or2  I488_045(w_488_045, w_334_337, w_235_177);
  and2 I488_102(w_488_102, w_416_427, w_477_032);
  or2  I489_025(w_489_025, w_247_162, w_377_087);
  or2  I489_094(w_489_094, w_291_007, w_199_373);
  not1 I489_384(w_489_384, w_172_005);
  not1 I489_395(w_489_395, w_192_114);
  and2 I490_012(w_490_012, w_335_098, w_230_157);
  not1 I490_019(w_490_019, w_153_044);
  or2  I490_067(w_490_067, w_053_054, w_084_014);
  or2  I490_089(w_490_089, w_456_193, w_244_229);
  not1 I490_093(w_490_093, w_365_128);
  not1 I491_021(w_491_021, w_461_637);
  or2  I491_022(w_491_022, w_062_517, w_146_323);
  and2 I491_040(w_491_040, w_223_079, w_067_146);
  or2  I491_077(w_491_077, w_295_227, w_306_106);
  nand2 I492_157(w_492_157, w_408_005, w_096_001);
  and2 I492_275(w_492_275, w_224_095, w_323_269);
  or2  I492_319(w_492_319, w_420_161, w_274_221);
  and2 I492_323(w_492_323, w_184_007, w_339_008);
  nand2 I493_026(w_493_026, w_487_319, w_397_141);
  and2 I493_038(w_493_038, w_258_411, w_316_219);
  and2 I493_044(w_493_044, w_328_153, w_141_093);
  not1 I493_050(w_493_050, w_043_026);
  not1 I493_093(w_493_093, w_066_405);
  not1 I493_095(w_493_095, w_464_281);
  or2  I493_103(w_493_103, w_455_172, w_379_186);
  nand2 I493_139(w_493_139, w_168_028, w_402_068);
  and2 I494_028(w_494_028, w_096_005, w_005_103);
  and2 I494_046(w_494_046, w_186_440, w_262_381);
  or2  I494_241(w_494_241, w_061_184, w_280_258);
  or2  I495_026(w_495_026, w_430_484, w_217_074);
  and2 I495_096(w_495_096, w_042_279, w_171_162);
  and2 I495_128(w_495_128, w_467_251, w_177_006);
  not1 I495_164(w_495_164, w_481_039);
  and2 I495_183(w_495_183, w_014_256, w_033_391);
  and2 I495_343(w_495_343, w_285_041, w_386_188);
  nand2 I495_435(w_495_435, w_091_109, w_092_162);
  or2  I496_077(w_496_077, w_253_008, w_457_107);
  or2  I496_447(w_496_447, w_474_307, w_030_319);
  nand2 I496_598(w_496_600, w_496_599, w_052_000);
  and2 I496_599(w_496_601, w_496_600, w_405_071);
  and2 I496_600(w_496_602, w_496_601, w_328_110);
  and2 I496_601(w_496_603, w_260_159, w_496_602);
  and2 I496_602(w_496_604, w_496_603, w_004_408);
  and2 I496_603(w_496_599, w_496_604, w_450_070);
  not1 I497_078(w_497_078, w_127_071);
  and2 I497_107(w_497_107, w_066_335, w_049_033);
  or2  I498_120(w_498_120, w_085_141, w_240_090);
  or2  I498_170(w_498_170, w_124_001, w_023_200);
  not1 I498_415(w_498_415, w_279_253);
  not1 I498_619(w_498_619, w_238_189);
  nand2 I499_189(w_499_189, w_101_020, w_468_025);
  nand2 I499_222(w_499_222, w_371_000, w_343_138);
  or2  I499_376(w_499_376, w_133_313, w_319_278);
  nand2 I499_433(w_499_433, w_215_533, w_180_001);
  not1 I499_548(w_499_548, w_113_049);
  not1 I499_573(w_499_573, w_134_474);
  and2 I499_583(w_499_583, w_446_298, w_480_075);
  nand2 I500_020(w_500_020, w_360_482, w_016_006);
  and2 I500_064(w_500_064, w_260_058, w_397_046);
  not1 I500_175(w_500_175, w_301_002);
  and2 I500_203(w_500_203, w_339_029, w_446_151);
  not1 I500_226(w_500_226, w_382_046);
  or2  I500_274(w_500_274, w_124_096, w_248_039);
  nand2 I500_302(w_500_302, w_257_075, w_165_051);
  or2  I500_353(w_500_353, w_030_016, w_180_002);
  and2 I501_013(w_501_013, w_163_078, w_183_244);
  nand2 I501_030(w_501_030, w_418_091, w_006_176);
  nand2 I502_349(w_502_349, w_117_016, w_376_251);
  and2 I502_372(w_502_372, w_156_005, w_394_070);
  or2  I502_416(w_502_416, w_188_225, w_370_020);
  nand2 I502_472(w_502_472, w_158_003, w_457_053);
  nand2 I502_539(w_502_539, w_086_201, w_351_336);
  not1 I502_661(w_502_663, w_502_662);
  or2  I502_662(w_502_664, w_461_173, w_502_663);
  and2 I502_663(w_502_665, w_502_664, w_129_353);
  and2 I502_664(w_502_666, w_502_665, w_026_310);
  and2 I502_665(w_502_667, w_050_010, w_502_666);
  or2  I502_666(w_502_662, w_502_682, w_502_667);
  or2  I502_667(w_502_672, w_502_671, w_226_475);
  or2  I502_668(w_502_673, w_502_672, w_500_175);
  not1 I502_669(w_502_674, w_502_673);
  not1 I502_670(w_502_675, w_502_674);
  nand2 I502_671(w_502_676, w_502_675, w_103_002);
  and2 I502_672(w_502_677, w_502_676, w_043_010);
  nand2 I502_673(w_502_678, w_178_006, w_502_677);
  or2  I502_674(w_502_679, w_063_519, w_502_678);
  and2 I502_675(w_502_680, w_408_005, w_502_679);
  not1 I502_676(w_502_671, w_502_662);
  and2 I502_677(w_502_682, w_133_003, w_502_680);
  and2 I502_678(w_502_685, w_362_019, w_502_684);
  or2  I502_679(w_502_686, w_007_173, w_502_685);
  or2  I502_680(w_502_687, w_502_686, w_070_035);
  nand2 I502_681(w_502_688, w_502_703, w_502_687);
  and2 I502_682(w_502_689, w_151_215, w_502_688);
  and2 I502_683(w_502_690, w_502_689, w_124_281);
  not1 I502_684(w_502_691, w_502_690);
  and2 I502_685(w_502_692, w_238_264, w_502_691);
  or2  I502_686(w_502_684, w_502_692, w_356_044);
  nand2 I502_687(w_502_697, w_008_302, w_502_696);
  nand2 I502_688(w_502_698, w_502_697, w_248_099);
  and2 I502_689(w_502_699, w_502_698, w_006_165);
  and2 I502_690(w_502_700, w_502_699, w_075_153);
  and2 I502_691(w_502_701, w_502_700, w_198_076);
  not1 I502_692(w_502_696, w_502_688);
  and2 I502_693(w_502_703, w_237_084, w_502_701);
  and2 I503_015(w_503_015, w_301_046, w_225_194);
  or2  I503_190(w_503_190, w_301_153, w_251_047);
  not1 I503_202(w_503_202, w_218_334);
  or2  I503_252(w_503_252, w_389_087, w_026_117);
  not1 I503_483(w_503_484, w_503_483);
  nand2 I503_484(w_503_485, w_503_484, w_146_168);
  and2 I503_485(w_503_486, w_439_039, w_503_485);
  or2  I503_486(w_503_487, w_159_018, w_503_486);
  and2 I503_487(w_503_488, w_503_487, w_047_249);
  not1 I503_488(w_503_489, w_503_488);
  not1 I503_489(w_503_490, w_503_489);
  nand2 I503_490(w_503_491, w_407_133, w_503_490);
  and2 I503_491(w_503_492, w_503_491, w_414_325);
  not1 I503_492(w_503_483, w_503_492);
  or2  I504_027(w_504_027, w_256_097, w_363_056);
  or2  I504_031(w_504_031, w_110_289, w_182_026);
  and2 I504_053(w_504_053, w_487_141, w_497_078);
  nand2 I505_066(w_505_066, w_294_046, w_274_143);
  nand2 I505_074(w_505_074, w_222_226, w_038_531);
  and2 I505_236(w_505_236, w_409_153, w_397_137);
  and2 I506_071(w_506_071, w_124_171, w_130_023);
  nand2 I506_153(w_506_153, w_428_010, w_182_009);
  and2 I506_261(w_506_261, w_435_085, w_404_588);
  not1 I506_513(w_506_513, w_253_060);
  nand2 I506_594(w_506_594, w_425_214, w_150_200);
  or2  I506_611(w_506_611, w_477_034, w_179_044);
  or2  I506_631(w_506_633, w_506_632, w_191_082);
  and2 I506_632(w_506_634, w_506_633, w_266_324);
  or2  I506_633(w_506_632, w_506_634, w_506_644);
  or2  I506_634(w_506_639, w_309_215, w_506_638);
  or2  I506_635(w_506_640, w_506_639, w_249_280);
  and2 I506_636(w_506_641, w_506_640, w_168_315);
  and2 I506_637(w_506_642, w_506_641, w_137_185);
  not1 I506_638(w_506_638, w_506_632);
  and2 I506_639(w_506_644, w_447_093, w_506_642);
  nand2 I507_012(w_507_012, w_275_090, w_393_102);
  or2  I507_016(w_507_016, w_028_222, w_239_000);
  not1 I507_035(w_507_035, w_110_290);
  nand2 I507_046(w_507_046, w_342_217, w_022_185);
  nand2 I508_005(w_508_005, w_333_222, w_267_055);
  nand2 I508_074(w_508_074, w_002_237, w_019_019);
  or2  I508_172(w_508_172, w_330_116, w_036_097);
  nand2 I508_173(w_508_173, w_130_252, w_464_668);
  and2 I508_396(w_508_396, w_161_272, w_263_101);
  not1 I509_075(w_509_075, w_440_037);
  not1 I509_086(w_509_088, w_509_087);
  and2 I509_087(w_509_089, w_382_563, w_509_088);
  or2  I509_088(w_509_090, w_509_104, w_509_089);
  not1 I509_089(w_509_091, w_509_090);
  and2 I509_090(w_509_092, w_509_091, w_467_367);
  and2 I509_091(w_509_087, w_509_092, w_172_042);
  not1 I509_092(w_509_097, w_509_096);
  nand2 I509_093(w_509_098, w_509_097, w_265_237);
  and2 I509_094(w_509_099, w_141_044, w_509_098);
  not1 I509_095(w_509_100, w_509_099);
  or2  I509_096(w_509_101, w_509_100, w_107_211);
  and2 I509_097(w_509_102, w_509_101, w_016_006);
  not1 I509_098(w_509_096, w_509_090);
  and2 I509_099(w_509_104, w_191_074, w_509_102);
  not1 I510_136(w_510_136, w_102_597);
  not1 I510_292(w_510_292, w_159_037);
  nand2 I510_447(w_510_447, w_458_038, w_103_156);
  or2  I510_595(w_510_595, w_408_004, w_017_086);
  and2 I510_748(w_510_748, w_246_482, w_332_224);
  or2  I511_028(w_511_028, w_158_002, w_011_148);
  or2  I511_186(w_511_186, w_059_184, w_338_022);
  nand2 I511_240(w_511_240, w_159_039, w_435_085);
  nand2 I511_326(w_511_326, w_069_003, w_468_137);
  and2 I511_396(w_511_396, w_370_095, w_367_125);
  nand2 I512_059(w_512_059, w_357_460, w_322_013);
  not1 I512_088(w_512_088, w_174_066);
  and2 I512_098(w_512_098, w_292_554, w_075_065);
  and2 I512_124(w_512_124, w_080_287, w_224_083);
  and2 I512_157(w_512_157, w_228_146, w_423_052);
  and2 I512_434(w_512_434, w_129_313, w_059_060);
  nand2 I512_451(w_512_451, w_361_221, w_200_106);
  and2 I513_076(w_513_076, w_252_280, w_214_206);
  nand2 I513_232(w_513_232, w_241_029, w_047_007);
  not1 I513_378(w_513_378, w_176_158);
  nand2 I513_448(w_513_448, w_208_354, w_384_046);
  or2  I513_499(w_513_499, w_172_046, w_420_587);
  not1 I513_576(w_513_576, w_254_000);
  not1 I514_083(w_514_083, w_073_245);
  nand2 I514_170(w_514_170, w_475_190, w_068_009);
  or2  I514_191(w_514_191, w_234_111, w_430_092);
  not1 I514_456(w_514_456, w_017_399);
  and2 I515_066(w_515_066, w_500_020, w_140_092);
  nand2 I515_094(w_515_094, w_168_126, w_054_590);
  not1 I515_172(w_515_172, w_401_178);
  and2 I515_371(w_515_371, w_000_485, w_482_434);
  or2  I516_079(w_516_079, w_508_172, w_448_264);
  not1 I516_096(w_516_096, w_480_102);
  or2  I516_329(w_516_329, w_161_446, w_247_159);
  or2  I516_406(w_516_406, w_338_003, w_282_298);
  and2 I517_005(w_517_005, w_195_006, w_230_060);
  or2  I517_052(w_517_052, w_499_433, w_046_120);
  nand2 I517_098(w_517_098, w_227_163, w_002_535);
  not1 I517_227(w_517_227, w_284_005);
  nand2 I518_010(w_518_010, w_097_201, w_510_292);
  nand2 I518_057(w_518_057, w_315_724, w_145_066);
  nand2 I518_062(w_518_062, w_457_089, w_132_384);
  or2  I519_022(w_519_022, w_507_046, w_308_155);
  and2 I519_041(w_519_041, w_021_117, w_166_081);
  or2  I520_053(w_520_053, w_454_119, w_294_009);
  nand2 I520_109(w_520_109, w_051_162, w_039_117);
  not1 I520_202(w_520_202, w_354_113);
  and2 I520_253(w_520_253, w_059_288, w_154_110);
  not1 I520_292(w_520_294, w_520_293);
  and2 I520_293(w_520_295, w_520_294, w_520_305);
  not1 I520_294(w_520_293, w_520_295);
  nand2 I520_295(w_520_300, w_520_299, w_422_008);
  nand2 I520_296(w_520_301, w_520_300, w_215_434);
  or2  I520_297(w_520_302, w_187_020, w_520_301);
  and2 I520_298(w_520_303, w_274_149, w_520_302);
  not1 I520_299(w_520_299, w_520_295);
  and2 I520_300(w_520_305, w_011_242, w_520_303);
  nand2 I521_058(w_521_058, w_318_003, w_013_144);
  nand2 I521_151(w_521_151, w_495_183, w_047_399);
  and2 I521_322(w_521_322, w_418_068, w_169_365);
  or2  I521_334(w_521_334, w_213_392, w_478_177);
  and2 I522_092(w_522_092, w_327_344, w_091_153);
  not1 I522_256(w_522_256, w_157_162);
  nand2 I522_397(w_522_397, w_316_257, w_376_176);
  not1 I522_505(w_522_505, w_283_043);
  or2  I522_539(w_522_539, w_229_323, w_417_075);
  not1 I523_003(w_523_003, w_004_046);
  nand2 I523_065(w_523_065, w_433_398, w_449_138);
  or2  I523_087(w_523_087, w_063_424, w_450_104);
  nand2 I523_190(w_523_190, w_254_057, w_199_235);
  and2 I523_473(w_523_473, w_353_570, w_110_237);
  or2  I524_346(w_524_346, w_386_115, w_341_351);
  nand2 I524_444(w_524_444, w_192_059, w_459_109);
  and2 I524_591(w_524_591, w_385_213, w_046_646);
  not1 I524_595(w_524_595, w_390_187);
  not1 I524_612(w_524_612, w_256_484);
  nand2 I525_007(w_525_007, w_036_024, w_512_059);
  not1 I525_029(w_525_029, w_167_078);
  or2  I525_081(w_525_081, w_117_059, w_140_178);
  not1 I525_095(w_525_095, w_096_004);
  or2  I526_153(w_526_153, w_235_046, w_102_035);
  nand2 I527_061(w_527_061, w_071_066, w_226_138);
  and2 I527_082(w_527_082, w_103_140, w_177_310);
  and2 I527_096(w_527_096, w_109_229, w_277_268);
  nand2 I527_197(w_527_197, w_327_363, w_233_204);
  not1 I527_223(w_527_223, w_495_343);
  not1 I527_350(w_527_350, w_479_072);
  not1 I527_526(w_527_526, w_195_236);
  and2 I528_015(w_528_015, w_145_032, w_442_045);
  or2  I528_017(w_528_017, w_325_238, w_104_067);
  and2 I528_039(w_528_039, w_289_574, w_366_174);
  and2 I528_046(w_528_046, w_488_017, w_394_107);
  or2  I529_000(w_529_000, w_284_102, w_086_185);
  not1 I529_002(w_529_002, w_522_256);
  nand2 I529_004(w_529_004, w_016_007, w_408_004);
  nand2 I530_042(w_530_042, w_259_457, w_122_103);
  nand2 I530_096(w_530_096, w_155_001, w_051_106);
  not1 I530_147(w_530_147, w_031_601);
  and2 I530_182(w_530_182, w_325_000, w_235_141);
  and2 I530_219(w_530_219, w_108_031, w_047_342);
  or2  I531_012(w_531_012, w_369_524, w_351_095);
  and2 I531_317(w_531_317, w_496_447, w_348_114);
  nand2 I531_580(w_531_580, w_084_001, w_123_101);
  nand2 I532_176(w_532_176, w_106_032, w_307_093);
  or2  I532_222(w_532_222, w_102_199, w_069_140);
  nand2 I532_242(w_532_244, w_532_243, w_206_119);
  not1 I532_243(w_532_245, w_532_244);
  and2 I532_244(w_532_246, w_532_245, w_360_353);
  or2  I532_245(w_532_247, w_532_246, w_422_005);
  not1 I532_246(w_532_248, w_532_247);
  or2  I532_247(w_532_249, w_532_248, w_282_387);
  not1 I532_248(w_532_250, w_532_249);
  not1 I532_249(w_532_251, w_532_250);
  not1 I532_250(w_532_252, w_532_251);
  nand2 I532_251(w_532_253, w_532_252, w_306_281);
  and2 I532_252(w_532_254, w_532_266, w_532_253);
  and2 I532_253(w_532_243, w_532_254, w_082_502);
  or2  I532_254(w_532_259, w_165_109, w_532_258);
  nand2 I532_255(w_532_260, w_291_123, w_532_259);
  not1 I532_256(w_532_261, w_532_260);
  or2  I532_257(w_532_262, w_481_054, w_532_261);
  and2 I532_258(w_532_263, w_477_041, w_532_262);
  and2 I532_259(w_532_264, w_078_520, w_532_263);
  not1 I532_260(w_532_258, w_532_254);
  and2 I532_261(w_532_266, w_103_149, w_532_264);
  or2  I533_089(w_533_089, w_254_037, w_529_004);
  or2  I533_110(w_533_110, w_405_132, w_057_121);
  or2  I533_169(w_533_169, w_114_189, w_024_342);
  or2  I533_187(w_533_187, w_030_348, w_354_048);
  nand2 I533_253(w_533_253, w_460_040, w_070_044);
  and2 I533_329(w_533_329, w_359_075, w_107_396);
  nand2 I533_361(w_533_361, w_422_013, w_233_037);
  nand2 I533_532(w_533_532, w_320_218, w_201_268);
  not1 I533_550(w_533_550, w_446_438);
  and2 I534_003(w_534_003, w_224_113, w_211_023);
  and2 I534_011(w_534_011, w_152_200, w_294_019);
  and2 I534_016(w_534_018, w_534_017, w_073_516);
  nand2 I534_017(w_534_019, w_481_198, w_534_018);
  and2 I534_018(w_534_020, w_109_407, w_534_019);
  nand2 I534_019(w_534_021, w_058_562, w_534_020);
  or2  I534_020(w_534_022, w_534_021, w_468_105);
  nand2 I534_021(w_534_023, w_534_022, w_150_378);
  and2 I534_022(w_534_024, w_534_023, w_161_183);
  nand2 I534_023(w_534_017, w_327_364, w_534_024);
  not1 I535_000(w_535_000, w_186_131);
  or2  I535_114(w_535_114, w_071_299, w_205_217);
  not1 I535_119(w_535_119, w_122_094);
  or2  I535_180(w_535_180, w_157_058, w_189_463);
  not1 I535_189(w_535_189, w_142_205);
  or2  I535_202(w_535_202, w_120_343, w_350_049);
  nand2 I535_252(w_535_252, w_261_034, w_522_539);
  and2 I535_261(w_535_263, w_535_262, w_235_115);
  and2 I535_262(w_535_264, w_535_263, w_389_279);
  not1 I535_263(w_535_265, w_535_264);
  and2 I535_264(w_535_266, w_343_478, w_535_265);
  nand2 I535_265(w_535_267, w_535_266, w_471_190);
  or2  I535_266(w_535_268, w_351_240, w_535_267);
  and2 I535_267(w_535_269, w_535_278, w_535_268);
  and2 I535_268(w_535_262, w_535_269, w_481_280);
  nand2 I535_269(w_535_274, w_321_303, w_535_273);
  and2 I535_270(w_535_275, w_535_274, w_106_023);
  and2 I535_271(w_535_276, w_535_275, w_281_044);
  not1 I535_272(w_535_273, w_535_269);
  and2 I535_273(w_535_278, w_292_433, w_535_276);
  or2  I535_274(w_535_281, w_038_116, w_535_280);
  or2  I535_275(w_535_282, w_475_293, w_535_281);
  not1 I535_276(w_535_283, w_535_282);
  and2 I535_277(w_535_284, w_535_283, w_485_143);
  and2 I535_278(w_535_285, w_403_289, w_535_284);
  not1 I535_279(w_535_286, w_535_285);
  and2 I535_280(w_535_287, w_535_299, w_535_286);
  and2 I535_281(w_535_288, w_434_061, w_535_287);
  or2  I535_282(w_535_280, w_535_288, w_434_335);
  or2  I535_283(w_535_293, w_335_151, w_535_292);
  and2 I535_284(w_535_294, w_535_293, w_176_085);
  nand2 I535_285(w_535_295, w_349_177, w_535_294);
  not1 I535_286(w_535_296, w_535_295);
  and2 I535_287(w_535_297, w_050_470, w_535_296);
  not1 I535_288(w_535_292, w_535_287);
  and2 I535_289(w_535_299, w_401_079, w_535_297);
  or2  I536_022(w_536_022, w_417_116, w_053_085);
  and2 I536_040(w_536_040, w_025_287, w_516_406);
  nand2 I537_029(w_537_029, w_320_389, w_383_240);
  not1 I537_032(w_537_032, w_163_036);
  not1 I537_053(w_537_053, w_388_100);
  nand2 I537_056(w_537_056, w_211_028, w_446_533);
  and2 I537_154(w_537_154, w_502_416, w_193_131);
  not1 I537_220(w_537_220, w_080_183);
  and2 I537_248(w_537_248, w_507_012, w_357_302);
  not1 I537_264(w_537_264, w_265_073);
  nand2 I538_039(w_538_039, w_137_003, w_124_143);
  nand2 I538_046(w_538_046, w_080_430, w_334_367);
  nand2 I538_190(w_538_190, w_167_041, w_462_016);
  or2  I538_262(w_538_262, w_438_084, w_169_101);
  or2  I539_321(w_539_321, w_105_327, w_029_104);
  or2  I539_387(w_539_387, w_451_064, w_425_362);
  nand2 I539_388(w_539_388, w_486_038, w_419_139);
  not1 I539_422(w_539_422, w_515_371);
  or2  I539_491(w_539_491, w_301_027, w_146_227);
  or2  I539_538(w_539_538, w_037_081, w_283_064);
  or2  I539_723(w_539_723, w_225_204, w_347_117);
  and2 I540_053(w_540_053, w_205_053, w_086_134);
  or2  I540_118(w_540_118, w_071_145, w_227_160);
  and2 I541_024(w_541_024, w_019_018, w_476_235);
  and2 I541_066(w_541_066, w_471_169, w_137_469);
  nand2 I542_007(w_542_007, w_067_052, w_242_134);
  or2  I542_053(w_542_053, w_262_073, w_409_455);
  nand2 I542_058(w_542_058, w_460_003, w_147_097);
  not1 I542_061(w_542_061, w_429_003);
  nand2 I542_116(w_542_116, w_265_029, w_179_745);
  not1 I542_331(w_542_331, w_478_275);
  and2 I543_105(w_543_105, w_469_080, w_128_111);
  and2 I543_210(w_543_210, w_447_125, w_542_058);
  and2 I543_769(w_543_771, w_543_770, w_370_056);
  nand2 I543_770(w_543_772, w_543_771, w_053_081);
  not1 I543_771(w_543_773, w_543_772);
  and2 I543_772(w_543_774, w_543_788, w_543_773);
  not1 I543_773(w_543_775, w_543_774);
  not1 I543_774(w_543_776, w_543_775);
  and2 I543_775(w_543_777, w_543_776, w_500_302);
  or2  I543_776(w_543_778, w_110_386, w_543_777);
  nand2 I543_777(w_543_779, w_209_322, w_543_778);
  and2 I543_778(w_543_780, w_137_076, w_543_779);
  or2  I543_779(w_543_770, w_383_350, w_543_780);
  or2  I543_780(w_543_785, w_173_030, w_543_784);
  and2 I543_781(w_543_786, w_158_000, w_543_785);
  not1 I543_782(w_543_784, w_543_774);
  and2 I543_783(w_543_788, w_466_136, w_543_786);
  nand2 I544_146(w_544_146, w_175_221, w_404_196);
  nand2 I544_153(w_544_153, w_077_481, w_375_171);
  nand2 I545_117(w_545_117, w_148_215, w_513_232);
  nand2 I545_151(w_545_151, w_181_123, w_314_077);
  nand2 I545_345(w_545_345, w_277_020, w_002_482);
  not1 I545_349(w_545_349, w_274_144);
  not1 I546_073(w_546_073, w_144_010);
  nand2 I546_086(w_546_086, w_445_135, w_376_055);
  not1 I546_385(w_546_385, w_441_407);
  or2  I546_450(w_546_450, w_110_148, w_147_146);
  not1 I546_517(w_546_519, w_546_518);
  not1 I546_518(w_546_520, w_546_519);
  not1 I546_519(w_546_521, w_546_520);
  or2  I546_520(w_546_522, w_546_521, w_305_077);
  not1 I546_521(w_546_523, w_546_522);
  and2 I546_522(w_546_524, w_546_523, w_489_094);
  and2 I546_523(w_546_518, w_475_193, w_546_524);
  nand2 I547_002(w_547_002, w_178_015, w_250_605);
  or2  I547_024(w_547_024, w_167_100, w_295_275);
  or2  I547_031(w_547_031, w_296_129, w_526_153);
  or2  I547_032(w_547_032, w_385_106, w_252_247);
  and2 I547_034(w_547_034, w_065_496, w_401_230);
  or2  I547_035(w_547_035, w_099_169, w_331_111);
  nand2 I547_045(w_547_045, w_049_217, w_237_111);
  not1 I548_060(w_548_060, w_136_013);
  or2  I548_192(w_548_192, w_178_015, w_271_416);
  and2 I548_264(w_548_264, w_074_265, w_489_395);
  nand2 I549_047(w_549_047, w_404_648, w_167_108);
  and2 I549_107(w_549_107, w_450_107, w_358_066);
  not1 I549_130(w_549_130, w_444_520);
  and2 I550_122(w_550_122, w_238_052, w_120_038);
  not1 I550_260(w_550_260, w_376_251);
  not1 I551_007(w_551_007, w_211_012);
  or2  I551_012(w_551_012, w_129_023, w_317_249);
  or2  I551_031(w_551_031, w_119_043, w_196_141);
  nand2 I551_088(w_551_088, w_308_107, w_513_378);
  or2  I551_109(w_551_109, w_200_282, w_176_059);
  nand2 I552_006(w_552_006, w_098_011, w_302_338);
  and2 I552_100(w_552_100, w_366_238, w_337_072);
  and2 I552_304(w_552_304, w_267_131, w_205_367);
  not1 I553_015(w_553_015, w_468_021);
  or2  I553_020(w_553_020, w_455_418, w_271_072);
  and2 I553_027(w_553_027, w_492_157, w_161_134);
  or2  I553_031(w_553_031, w_338_010, w_436_562);
  not1 I554_069(w_554_069, w_322_022);
  nand2 I555_067(w_555_067, w_220_119, w_169_380);
  or2  I555_293(w_555_293, w_529_002, w_387_252);
  and2 I556_035(w_556_035, w_240_101, w_252_394);
  not1 I556_212(w_556_212, w_079_024);
  or2  I556_270(w_556_270, w_544_153, w_399_163);
  nand2 I556_324(w_556_324, w_029_106, w_170_198);
  or2  I556_463(w_556_463, w_386_161, w_122_022);
  nand2 I557_047(w_557_047, w_040_601, w_465_208);
  nand2 I557_050(w_557_050, w_439_038, w_510_595);
  or2  I557_062(w_557_062, w_229_136, w_419_308);
  nand2 I557_111(w_557_111, w_495_026, w_325_272);
  nand2 I557_167(w_557_167, w_523_473, w_524_444);
  or2  I557_419(w_557_419, w_479_314, w_013_088);
  and2 I557_428(w_557_430, w_415_079, w_557_429);
  not1 I557_429(w_557_431, w_557_430);
  and2 I557_430(w_557_432, w_315_171, w_557_431);
  nand2 I557_431(w_557_429, w_557_432, w_330_247);
  or2  I558_030(w_558_030, w_075_152, w_477_022);
  not1 I558_122(w_558_122, w_495_435);
  or2  I558_151(w_558_151, w_170_423, w_343_605);
  nand2 I559_020(w_559_020, w_129_088, w_385_427);
  or2  I559_028(w_559_028, w_029_061, w_044_030);
  and2 I559_040(w_559_040, w_020_518, w_459_035);
  nand2 I560_071(w_560_071, w_523_065, w_455_026);
  or2  I560_106(w_560_106, w_074_105, w_021_098);
  nand2 I560_149(w_560_149, w_488_102, w_525_081);
  and2 I560_512(w_560_512, w_518_057, w_015_461);
  not1 I560_543(w_560_543, w_383_112);
  or2  I561_038(w_561_038, w_315_524, w_452_112);
  and2 I561_079(w_561_079, w_001_035, w_199_106);
  or2  I561_175(w_561_175, w_031_001, w_163_486);
  not1 I561_205(w_561_205, w_396_045);
  and2 I561_308(w_561_308, w_501_030, w_138_096);
  not1 I561_343(w_561_343, w_537_053);
  not1 I562_147(w_562_147, w_151_009);
  or2  I562_429(w_562_429, w_451_133, w_276_110);
  and2 I562_660(w_562_660, w_294_110, w_162_020);
  or2  I563_022(w_563_022, w_273_075, w_191_331);
  nand2 I563_052(w_563_052, w_548_192, w_157_121);
  and2 I563_470(w_563_470, w_464_676, w_101_104);
  or2  I564_007(w_564_007, w_440_064, w_132_435);
  or2  I564_065(w_564_065, w_208_169, w_177_288);
  not1 I564_097(w_564_097, w_165_071);
  nand2 I564_279(w_564_281, w_564_280, w_467_167);
  and2 I564_280(w_564_282, w_564_281, w_440_079);
  not1 I564_281(w_564_283, w_564_282);
  or2  I564_282(w_564_284, w_564_283, w_193_296);
  nand2 I564_283(w_564_285, w_446_406, w_564_284);
  and2 I564_284(w_564_286, w_480_046, w_564_285);
  and2 I564_285(w_564_287, w_564_286, w_240_038);
  or2  I564_286(w_564_288, w_564_287, w_367_160);
  and2 I564_287(w_564_289, w_418_045, w_564_288);
  not1 I564_288(w_564_290, w_564_289);
  and2 I564_289(w_564_291, w_564_290, w_205_000);
  not1 I564_290(w_564_280, w_564_291);
  and2 I565_008(w_565_008, w_088_121, w_484_008);
  not1 I565_009(w_565_009, w_506_153);
  not1 I565_020(w_565_020, w_328_037);
  nand2 I566_094(w_566_094, w_450_103, w_151_276);
  and2 I566_198(w_566_198, w_299_316, w_029_085);
  not1 I567_003(w_567_003, w_556_463);
  or2  I567_010(w_567_010, w_495_128, w_171_228);
  and2 I567_014(w_567_014, w_528_017, w_274_126);
  not1 I567_016(w_567_016, w_564_097);
  or2  I567_020(w_567_020, w_391_100, w_547_034);
  or2  I567_033(w_567_033, w_445_021, w_344_042);
  or2  I567_040(w_567_040, w_476_513, w_420_673);
  or2  I567_042(w_567_042, w_269_565, w_385_124);
  or2  I568_227(w_568_227, w_435_075, w_508_173);
  and2 I568_367(w_568_367, w_062_211, w_497_107);
  not1 I568_499(w_568_499, w_189_513);
  nand2 I569_040(w_569_040, w_206_010, w_460_089);
  and2 I569_133(w_569_133, w_127_008, w_193_327);
  not1 I570_085(w_570_085, w_029_039);
  not1 I570_197(w_570_199, w_570_198);
  not1 I570_198(w_570_200, w_570_199);
  not1 I570_199(w_570_201, w_570_200);
  not1 I570_200(w_570_202, w_570_201);
  and2 I570_201(w_570_203, w_570_202, w_310_258);
  and2 I570_202(w_570_204, w_570_203, w_281_119);
  or2  I570_203(w_570_205, w_570_204, w_190_001);
  and2 I570_204(w_570_206, w_570_220, w_570_205);
  nand2 I570_205(w_570_198, w_570_206, w_214_206);
  or2  I570_206(w_570_211, w_570_210, w_307_350);
  not1 I570_207(w_570_212, w_570_211);
  and2 I570_208(w_570_213, w_393_084, w_570_212);
  not1 I570_209(w_570_214, w_570_213);
  not1 I570_210(w_570_215, w_570_214);
  nand2 I570_211(w_570_216, w_366_072, w_570_215);
  nand2 I570_212(w_570_217, w_210_061, w_570_216);
  and2 I570_213(w_570_218, w_242_082, w_570_217);
  not1 I570_214(w_570_210, w_570_206);
  and2 I570_215(w_570_220, w_279_138, w_570_218);
  and2 I571_075(w_571_075, w_152_621, w_409_408);
  not1 I571_130(w_571_130, w_138_024);
  not1 I571_402(w_571_402, w_457_132);
  and2 I571_624(w_570_208, w_479_088, w_570_198);
  or2  I572_107(w_572_107, w_304_258, w_294_017);
  and2 I572_131(w_572_131, w_570_208, w_543_210);
  or2  I572_140(w_572_140, w_542_053, w_432_218);
  nand2 I573_020(w_573_020, w_060_290, w_146_088);
  not1 I573_043(w_573_043, w_172_013);
  not1 I573_058(w_573_058, w_549_130);
  and2 I573_208(w_573_208, w_263_104, w_481_104);
  not1 I573_223(w_573_223, w_558_030);
  or2  I573_324(w_573_324, w_355_038, w_533_253);
  and2 I574_164(w_574_164, w_052_012, w_097_088);
  nand2 I574_265(w_574_265, w_080_407, w_547_024);
  nand2 I574_373(w_574_373, w_163_509, w_134_135);
  nand2 I575_000(w_575_000, w_281_365, w_186_140);
  nand2 I575_053(w_575_053, w_539_422, w_126_116);
  or2  I575_064(w_575_064, w_537_220, w_080_153);
  or2  I575_065(w_575_065, w_123_364, w_271_555);
  or2  I575_094(w_575_094, w_520_253, w_147_100);
  or2  I575_096(w_575_096, w_215_124, w_336_025);
  nand2 I575_160(w_575_160, w_439_313, w_183_092);
  or2  I575_178(w_575_178, w_090_066, w_309_187);
  or2  I575_207(w_575_207, w_158_000, w_268_152);
  not1 I576_111(w_576_111, w_135_191);
  nand2 I576_172(w_576_172, w_019_001, w_393_109);
  and2 I576_288(w_576_290, w_139_020, w_576_289);
  and2 I576_289(w_576_291, w_576_290, w_457_139);
  nand2 I576_290(w_576_292, w_134_323, w_576_291);
  nand2 I576_291(w_576_293, w_492_323, w_576_292);
  and2 I576_292(w_576_294, w_576_293, w_375_142);
  and2 I576_293(w_576_295, w_576_294, w_453_090);
  or2  I576_294(w_576_296, w_173_013, w_576_295);
  not1 I576_295(w_576_297, w_576_296);
  and2 I576_296(w_576_298, w_576_297, w_547_032);
  nand2 I576_297(w_576_289, w_341_035, w_576_298);
  and2 I577_031(w_577_031, w_025_171, w_537_248);
  or2  I577_485(w_577_485, w_011_324, w_454_158);
  or2  I577_496(w_577_496, w_340_004, w_551_109);
  and2 I578_007(w_578_007, w_126_142, w_032_352);
  nand2 I578_284(w_578_284, w_023_023, w_044_657);
  or2  I578_543(w_578_543, w_165_050, w_152_387);
  or2  I578_724(w_578_724, w_466_214, w_546_385);
  and2 I579_358(w_579_358, w_047_327, w_388_025);
  nand2 I579_461(w_579_461, w_068_328, w_388_159);
  not1 I579_647(w_579_647, w_180_012);
  nand2 I580_031(w_580_031, w_093_016, w_230_233);
  and2 I580_420(w_580_420, w_304_500, w_487_127);
  nand2 I581_400(w_581_400, w_551_109, w_482_287);
  or2  I582_245(w_582_245, w_053_115, w_194_077);
  not1 I582_461(w_582_461, w_379_071);
  not1 I582_657(w_582_657, w_279_124);
  nand2 I582_708(w_582_708, w_074_194, w_263_119);
  nand2 I583_002(w_583_002, w_005_260, w_551_088);
  nand2 I583_023(w_583_023, w_037_309, w_567_016);
  not1 I583_075(w_583_075, w_470_504);
  or2  I583_099(w_583_101, w_583_100, w_583_117);
  and2 I583_100(w_583_102, w_583_101, w_048_007);
  and2 I583_101(w_583_100, w_583_102, w_125_084);
  or2  I583_102(w_583_107, w_321_282, w_583_106);
  nand2 I583_103(w_583_108, w_583_107, w_287_315);
  or2  I583_104(w_583_109, w_583_108, w_259_472);
  nand2 I583_105(w_583_110, w_437_010, w_583_109);
  nand2 I583_106(w_583_111, w_373_057, w_583_110);
  and2 I583_107(w_583_112, w_583_111, w_103_048);
  not1 I583_108(w_583_113, w_583_112);
  not1 I583_109(w_583_114, w_583_113);
  and2 I583_110(w_583_115, w_103_137, w_583_114);
  not1 I583_111(w_583_106, w_583_101);
  and2 I583_112(w_583_117, w_219_656, w_583_115);
  nand2 I584_024(w_584_024, w_191_136, w_332_261);
  nand2 I584_255(w_584_255, w_395_290, w_361_070);
  or2  I584_341(w_584_341, w_195_209, w_317_264);
  not1 I584_544(w_584_544, w_201_062);
  or2  I584_574(w_584_574, w_170_226, w_308_022);
  nand2 I584_666(w_584_666, w_478_381, w_458_072);
  not1 I584_712(w_584_712, w_200_407);
  or2  I585_046(w_585_046, w_128_130, w_134_002);
  nand2 I585_101(w_585_101, w_220_195, w_364_027);
  or2  I585_554(w_585_554, w_293_325, w_567_020);
  or2  I585_731(w_585_733, w_565_008, w_585_732);
  nand2 I585_732(w_585_734, w_585_753, w_585_733);
  or2  I585_733(w_585_735, w_585_734, w_511_326);
  or2  I585_734(w_585_736, w_177_102, w_585_735);
  not1 I585_735(w_585_737, w_585_736);
  and2 I585_736(w_585_738, w_079_052, w_585_737);
  not1 I585_737(w_585_732, w_585_738);
  and2 I585_738(w_585_743, w_585_742, w_430_422);
  nand2 I585_739(w_585_744, w_291_129, w_585_743);
  and2 I585_740(w_585_745, w_260_282, w_585_744);
  not1 I585_741(w_585_746, w_585_745);
  and2 I585_742(w_585_747, w_585_746, w_295_308);
  and2 I585_743(w_585_748, w_585_747, w_530_182);
  or2  I585_744(w_585_749, w_460_237, w_585_748);
  and2 I585_745(w_585_750, w_585_749, w_532_176);
  and2 I585_746(w_585_751, w_585_750, w_332_451);
  not1 I585_747(w_585_742, w_585_734);
  and2 I585_748(w_585_753, w_378_111, w_585_751);
  nand2 I585_749(w_585_756, w_263_028, w_585_755);
  nand2 I585_750(w_585_757, w_459_216, w_585_756);
  not1 I585_751(w_585_758, w_585_757);
  not1 I585_752(w_585_759, w_585_758);
  nand2 I585_753(w_585_760, w_585_759, w_281_307);
  or2  I585_754(w_585_761, w_562_660, w_585_760);
  and2 I585_755(w_585_762, w_585_761, w_171_611);
  nand2 I585_756(w_585_763, w_585_762, w_166_288);
  and2 I585_757(w_585_764, w_585_763, w_522_092);
  and2 I585_758(w_585_765, w_513_448, w_585_764);
  and2 I585_759(w_585_766, w_120_222, w_585_765);
  or2  I585_760(w_585_755, w_585_766, w_002_397);
  or2  I586_040(w_586_040, w_436_218, w_415_046);
  not1 I586_073(w_586_073, w_311_288);
  nand2 I586_090(w_586_090, w_417_060, w_045_269);
  nand2 I586_096(w_586_096, w_210_132, w_356_078);
  or2  I586_125(w_586_125, w_264_310, w_195_072);
  or2  I586_230(w_586_231, w_586_230, w_421_047);
  or2  I586_231(w_586_232, w_582_657, w_586_231);
  and2 I586_232(w_586_233, w_165_007, w_586_232);
  not1 I586_233(w_586_234, w_586_233);
  not1 I586_234(w_586_235, w_586_234);
  and2 I586_235(w_586_236, w_051_244, w_586_235);
  and2 I586_236(w_586_230, w_579_461, w_586_236);
  not1 I587_009(w_587_009, w_359_198);
  nand2 I587_090(w_587_090, w_490_089, w_528_017);
  nand2 I587_141(w_587_141, w_113_015, w_420_607);
  nand2 I587_230(w_587_230, w_043_033, w_337_412);
  not1 I587_313(w_587_313, w_106_096);
  not1 I588_111(w_588_111, w_020_042);
  and2 I588_153(w_588_153, w_177_085, w_554_069);
  and2 I588_164(w_588_164, w_043_038, w_469_024);
  not1 I589_007(w_589_007, w_200_448);
  not1 I589_022(w_589_022, w_479_185);
  not1 I589_092(w_589_092, w_342_047);
  or2  I589_154(w_589_154, w_267_276, w_505_074);
  not1 I589_331(w_589_331, w_519_041);
  not1 I590_003(w_590_003, w_284_145);
  nand2 I590_026(w_590_026, w_375_032, w_389_234);
  not1 I590_161(w_590_161, w_035_074);
  and2 I591_057(w_591_057, w_052_022, w_398_067);
  nand2 I591_101(w_591_101, w_423_092, w_579_358);
  and2 I591_190(w_591_190, w_300_139, w_328_120);
  and2 I591_221(w_591_223, w_591_222, w_452_300);
  or2  I591_222(w_591_224, w_591_239, w_591_223);
  not1 I591_223(w_591_225, w_591_224);
  or2  I591_224(w_591_226, w_591_225, w_537_264);
  and2 I591_225(w_591_227, w_317_162, w_591_226);
  or2  I591_226(w_591_222, w_320_019, w_591_227);
  or2  I591_227(w_591_232, w_423_057, w_591_231);
  and2 I591_228(w_591_233, w_463_192, w_591_232);
  not1 I591_229(w_591_234, w_591_233);
  nand2 I591_230(w_591_235, w_268_038, w_591_234);
  not1 I591_231(w_591_236, w_591_235);
  and2 I591_232(w_591_237, w_299_015, w_591_236);
  not1 I591_233(w_591_231, w_591_224);
  and2 I591_234(w_591_239, w_231_220, w_591_237);
  or2  I592_177(w_592_177, w_300_085, w_533_329);
  or2  I592_233(w_592_233, w_360_373, w_274_100);
  nand2 I592_491(w_592_491, w_110_335, w_138_309);
  and2 I593_079(w_593_079, w_014_032, w_273_054);
  not1 I593_161(w_593_161, w_245_507);
  and2 I594_104(w_594_104, w_412_202, w_457_164);
  nand2 I594_121(w_594_121, w_234_145, w_120_104);
  not1 I595_029(w_595_029, w_286_275);
  not1 I595_130(w_595_130, w_508_396);
  and2 I595_157(w_595_157, w_464_242, w_506_513);
  or2  I595_246(w_595_246, w_137_164, w_175_103);
  nand2 I596_010(w_596_010, w_180_015, w_354_112);
  nand2 I596_068(w_596_068, w_323_089, w_286_037);
  nand2 I596_137(w_596_137, w_225_051, w_239_000);
  not1 I596_405(w_596_405, w_123_056);
  not1 I597_258(w_597_258, w_359_089);
  not1 I598_010(w_598_010, w_575_000);
  and2 I598_017(w_598_017, w_434_382, w_490_019);
  or2  I598_028(w_598_028, w_383_618, w_336_209);
  not1 I599_018(w_599_018, w_048_010);
  nand2 I599_025(w_599_025, w_125_059, w_573_058);
  or2  I599_032(w_599_032, w_493_103, w_376_055);
  or2  I600_084(w_600_084, w_240_125, w_362_031);
  or2  I600_130(w_600_130, w_026_709, w_314_174);
  not1 I600_264(w_600_264, w_131_511);
  and2 I600_697(w_600_697, w_224_331, w_563_022);
  or2  I601_071(w_601_071, w_353_137, w_425_247);
  not1 I601_073(w_601_073, w_259_551);
  nand2 I601_077(w_601_077, w_493_038, w_416_168);
  nand2 I601_123(w_601_123, w_286_130, w_502_539);
  not1 I601_384(w_601_384, w_006_093);
  nand2 I601_583(w_601_583, w_349_214, w_420_673);
  nand2 I602_005(w_602_005, w_089_160, w_436_224);
  not1 I602_296(w_602_296, w_157_101);
  or2  I603_090(w_603_090, w_406_280, w_207_086);
  nand2 I603_123(w_603_123, w_600_130, w_563_470);
  and2 I603_163(w_603_163, w_060_194, w_362_337);
  and2 I603_183(w_603_185, w_603_184, w_549_107);
  and2 I603_184(w_603_186, w_603_185, w_603_197);
  not1 I603_185(w_603_184, w_603_186);
  not1 I603_186(w_603_191, w_603_190);
  not1 I603_187(w_603_192, w_603_191);
  or2  I603_188(w_603_193, w_406_282, w_603_192);
  nand2 I603_189(w_603_194, w_603_193, w_582_461);
  and2 I603_190(w_603_195, w_603_194, w_226_401);
  not1 I603_191(w_603_190, w_603_186);
  and2 I603_192(w_603_197, w_009_583, w_603_195);
  not1 I604_108(w_604_108, w_098_003);
  and2 I604_237(w_604_237, w_593_161, w_524_346);
  nand2 I605_212(w_605_212, w_320_297, w_490_012);
  not1 I605_658(w_605_658, w_503_252);
  or2  I607_016(w_607_016, w_171_363, w_166_040);
  not1 I608_014(w_608_014, w_511_240);
  not1 I608_218(w_608_218, w_218_576);
  or2  I608_359(w_608_359, w_207_198, w_445_012);
  not1 I608_384(w_608_384, w_209_018);
  or2  I609_050(w_609_050, w_403_216, w_561_308);
  and2 I609_187(w_609_187, w_217_020, w_045_239);
  and2 I609_233(w_609_233, w_568_499, w_039_072);
  nand2 I610_041(w_610_041, w_557_062, w_222_521);
  or2  I610_051(w_610_051, w_372_033, w_584_712);
  or2  I610_104(w_610_104, w_123_172, w_308_115);
  nand2 I611_282(w_611_282, w_574_373, w_530_147);
  nand2 I611_485(w_611_485, w_425_000, w_561_079);
  nand2 I612_076(w_612_076, w_177_258, w_213_466);
  and2 I612_103(w_612_103, w_531_012, w_567_014);
  or2  I613_009(w_613_009, w_014_195, w_570_085);
  nand2 I613_024(w_613_024, w_385_089, w_028_234);
  or2  I613_030(w_613_030, w_012_009, w_308_067);
  not1 I613_089(w_613_089, w_513_076);
  or2  I614_253(w_614_253, w_124_035, w_499_376);
  nand2 I614_334(w_614_334, w_466_066, w_401_244);
  nand2 I615_023(w_615_023, w_138_125, w_275_049);
  nand2 I615_033(w_615_033, w_006_122, w_488_021);
  and2 I615_034(w_615_034, w_372_031, w_173_018);
  and2 I615_052(w_615_052, w_134_018, w_437_429);
  nand2 I615_067(w_615_067, w_333_314, w_386_080);
  not1 I615_078(w_615_078, w_490_067);
  or2  I615_079(w_615_079, w_379_099, w_537_154);
  or2  I616_232(w_616_232, w_586_090, w_373_092);
  not1 I616_388(w_616_388, w_561_038);
  or2  I617_086(w_617_086, w_199_040, w_523_087);
  nand2 I617_233(w_617_233, w_269_171, w_412_076);
  nand2 I618_009(w_618_009, w_232_332, w_153_030);
  not1 I618_048(w_618_048, w_475_296);
  or2  I618_060(w_618_060, w_051_246, w_579_647);
  not1 I619_167(w_619_167, w_167_050);
  nand2 I619_251(w_619_251, w_256_089, w_452_125);
  nand2 I619_510(w_619_510, w_314_032, w_185_140);
  and2 I620_002(w_620_002, w_618_009, w_174_010);
  nand2 I620_106(w_620_106, w_617_233, w_003_021);
  not1 I620_438(w_620_438, w_493_044);
  nand2 I620_440(w_620_440, w_429_137, w_206_002);
  or2  I621_230(w_621_230, w_500_203, w_204_011);
  or2  I621_444(w_621_444, w_132_094, w_117_012);
  or2  I622_033(w_622_033, w_282_236, w_039_513);
  or2  I622_037(w_622_037, w_337_356, w_255_024);
  not1 I622_064(w_622_064, w_023_201);
  nand2 I622_074(w_622_074, w_296_041, w_347_016);
  and2 I623_081(w_623_081, w_428_181, w_440_040);
  not1 I623_364(w_623_364, w_002_328);
  not1 I624_018(w_624_018, w_235_079);
  nand2 I624_070(w_624_070, w_096_005, w_445_069);
  not1 I625_100(w_625_100, w_001_016);
  not1 I625_277(w_625_277, w_373_013);
  nand2 I626_011(w_626_011, w_187_015, w_451_006);
  and2 I626_319(w_626_319, w_126_144, w_287_334);
  nand2 I626_338(w_626_338, w_368_022, w_134_374);
  and2 I626_796(w_626_798, w_626_797, w_380_615);
  or2  I626_797(w_626_799, w_626_798, w_626_820);
  and2 I626_798(w_626_800, w_576_172, w_626_799);
  nand2 I626_799(w_626_801, w_480_029, w_626_800);
  or2  I626_800(w_626_802, w_081_005, w_626_801);
  not1 I626_801(w_626_803, w_626_802);
  and2 I626_802(w_626_804, w_626_803, w_127_027);
  not1 I626_803(w_626_797, w_626_804);
  nand2 I626_804(w_626_809, w_499_548, w_626_808);
  and2 I626_805(w_626_810, w_110_401, w_626_809);
  not1 I626_806(w_626_811, w_626_810);
  nand2 I626_807(w_626_812, w_163_489, w_626_811);
  nand2 I626_808(w_626_813, w_626_812, w_011_624);
  not1 I626_809(w_626_814, w_626_813);
  nand2 I626_810(w_626_815, w_626_814, w_596_010);
  and2 I626_811(w_626_816, w_626_815, w_406_004);
  and2 I626_812(w_626_817, w_626_816, w_058_504);
  and2 I626_813(w_626_818, w_626_817, w_401_246);
  not1 I626_814(w_626_808, w_626_799);
  and2 I626_815(w_626_820, w_512_434, w_626_818);
  or2  I626_816(w_626_823, w_626_822, w_484_249);
  or2  I626_817(w_626_824, w_626_823, w_355_071);
  or2  I626_818(w_626_825, w_626_824, w_412_398);
  nand2 I626_819(w_626_826, w_626_825, w_181_169);
  nand2 I626_820(w_626_827, w_626_826, w_336_002);
  not1 I626_821(w_626_828, w_626_827);
  not1 I626_822(w_626_829, w_626_828);
  and2 I626_823(w_626_830, w_626_829, w_290_005);
  and2 I626_824(w_626_831, w_071_188, w_626_830);
  not1 I626_825(w_626_832, w_626_831);
  and2 I626_826(w_626_833, w_344_061, w_626_832);
  not1 I626_827(w_626_822, w_626_833);
  or2  I628_056(w_628_056, w_180_011, w_286_136);
  nand2 I628_074(w_628_074, w_573_043, w_399_118);
  not1 I628_151(w_628_151, w_468_079);
  nand2 I629_146(w_629_146, w_288_420, w_194_170);
  not1 I629_161(w_629_161, w_527_223);
  not1 I629_191(w_629_191, w_308_147);
  or2  I629_624(w_629_624, w_148_164, w_589_007);
  and2 I630_049(w_630_049, w_444_585, w_559_020);
  and2 I630_052(w_630_052, w_426_017, w_006_248);
  and2 I631_130(w_631_130, w_023_114, w_316_450);
  and2 I631_326(w_631_326, w_589_092, w_224_178);
  or2  I633_039(w_633_039, w_545_349, w_153_029);
  nand2 I633_744(w_633_744, w_065_537, w_043_005);
  not1 I634_179(w_634_179, w_010_759);
  nand2 I634_264(w_634_264, w_493_050, w_107_355);
  nand2 I634_295(w_634_295, w_628_056, w_319_289);
  and2 I635_039(w_635_039, w_252_306, w_270_335);
  or2  I635_156(w_635_156, w_620_106, w_096_002);
  not1 I635_170(w_635_170, w_079_003);
  not1 I635_484(w_635_484, w_165_110);
  nand2 I636_078(w_636_078, w_103_026, w_483_358);
  nand2 I636_112(w_636_112, w_107_103, w_601_073);
  nand2 I636_159(w_636_159, w_033_618, w_183_270);
  or2  I637_003(w_637_003, w_445_025, w_075_138);
  and2 I637_010(w_637_010, w_091_036, w_624_018);
  or2  I637_242(w_637_242, w_482_175, w_192_099);
  nand2 I638_261(w_638_261, w_434_098, w_414_089);
  or2  I638_350(w_638_350, w_225_180, w_122_081);
  nand2 I638_380(w_638_380, w_620_440, w_354_010);
  or2  I638_423(w_638_423, w_265_418, w_448_260);
  or2  I638_470(w_638_470, w_487_101, w_216_301);
  or2  I639_000(w_639_000, w_384_149, w_466_296);
  nand2 I639_018(w_639_018, w_454_305, w_467_177);
  and2 I640_029(w_640_029, w_561_175, w_451_105);
  and2 I640_267(w_640_267, w_367_035, w_572_107);
  nand2 I640_443(w_640_443, w_318_004, w_187_013);
  nand2 I640_456(w_640_456, w_140_074, w_638_423);
  and2 I640_532(w_640_532, w_372_038, w_076_161);
  nand2 I640_598(w_640_598, w_267_014, w_034_057);
  nand2 I640_653(w_640_653, w_439_116, w_431_210);
  and2 I641_058(w_641_058, w_523_003, w_293_101);
  and2 I641_063(w_641_063, w_475_511, w_401_008);
  and2 I641_072(w_641_072, w_492_319, w_623_081);
  and2 I642_569(w_642_569, w_427_059, w_344_455);
  or2  I643_008(w_643_008, w_591_190, w_011_117);
  and2 I643_030(w_643_030, w_339_039, w_423_019);
  and2 I643_303(w_643_303, w_317_014, w_059_057);
  not1 I644_011(w_644_011, w_420_483);
  or2  I645_314(w_645_314, w_447_160, w_084_014);
  and2 I646_003(w_646_003, w_354_039, w_116_224);
  or2  I646_007(w_646_007, w_074_209, w_639_018);
  or2  I646_009(w_646_009, w_048_003, w_325_139);
  and2 I646_013(w_646_013, w_021_068, w_004_221);
  or2  I647_193(w_647_193, w_517_098, w_231_322);
  and2 I647_200(w_647_200, w_228_343, w_610_051);
  not1 I647_366(w_647_366, w_454_039);
  not1 I647_367(w_647_367, w_173_009);
  and2 I647_393(w_647_393, w_138_093, w_267_217);
  or2  I647_446(w_647_446, w_310_557, w_643_008);
  or2  I647_488(w_647_488, w_052_008, w_615_034);
  or2  I648_040(w_648_040, w_143_209, w_364_013);
  nand2 I648_041(w_648_041, w_236_199, w_466_053);
  or2  I648_079(w_648_079, w_465_165, w_135_457);
  and2 I649_021(w_649_021, w_211_003, w_227_612);
  or2  I649_026(w_649_026, w_048_013, w_561_205);
  not1 I649_029(w_649_031, w_649_030);
  not1 I649_030(w_649_032, w_649_031);
  or2  I649_031(w_649_033, w_649_032, w_621_444);
  not1 I649_032(w_649_034, w_649_033);
  and2 I649_033(w_649_035, w_649_034, w_441_505);
  or2  I649_034(w_649_030, w_649_035, w_649_049);
  not1 I649_035(w_649_040, w_649_039);
  or2  I649_036(w_649_041, w_433_213, w_649_040);
  or2  I649_037(w_649_042, w_649_041, w_300_261);
  nand2 I649_038(w_649_043, w_649_042, w_442_123);
  and2 I649_039(w_649_044, w_649_043, w_563_052);
  not1 I649_040(w_649_045, w_649_044);
  nand2 I649_041(w_649_046, w_649_045, w_647_366);
  and2 I649_042(w_649_047, w_257_101, w_649_046);
  not1 I649_043(w_649_039, w_649_030);
  and2 I649_044(w_649_049, w_527_526, w_649_047);
  not1 I650_341(w_650_341, w_619_167);
  not1 I650_578(w_650_578, w_527_197);
  nand2 I650_741(w_650_741, w_270_037, w_201_141);
  not1 I651_019(w_651_019, w_628_151);
  or2  I651_337(w_651_337, w_506_594, w_350_022);
  not1 I651_464(w_651_464, w_590_003);
  not1 I652_014(w_652_014, w_552_304);
  and2 I652_020(w_652_020, w_076_036, w_269_019);
  or2  I652_030(w_652_030, w_193_190, w_175_208);
  or2  I652_041(w_652_041, w_131_432, w_535_202);
  nand2 I652_042(w_652_042, w_530_096, w_148_611);
  and2 I652_061(w_652_061, w_142_129, w_219_644);
  nand2 I653_035(w_653_035, w_652_030, w_244_071);
  nand2 I653_063(w_653_063, w_350_094, w_168_359);
  nand2 I653_094(w_653_094, w_184_112, w_575_160);
  or2  I653_188(w_653_188, w_394_080, w_539_538);
  not1 I653_262(w_653_262, w_000_102);
  and2 I654_153(w_654_153, w_027_187, w_261_005);
  not1 I654_308(w_654_308, w_407_356);
  nand2 I654_336(w_654_336, w_468_035, w_243_072);
  and2 I654_410(w_654_412, w_138_192, w_654_411);
  and2 I654_411(w_654_413, w_654_412, w_280_098);
  not1 I654_412(w_654_414, w_654_413);
  nand2 I654_413(w_654_415, w_654_414, w_148_698);
  not1 I654_414(w_654_416, w_654_415);
  and2 I654_415(w_654_417, w_654_416, w_615_052);
  not1 I654_416(w_654_411, w_654_417);
  and2 I655_478(w_655_478, w_092_690, w_286_190);
  and2 I656_067(w_656_067, w_418_029, w_477_070);
  nand2 I656_087(w_656_087, w_504_031, w_312_023);
  and2 I656_298(w_656_298, w_120_060, w_244_081);
  and2 I656_348(w_656_348, w_467_284, w_091_041);
  or2  I656_595(w_656_597, w_356_043, w_656_596);
  or2  I656_596(w_656_598, w_261_100, w_656_597);
  nand2 I656_597(w_656_599, w_621_230, w_656_598);
  or2  I656_598(w_656_600, w_402_032, w_656_599);
  nand2 I656_599(w_656_601, w_624_070, w_656_600);
  nand2 I656_600(w_656_602, w_656_601, w_221_071);
  nand2 I656_601(w_656_603, w_656_602, w_079_054);
  and2 I656_602(w_656_604, w_045_367, w_656_603);
  or2  I656_603(w_656_605, w_656_604, w_546_450);
  not1 I656_604(w_656_606, w_656_605);
  and2 I656_605(w_656_607, w_462_400, w_656_606);
  not1 I656_606(w_656_596, w_656_607);
  not1 I658_054(w_658_054, w_093_067);
  not1 I658_094(w_658_094, w_587_141);
  or2  I658_262(w_658_262, w_435_156, w_353_047);
  or2  I659_239(w_659_239, w_533_532, w_204_473);
  nand2 I660_000(w_660_000, w_020_118, w_305_239);
  not1 I660_001(w_660_001, w_588_164);
  and2 I661_018(w_661_018, w_277_293, w_247_079);
  or2  I661_049(w_661_049, w_169_106, w_597_258);
  not1 I662_321(w_662_321, w_575_178);
  not1 I663_023(w_663_023, w_302_495);
  and2 I663_060(w_663_060, w_092_159, w_472_163);
  and2 I663_070(w_663_070, w_635_039, w_519_022);
  and2 I663_094(w_663_094, w_417_083, w_109_213);
  or2  I664_018(w_664_018, w_393_113, w_136_024);
  nand2 I664_103(w_664_103, w_560_071, w_398_043);
  or2  I664_123(w_664_123, w_294_000, w_159_007);
  nand2 I664_155(w_664_155, w_035_013, w_378_022);
  and2 I665_027(w_665_027, w_596_068, w_234_159);
  and2 I665_424(w_665_424, w_039_039, w_423_038);
  not1 I666_406(w_666_406, w_581_400);
  not1 I666_445(w_666_445, w_617_086);
  nand2 I667_051(w_667_051, w_336_177, w_289_257);
  and2 I667_625(w_667_625, w_036_097, w_018_008);
  and2 I668_171(w_668_171, w_192_008, w_450_067);
  nand2 I669_108(w_669_108, w_503_190, w_334_139);
  not1 I669_152(w_669_152, w_432_136);
  and2 I669_254(w_669_254, w_149_075, w_272_040);
  not1 I669_261(w_669_261, w_639_000);
  nand2 I669_298(w_669_298, w_036_175, w_598_010);
  nand2 I669_307(w_669_307, w_419_240, w_095_053);
  not1 I670_022(w_670_022, w_280_687);
  nand2 I670_024(w_670_024, w_135_089, w_486_111);
  not1 I670_045(w_670_045, w_339_022);
  nand2 I671_371(w_671_371, w_500_226, w_131_120);
  nand2 I673_161(w_673_161, w_174_096, w_591_057);
  not1 I673_278(w_673_278, w_482_327);
  or2  I673_419(w_673_419, w_330_042, w_557_047);
  nand2 I674_172(w_674_172, w_116_122, w_231_009);
  and2 I674_360(w_674_360, w_411_581, w_277_364);
  and2 I675_109(w_675_109, w_054_155, w_072_156);
  not1 I675_146(w_675_146, w_628_074);
  and2 I675_252(w_675_252, w_485_072, w_033_291);
  nand2 I675_318(w_675_318, w_252_368, w_279_171);
  not1 I676_185(w_676_185, w_410_048);
  not1 I676_222(w_676_222, w_010_235);
  nand2 I676_258(w_676_258, w_667_625, w_298_073);
  not1 I677_020(w_677_020, w_185_103);
  and2 I677_131(w_677_131, w_303_121, w_325_035);
  nand2 I678_049(w_678_049, w_525_007, w_008_033);
  not1 I678_201(w_678_201, w_670_045);
  nand2 I678_225(w_678_225, w_049_231, w_252_229);
  and2 I678_454(w_678_454, w_359_154, w_516_079);
  not1 I679_286(w_679_286, w_034_021);
  and2 I679_443(w_679_443, w_126_193, w_164_004);
  nand2 I679_618(w_679_618, w_052_023, w_261_032);
  and2 I680_105(w_680_105, w_546_073, w_013_166);
  and2 I680_186(w_680_186, w_491_022, w_337_225);
  or2  I681_081(w_681_081, w_397_019, w_404_022);
  not1 I681_252(w_681_252, w_282_327);
  not1 I681_320(w_681_320, w_494_046);
  not1 I682_371(w_682_371, w_430_534);
  or2  I682_399(w_682_399, w_286_377, w_298_099);
  or2  I682_472(w_682_472, w_368_081, w_654_308);
  or2  I682_543(w_682_543, w_024_197, w_482_003);
  not1 I682_715(w_682_717, w_682_716);
  and2 I682_716(w_682_718, w_682_717, w_682_732);
  nand2 I682_717(w_682_716, w_399_098, w_682_718);
  or2  I682_718(w_682_723, w_682_722, w_039_561);
  not1 I682_719(w_682_724, w_682_723);
  nand2 I682_720(w_682_725, w_682_724, w_160_465);
  nand2 I682_721(w_682_726, w_682_725, w_652_061);
  and2 I682_722(w_682_727, w_682_726, w_507_035);
  or2  I682_723(w_682_728, w_682_727, w_398_058);
  nand2 I682_724(w_682_729, w_682_728, w_158_004);
  and2 I682_725(w_682_730, w_682_729, w_637_010);
  not1 I682_726(w_682_722, w_682_718);
  and2 I682_727(w_682_732, w_181_205, w_682_730);
  or2  I683_089(w_683_089, w_499_583, w_003_068);
  not1 I683_112(w_683_112, w_372_008);
  or2  I683_230(w_683_230, w_476_274, w_643_030);
  and2 I683_259(w_683_259, w_202_286, w_140_027);
  and2 I685_294(w_685_294, w_239_000, w_427_051);
  or2  I685_299(w_685_299, w_116_118, w_192_153);
  and2 I686_011(w_686_011, w_211_021, w_238_000);
  or2  I686_026(w_686_026, w_270_017, w_247_183);
  not1 I686_102(w_686_102, w_116_004);
  nand2 I686_107(w_686_107, w_281_133, w_175_156);
  and2 I687_198(w_687_198, w_242_000, w_601_583);
  not1 I688_036(w_688_036, w_120_516);
  or2  I688_387(w_688_387, w_303_080, w_604_108);
  or2  I688_501(w_688_501, w_251_130, w_664_103);
  or2  I688_748(w_688_750, w_688_770, w_688_749);
  not1 I688_749(w_688_751, w_688_750);
  not1 I688_750(w_688_752, w_688_751);
  or2  I688_751(w_688_753, w_688_752, w_163_307);
  nand2 I688_752(w_688_754, w_688_753, w_573_324);
  and2 I688_753(w_688_755, w_688_754, w_110_279);
  nand2 I688_754(w_688_756, w_688_755, w_488_102);
  and2 I688_755(w_688_757, w_474_160, w_688_756);
  or2  I688_756(w_688_749, w_688_757, w_584_341);
  and2 I688_757(w_688_762, w_301_091, w_688_761);
  and2 I688_758(w_688_763, w_688_762, w_134_122);
  and2 I688_759(w_688_764, w_688_763, w_165_079);
  nand2 I688_760(w_688_765, w_393_194, w_688_764);
  or2  I688_761(w_688_766, w_257_318, w_688_765);
  or2  I688_762(w_688_767, w_092_489, w_688_766);
  and2 I688_763(w_688_768, w_675_146, w_688_767);
  not1 I688_764(w_688_761, w_688_750);
  and2 I688_765(w_688_770, w_303_059, w_688_768);
  and2 I689_090(w_689_090, w_567_003, w_159_078);
  and2 I689_226(w_689_226, w_065_327, w_673_278);
  and2 I689_227(w_689_227, w_098_063, w_110_026);
  and2 I689_232(w_689_234, w_689_233, w_113_029);
  nand2 I689_233(w_689_235, w_689_234, w_646_009);
  not1 I689_234(w_689_236, w_689_235);
  nand2 I689_235(w_689_237, w_484_329, w_689_236);
  nand2 I689_236(w_689_238, w_689_237, w_098_061);
  and2 I689_237(w_689_239, w_203_015, w_689_238);
  nand2 I689_238(w_689_240, w_689_239, w_661_018);
  and2 I689_239(w_689_241, w_689_240, w_161_565);
  and2 I689_240(w_689_233, w_689_241, w_005_100);
  and2 I690_025(w_690_025, w_601_077, w_286_380);
  not1 I690_051(w_690_053, w_690_052);
  and2 I690_052(w_690_054, w_411_567, w_690_053);
  and2 I690_053(w_690_055, w_484_349, w_690_054);
  and2 I690_054(w_690_056, w_690_055, w_609_233);
  or2  I690_055(w_690_052, w_419_155, w_690_056);
  or2  I691_005(w_691_005, w_611_282, w_051_017);
  or2  I691_139(w_691_139, w_590_026, w_331_247);
  nand2 I692_155(w_692_155, w_383_018, w_619_510);
  not1 I692_168(w_692_168, w_303_095);
  and2 I693_031(w_693_031, w_630_052, w_626_319);
  not1 I693_163(w_693_163, w_569_133);
  nand2 I693_193(w_693_193, w_647_193, w_223_201);
  not1 I693_292(w_693_292, w_021_091);
  nand2 I693_319(w_693_319, w_106_170, w_047_024);
  nand2 I693_324(w_693_324, w_652_014, w_650_578);
  or2  I694_002(w_694_002, w_575_094, w_077_378);
  or2  I694_018(w_694_018, w_529_000, w_688_387);
  not1 I694_021(w_694_021, w_490_093);
  nand2 I694_029(w_694_029, w_076_145, w_547_002);
  not1 I695_052(w_695_052, w_151_068);
  nand2 I695_312(w_695_314, w_695_325, w_695_313);
  nand2 I695_313(w_695_315, w_695_314, w_575_064);
  and2 I695_314(w_695_316, w_309_193, w_695_315);
  and2 I695_315(w_695_313, w_206_087, w_695_316);
  or2  I695_316(w_695_321, w_695_320, w_688_036);
  and2 I695_317(w_695_322, w_327_440, w_695_321);
  and2 I695_318(w_695_323, w_695_322, w_673_419);
  not1 I695_319(w_695_320, w_695_314);
  and2 I695_320(w_695_325, w_015_647, w_695_323);
  and2 I696_115(w_696_115, w_057_215, w_200_127);
  not1 I697_033(w_697_033, w_319_200);
  or2  I697_187(w_697_187, w_404_182, w_674_172);
  or2  I697_213(w_697_213, w_010_351, w_401_158);
  not1 I699_036(w_699_036, w_088_119);
  not1 I699_231(w_699_231, w_444_425);
  or2  I699_724(w_699_724, w_370_051, w_028_183);
  and2 I701_033(w_701_033, w_603_090, w_432_300);
  or2  I701_054(w_701_054, w_694_002, w_013_157);
  not1 I701_157(w_701_157, w_023_040);
  not1 I702_148(w_702_148, w_217_006);
  nand2 I703_135(w_703_135, w_135_111, w_291_110);
  or2  I703_220(w_703_220, w_309_380, w_194_132);
  not1 I703_306(w_703_306, w_644_011);
  or2  I704_043(w_704_043, w_106_127, w_699_036);
  not1 I704_140(w_704_140, w_322_015);
  and2 I704_721(w_704_723, w_704_722, w_333_158);
  or2  I704_722(w_704_724, w_704_723, w_326_077);
  not1 I704_723(w_704_725, w_704_724);
  not1 I704_724(w_704_726, w_704_725);
  not1 I704_725(w_704_727, w_704_726);
  or2  I704_726(w_704_728, w_365_045, w_704_727);
  and2 I704_727(w_704_729, w_704_728, w_506_611);
  or2  I704_728(w_704_730, w_157_064, w_704_729);
  or2  I704_729(w_704_731, w_238_395, w_704_730);
  and2 I704_730(w_704_732, w_704_731, w_535_252);
  not1 I704_731(w_704_722, w_704_732);
  nand2 I705_453(w_705_455, w_705_454, w_224_524);
  and2 I705_454(w_705_456, w_622_064, w_705_455);
  or2  I705_455(w_705_457, w_648_040, w_705_456);
  and2 I705_456(w_705_458, w_705_457, w_447_336);
  nand2 I705_457(w_705_459, w_705_458, w_694_021);
  nand2 I705_458(w_705_460, w_705_459, w_649_021);
  nand2 I705_459(w_705_461, w_047_320, w_705_460);
  not1 I705_460(w_705_462, w_705_461);
  and2 I705_461(w_705_463, w_292_033, w_705_462);
  not1 I705_462(w_705_454, w_705_463);
  nand2 I706_205(w_706_205, w_227_485, w_424_228);
  nand2 I706_227(w_706_227, w_095_031, w_515_172);
  not1 I707_117(w_707_117, w_545_151);
  nand2 I707_118(w_707_118, w_566_198, w_484_326);
  and2 I708_064(w_708_064, w_226_219, w_636_078);
  not1 I708_269(w_708_269, w_429_259);
  not1 I709_559(w_709_559, w_126_120);
  not1 I710_119(w_710_119, w_390_148);
  and2 I711_004(w_711_004, w_457_154, w_117_046);
  and2 I711_018(w_711_018, w_415_283, w_638_261);
  and2 I711_030(w_711_030, w_594_104, w_242_090);
  nand2 I711_048(w_711_048, w_665_424, w_121_134);
  nand2 I711_050(w_711_052, w_711_051, w_014_234);
  or2  I711_051(w_711_053, w_711_052, w_308_123);
  and2 I711_052(w_711_054, w_711_067, w_711_053);
  and2 I711_053(w_711_051, w_360_150, w_711_054);
  or2  I711_054(w_711_059, w_179_416, w_711_058);
  not1 I711_055(w_711_060, w_711_059);
  nand2 I711_056(w_711_061, w_659_239, w_711_060);
  and2 I711_057(w_711_062, w_079_059, w_711_061);
  nand2 I711_058(w_711_063, w_488_037, w_711_062);
  and2 I711_059(w_711_064, w_593_079, w_711_063);
  and2 I711_060(w_711_065, w_711_064, w_245_035);
  not1 I711_061(w_711_058, w_711_054);
  and2 I711_062(w_711_067, w_556_270, w_711_065);
  not1 I712_033(w_712_033, w_205_462);
  or2  I712_065(w_712_065, w_386_015, w_200_214);
  and2 I714_000(w_714_000, w_345_250, w_460_173);
  not1 I714_009(w_714_009, w_615_079);
  and2 I714_021(w_714_021, w_211_037, w_442_126);
  nand2 I714_046(w_714_046, w_124_094, w_163_243);
  and2 I716_018(w_716_018, w_039_256, w_130_035);
  nand2 I716_029(w_716_029, w_678_049, w_694_029);
  or2  I717_116(w_717_116, w_287_020, w_164_387);
  nand2 I718_123(w_718_123, w_413_083, w_636_159);
  or2  I718_200(w_718_200, w_537_032, w_524_591);
  or2  I718_258(w_718_258, w_552_100, w_191_033);
  nand2 I718_277(w_718_277, w_693_193, w_544_146);
  not1 I718_646(w_718_646, w_017_288);
  not1 I719_004(w_719_004, w_203_297);
  nand2 I719_150(w_719_150, w_613_030, w_136_014);
  or2  I719_250(w_719_250, w_542_007, w_574_265);
  nand2 I719_393(w_719_393, w_408_005, w_508_005);
  or2  I721_517(w_721_517, w_584_255, w_324_008);
  not1 I722_415(w_722_415, w_653_035);
  or2  I723_559(w_723_559, w_339_039, w_154_039);
  not1 I723_597(w_723_597, w_438_273);
  and2 I724_311(w_724_311, w_498_170, w_468_090);
  or2  I724_391(w_724_391, w_312_133, w_304_079);
  and2 I724_451(w_724_451, w_704_140, w_675_318);
  nand2 I725_058(w_725_058, w_484_346, w_701_157);
  and2 I725_102(w_725_102, w_125_397, w_683_230);
  not1 I725_342(w_725_342, w_322_005);
  not1 I726_165(w_726_165, w_238_195);
  or2  I726_379(w_726_379, w_054_258, w_457_054);
  or2  I726_437(w_726_437, w_538_190, w_028_362);
  nand2 I727_106(w_727_106, w_100_021, w_547_002);
  or2  I728_136(w_728_136, w_232_318, w_683_089);
  or2  I728_394(w_728_394, w_427_053, w_205_076);
  nand2 I728_548(w_728_548, w_680_186, w_530_219);
  nand2 I728_788(w_728_790, w_098_069, w_728_789);
  nand2 I728_789(w_728_791, w_728_790, w_093_050);
  not1 I728_790(w_728_792, w_728_791);
  or2  I728_791(w_728_793, w_728_792, w_551_012);
  or2  I728_792(w_728_794, w_728_793, w_653_094);
  not1 I728_793(w_728_795, w_728_794);
  nand2 I728_794(w_728_796, w_728_795, w_210_030);
  and2 I728_795(w_728_797, w_728_796, w_388_076);
  nand2 I728_796(w_728_789, w_573_223, w_728_797);
  or2  I729_360(w_729_360, w_427_050, w_356_001);
  or2  I730_122(w_730_122, w_663_070, w_066_290);
  or2  I730_150(w_730_150, w_154_002, w_468_070);
  not1 I730_158(w_730_160, w_730_159);
  nand2 I730_159(w_730_161, w_094_545, w_730_160);
  or2  I730_160(w_730_162, w_730_161, w_303_128);
  and2 I730_161(w_730_163, w_539_388, w_730_162);
  or2  I730_162(w_730_164, w_191_306, w_730_163);
  and2 I730_163(w_730_165, w_730_164, w_043_011);
  or2  I730_164(w_730_166, w_158_004, w_730_165);
  and2 I730_165(w_730_167, w_666_406, w_730_166);
  or2  I730_166(w_730_168, w_730_167, w_163_189);
  and2 I730_167(w_730_169, w_730_168, w_434_495);
  not1 I730_168(w_730_159, w_730_169);
  and2 I731_077(w_731_077, w_275_489, w_039_374);
  nand2 I731_087(w_731_087, w_022_279, w_614_253);
  and2 I731_103(w_731_103, w_313_231, w_209_255);
  nand2 I731_119(w_731_119, w_202_105, w_568_367);
  nand2 I731_122(w_731_122, w_414_241, w_647_488);
  nand2 I731_147(w_731_147, w_539_723, w_009_336);
  and2 I731_181(w_731_181, w_254_073, w_678_454);
  not1 I731_186(w_731_186, w_663_023);
  nand2 I731_200(w_731_201, w_731_200, w_553_031);
  or2  I731_201(w_731_202, w_731_201, w_500_353);
  and2 I731_202(w_731_203, w_731_202, w_731_216);
  not1 I731_203(w_731_200, w_731_203);
  not1 I731_204(w_731_208, w_731_207);
  nand2 I731_205(w_731_209, w_260_183, w_731_208);
  or2  I731_206(w_731_210, w_731_209, w_029_033);
  or2  I731_207(w_731_211, w_272_039, w_731_210);
  and2 I731_208(w_731_212, w_731_211, w_642_569);
  and2 I731_209(w_731_213, w_710_119, w_731_212);
  and2 I731_210(w_731_214, w_655_478, w_731_213);
  not1 I731_211(w_731_207, w_731_203);
  and2 I731_212(w_731_216, w_403_315, w_731_214);
  or2  I732_016(w_732_016, w_269_356, w_393_136);
  and2 I733_045(w_733_045, w_189_298, w_226_310);
  or2  I733_100(w_733_100, w_413_045, w_193_087);
  nand2 I733_108(w_733_108, w_600_264, w_488_045);
  or2  I734_086(w_734_086, w_586_096, w_491_021);
  and2 I734_104(w_734_104, w_223_141, w_032_090);
  and2 I735_051(w_735_051, w_123_149, w_608_014);
  and2 I736_059(w_736_059, w_656_298, w_587_090);
  not1 I736_091(w_736_091, w_354_082);
  nand2 I736_389(w_736_389, w_165_009, w_457_002);
  or2  I737_012(w_737_012, w_175_594, w_592_233);
  or2  I737_115(w_737_115, w_585_101, w_410_142);
  and2 I737_620(w_737_622, w_191_362, w_737_621);
  not1 I737_621(w_737_623, w_737_622);
  nand2 I737_622(w_737_624, w_737_623, w_189_513);
  not1 I737_623(w_737_625, w_737_624);
  and2 I737_624(w_737_626, w_737_636, w_737_625);
  and2 I737_625(w_737_621, w_737_626, w_149_636);
  not1 I737_626(w_737_631, w_737_630);
  or2  I737_627(w_737_632, w_737_631, w_370_031);
  and2 I737_628(w_737_633, w_537_056, w_737_632);
  and2 I737_629(w_737_634, w_726_437, w_737_633);
  not1 I737_630(w_737_630, w_737_626);
  and2 I737_631(w_737_636, w_721_517, w_737_634);
  not1 I739_093(w_739_093, w_230_027);
  and2 I739_105(w_739_105, w_001_017, w_307_343);
  or2  I740_115(w_740_115, w_440_057, w_130_211);
  or2  I740_318(w_740_318, w_669_254, w_533_089);
  not1 I741_144(w_741_144, w_075_020);
  not1 I742_030(w_742_030, w_310_071);
  or2  I743_021(w_743_021, w_527_350, w_134_200);
  or2  I743_031(w_743_031, w_707_118, w_333_011);
  and2 I743_117(w_743_119, w_743_118, w_227_475);
  nand2 I743_118(w_743_120, w_743_119, w_198_014);
  nand2 I743_119(w_743_121, w_743_120, w_555_067);
  not1 I743_120(w_743_122, w_743_121);
  not1 I743_121(w_743_123, w_743_122);
  nand2 I743_122(w_743_124, w_743_123, w_678_225);
  not1 I743_123(w_743_125, w_743_124);
  or2  I743_124(w_743_126, w_743_125, w_353_443);
  nand2 I743_125(w_743_127, w_743_126, w_575_096);
  and2 I743_126(w_743_128, w_743_127, w_539_491);
  and2 I743_127(w_743_129, w_743_138, w_743_128);
  and2 I743_128(w_743_118, w_743_129, w_725_058);
  nand2 I743_129(w_743_134, w_048_002, w_743_133);
  and2 I743_130(w_743_135, w_130_044, w_743_134);
  and2 I743_131(w_743_136, w_743_135, w_615_067);
  not1 I743_132(w_743_133, w_743_129);
  and2 I743_133(w_743_138, w_469_069, w_743_136);
  nand2 I744_058(w_744_058, w_433_409, w_420_519);
  nand2 I744_072(w_744_072, w_359_176, w_311_003);
  and2 I746_141(w_746_141, w_293_359, w_694_018);
  nand2 I746_633(w_746_635, w_746_634, w_075_046);
  and2 I746_634(w_746_636, w_086_034, w_746_635);
  or2  I746_635(w_746_637, w_650_741, w_746_636);
  not1 I746_636(w_746_638, w_746_637);
  or2  I746_637(w_746_639, w_284_040, w_746_638);
  nand2 I746_638(w_746_640, w_106_052, w_746_639);
  not1 I746_639(w_746_641, w_746_640);
  and2 I746_640(w_746_642, w_516_096, w_746_641);
  or2  I746_641(w_746_634, w_093_059, w_746_642);
  or2  I747_019(w_747_019, w_718_258, w_400_009);
  not1 I748_126(w_748_126, w_334_640);
  or2  I748_161(w_748_161, w_265_120, w_676_222);
  not1 I748_267(w_748_267, w_651_019);
  not1 I749_059(w_749_059, w_207_468);
  not1 I749_131(w_749_131, w_647_200);
  nand2 I749_176(w_749_176, w_616_232, w_342_311);
  nand2 I750_434(w_750_434, w_622_037, w_286_186);
  nand2 I750_448(w_750_448, w_410_085, w_527_096);
  or2  I751_282(w_751_282, w_291_001, w_377_065);
  not1 I751_314(w_751_314, w_740_115);
  and2 I751_322(w_751_322, w_424_087, w_113_025);
  or2  I752_418(w_752_418, w_398_050, w_198_024);
  not1 I753_377(w_753_377, w_402_135);
  not1 I753_543(w_753_543, w_029_070);
  or2  I754_136(w_754_136, w_286_393, w_265_645);
  not1 I754_167(w_754_167, w_131_140);
  nand2 I755_016(w_755_016, w_039_492, w_406_221);
  not1 I756_003(w_756_003, w_648_041);
  not1 I756_070(w_756_070, w_653_262);
  or2  I756_072(w_756_072, w_592_491, w_118_101);
  nand2 I756_471(w_756_473, w_620_438, w_756_472);
  and2 I756_472(w_756_474, w_756_473, w_615_023);
  nand2 I756_473(w_756_475, w_756_474, w_590_161);
  and2 I756_474(w_756_476, w_357_381, w_756_475);
  nand2 I756_475(w_756_472, w_533_187, w_756_476);
  not1 I757_133(w_757_133, w_133_028);
  not1 I758_227(w_758_227, w_361_354);
  nand2 I759_047(w_759_047, w_393_016, w_669_108);
  and2 I759_108(w_759_108, w_100_081, w_260_017);
  and2 I759_124(w_759_124, w_658_262, w_008_414);
  or2  I759_642(w_759_642, w_601_071, w_656_067);
  nand2 I759_649(w_759_649, w_264_599, w_194_078);
  or2  I761_018(w_761_018, w_569_040, w_363_123);
  nand2 I761_022(w_761_022, w_448_104, w_640_029);
  or2  I762_061(w_762_061, w_189_025, w_264_470);
  and2 I762_123(w_762_123, w_296_302, w_322_017);
  and2 I762_253(w_762_253, w_113_010, w_664_123);
  nand2 I764_054(w_764_054, w_631_326, w_139_016);
  not1 I764_241(w_764_241, w_599_025);
  not1 I764_379(w_764_381, w_764_380);
  nand2 I764_380(w_764_382, w_229_086, w_764_381);
  and2 I764_381(w_764_383, w_764_382, w_188_107);
  nand2 I764_382(w_764_384, w_454_079, w_764_383);
  not1 I764_383(w_764_385, w_764_384);
  nand2 I764_384(w_764_386, w_631_130, w_764_385);
  nand2 I764_385(w_764_387, w_764_386, w_308_064);
  and2 I764_386(w_764_388, w_247_181, w_764_387);
  or2  I764_387(w_764_380, w_039_111, w_764_388);
  not1 I765_198(w_765_198, w_404_606);
  nand2 I766_300(w_766_300, w_454_025, w_669_298);
  and2 I766_315(w_766_317, w_380_317, w_766_316);
  not1 I766_316(w_766_318, w_766_317);
  nand2 I766_317(w_766_319, w_766_318, w_460_040);
  nand2 I766_318(w_766_320, w_616_388, w_766_319);
  and2 I766_319(w_766_321, w_302_529, w_766_320);
  or2  I766_320(w_766_322, w_766_321, w_766_344);
  and2 I766_321(w_766_323, w_043_045, w_766_322);
  and2 I766_322(w_766_324, w_766_323, w_157_032);
  nand2 I766_323(w_766_325, w_646_007, w_766_324);
  not1 I766_324(w_766_326, w_766_325);
  and2 I766_325(w_766_327, w_398_023, w_766_326);
  or2  I766_326(w_766_316, w_766_327, w_567_033);
  not1 I766_327(w_766_332, w_766_331);
  nand2 I766_328(w_766_333, w_073_649, w_766_332);
  not1 I766_329(w_766_334, w_766_333);
  nand2 I766_330(w_766_335, w_766_334, w_685_299);
  nand2 I766_331(w_766_336, w_707_117, w_766_335);
  not1 I766_332(w_766_337, w_766_336);
  nand2 I766_333(w_766_338, w_766_337, w_086_181);
  nand2 I766_334(w_766_339, w_464_299, w_766_338);
  not1 I766_335(w_766_340, w_766_339);
  nand2 I766_336(w_766_341, w_353_106, w_766_340);
  and2 I766_337(w_766_342, w_766_341, w_683_112);
  not1 I766_338(w_766_331, w_766_322);
  and2 I766_339(w_766_344, w_315_523, w_766_342);
  nand2 I767_284(w_767_284, w_105_052, w_665_027);
  and2 I768_275(w_768_277, w_768_276, w_768_296);
  not1 I768_276(w_768_278, w_768_277);
  nand2 I768_277(w_768_279, w_768_278, w_465_019);
  and2 I768_278(w_768_280, w_768_279, w_396_025);
  not1 I768_279(w_768_281, w_768_280);
  or2  I768_280(w_768_282, w_251_089, w_768_281);
  or2  I768_281(w_768_283, w_283_137, w_768_282);
  nand2 I768_282(w_768_284, w_768_283, w_061_160);
  or2  I768_283(w_768_285, w_768_284, w_428_124);
  nand2 I768_284(w_768_286, w_208_231, w_768_285);
  and2 I768_285(w_768_287, w_768_286, w_633_744);
  nand2 I768_286(w_768_276, w_513_576, w_768_287);
  and2 I768_287(w_768_292, w_768_291, w_392_245);
  or2  I768_288(w_768_293, w_768_292, w_731_119);
  and2 I768_289(w_768_294, w_768_293, w_729_360);
  not1 I768_290(w_768_291, w_768_277);
  and2 I768_291(w_768_296, w_371_000, w_768_294);
  nand2 I770_055(w_770_055, w_759_124, w_499_189);
  nand2 I770_072(w_770_072, w_394_040, w_211_005);
  not1 I772_073(w_772_073, w_105_249);
  nand2 I772_264(w_772_266, w_772_265, w_697_213);
  nand2 I772_265(w_772_267, w_772_283, w_772_266);
  and2 I772_266(w_772_268, w_772_267, w_284_123);
  not1 I772_267(w_772_269, w_772_268);
  or2  I772_268(w_772_270, w_449_218, w_772_269);
  and2 I772_269(w_772_271, w_582_245, w_772_270);
  and2 I772_270(w_772_272, w_077_240, w_772_271);
  or2  I772_271(w_772_273, w_429_236, w_772_272);
  and2 I772_272(w_772_274, w_772_273, w_446_025);
  not1 I772_273(w_772_265, w_772_274);
  nand2 I772_274(w_772_279, w_701_033, w_772_278);
  not1 I772_275(w_772_280, w_772_279);
  and2 I772_276(w_772_281, w_584_544, w_772_280);
  not1 I772_277(w_772_278, w_772_267);
  and2 I772_278(w_772_283, w_216_352, w_772_281);
  nand2 I773_230(w_773_231, w_773_230, w_381_284);
  or2  I773_231(w_773_232, w_773_231, w_598_028);
  or2  I773_232(w_773_233, w_514_083, w_773_232);
  or2  I773_233(w_773_234, w_214_175, w_773_233);
  nand2 I773_234(w_773_235, w_773_234, w_682_399);
  and2 I773_235(w_773_236, w_731_181, w_773_235);
  not1 I773_236(w_773_230, w_773_236);
  nand2 I774_008(w_774_008, w_397_092, w_360_414);
  and2 I775_193(w_775_193, w_294_031, w_462_524);
  not1 I776_012(w_776_012, w_596_405);
  nand2 I776_102(w_776_102, w_217_054, w_058_206);
  or2  I777_101(w_777_101, w_552_006, w_577_485);
  or2  I778_006(w_778_006, w_583_075, w_499_573);
  nand2 I779_209(w_779_209, w_693_031, w_483_777);
  not1 I779_213(w_779_213, w_749_059);
  nand2 I780_023(w_780_023, w_418_048, w_127_044);
  or2  I781_000(w_781_000, w_104_000, w_271_021);
  not1 I782_041(w_782_041, w_103_199);
  and2 I782_320(w_782_320, w_322_008, w_077_089);
  not1 I783_159(w_783_159, w_724_391);
  nand2 I783_184(w_783_184, w_310_165, w_068_009);
  nand2 I783_235(w_783_235, w_502_472, w_209_281);
  nand2 I784_109(w_784_109, w_383_092, w_547_031);
  or2  I784_272(w_784_272, w_371_000, w_405_182);
  or2  I784_375(w_784_375, w_432_313, w_675_252);
  not1 I784_522(w_784_524, w_784_523);
  and2 I784_523(w_784_525, w_784_534, w_784_524);
  not1 I784_524(w_784_523, w_784_525);
  not1 I784_525(w_784_530, w_784_529);
  and2 I784_526(w_784_531, w_633_039, w_784_530);
  and2 I784_527(w_784_532, w_784_531, w_782_041);
  not1 I784_528(w_784_529, w_784_525);
  and2 I784_529(w_784_534, w_703_220, w_784_532);
  or2  I784_530(w_784_537, w_784_536, w_423_075);
  nand2 I784_531(w_784_538, w_784_537, w_502_349);
  and2 I784_532(w_784_539, w_246_520, w_784_538);
  and2 I784_533(w_784_540, w_784_539, w_314_204);
  nand2 I784_534(w_784_541, w_784_540, w_719_004);
  not1 I784_535(w_784_542, w_784_541);
  not1 I784_536(w_784_543, w_784_542);
  and2 I784_537(w_784_544, w_209_140, w_784_543);
  and2 I784_538(w_784_545, w_784_544, w_161_121);
  nand2 I784_539(w_784_546, w_784_545, w_756_003);
  and2 I784_540(w_784_547, w_401_205, w_784_546);
  nand2 I784_541(w_784_536, w_784_547, w_339_028);
  not1 I785_011(w_785_011, w_232_103);
  and2 I786_008(w_786_008, w_210_124, w_075_116);
  and2 I786_009(w_786_009, w_661_049, w_312_363);
  and2 I787_032(w_787_032, w_487_002, w_215_139);
  and2 I788_008(w_788_008, w_538_046, w_731_147);
  and2 I788_021(w_788_021, w_383_450, w_129_293);
  and2 I788_095(w_788_095, w_326_179, w_605_212);
  or2  I788_134(w_788_134, w_258_153, w_354_004);
  nand2 I788_145(w_788_145, w_077_021, w_274_188);
  or2  I789_050(w_789_050, w_269_030, w_224_114);
  and2 I789_143(w_789_143, w_251_081, w_498_619);
  nand2 I789_340(w_789_340, w_670_022, w_536_022);
  nand2 I790_120(w_790_120, w_399_285, w_691_139);
  and2 I790_123(w_790_123, w_686_107, w_122_082);
  nand2 I790_297(w_790_297, w_772_073, w_584_574);
  and2 I790_401(w_790_401, w_577_031, w_658_094);
  and2 I791_006(w_791_006, w_107_349, w_711_030);
  and2 I792_343(w_792_343, w_206_070, w_479_325);
  not1 I793_014(w_793_014, w_630_049);
  or2  I793_040(w_793_040, w_339_012, w_214_225);
  nand2 I793_053(w_793_053, w_748_267, w_613_009);
  and2 I794_102(w_794_102, w_355_079, w_004_375);
  not1 I795_180(w_795_180, w_464_118);
  not1 I797_003(w_797_003, w_004_109);
  not1 I799_000(w_799_000, w_060_148);
  and2 I800_000(w_800_000, w_067_273, w_079_052);
  or2  I800_001(w_800_001, w_187_004, w_241_033);
  or2  I800_002(w_800_002, w_515_094, w_693_324);
  or2  I800_003(w_800_003, w_017_553, w_709_559);
  or2  I800_004(w_800_004, w_551_031, w_223_235);
  and2 I800_005(w_800_005, w_129_282, w_436_410);
  nand2 I800_006(w_800_006, w_405_073, w_748_126);
  not1 I800_007(w_800_007, w_465_224);
  and2 I800_008(w_800_008, w_259_345, w_341_774);
  nand2 I800_009(w_800_009, w_235_070, w_120_604);
  nand2 I800_010(w_800_010, w_029_009, w_565_009);
  not1 I800_011(w_800_011, w_788_021);
  not1 I800_012(w_800_012, w_117_048);
  not1 I800_013(w_800_013, w_079_027);
  nand2 I800_014(w_800_014, w_557_167, w_560_543);
  and2 I800_015(w_800_015, w_784_109, w_443_327);
  and2 I800_016(w_800_016, w_417_120, w_407_267);
  and2 I800_017(w_800_017, w_211_033, w_022_126);
  and2 I800_018(w_800_018, w_155_072, w_776_012);
  not1 I800_019(w_800_019, w_446_152);
  or2  I800_020(w_800_020, w_525_095, w_300_010);
  not1 I800_021(w_800_021, w_060_326);
  nand2 I800_022(w_800_022, w_396_065, w_718_277);
  or2  I800_023(w_800_023, w_688_501, w_692_155);
  not1 I800_024(w_800_024, w_456_127);
  and2 I800_025(w_800_025, w_134_230, w_575_207);
  nand2 I800_026(w_800_026, w_587_313, w_693_292);
  not1 I800_027(w_800_027, w_770_055);
  nand2 I800_028(w_800_028, w_605_658, w_451_240);
  or2  I800_029(w_800_029, w_048_015, w_403_325);
  and2 I800_030(w_800_030, w_291_099, w_024_219);
  or2  I800_031(w_800_031, w_480_057, w_045_167);
  and2 I800_032(w_800_032, w_620_002, w_095_051);
  nand2 I800_033(w_800_033, w_340_011, w_330_016);
  nand2 I800_034(w_800_034, w_369_115, w_677_020);
  not1 I800_035(w_800_035, w_362_420);
  or2  I800_036(w_800_036, w_317_298, w_629_161);
  or2  I800_037(w_800_037, w_653_063, w_302_049);
  or2  I800_038(w_800_038, w_347_053, w_641_063);
  nand2 I800_039(w_800_039, w_288_478, w_218_180);
  not1 I800_040(w_800_040, w_548_060);
  or2  I800_041(w_800_041, w_469_062, w_530_042);
  and2 I800_042(w_800_042, w_444_462, w_057_313);
  and2 I800_043(w_800_043, w_686_026, w_189_092);
  not1 I800_044(w_800_044, w_491_040);
  and2 I800_045(w_800_045, w_390_031, w_725_102);
  not1 I800_046(w_800_046, w_566_094);
  and2 I800_047(w_800_047, w_746_141, w_233_378);
  nand2 I800_048(w_800_048, w_702_148, w_357_296);
  and2 I800_049(w_800_049, w_353_311, w_118_030);
  nand2 I800_050(w_800_050, w_356_003, w_013_448);
  nand2 I800_051(w_800_051, w_056_037, w_515_066);
  or2  I800_052(w_800_052, w_793_040, w_723_559);
  and2 I800_053(w_800_053, w_056_057, w_126_095);
  nand2 I800_054(w_800_054, w_753_543, w_195_148);
  and2 I800_055(w_800_055, w_255_103, w_351_051);
  not1 I800_056(w_800_056, w_174_060);
  nand2 I800_057(w_800_057, w_187_030, w_310_244);
  or2  I800_058(w_800_058, w_378_112, w_622_074);
  nand2 I800_059(w_800_059, w_098_055, w_056_154);
  nand2 I800_060(w_800_060, w_534_011, w_586_040);
  not1 I800_061(w_800_061, w_781_000);
  not1 I800_062(w_800_062, w_589_022);
  or2  I800_063(w_800_063, w_514_456, w_656_348);
  nand2 I800_064(w_800_064, w_395_229, w_645_314);
  and2 I800_065(w_800_065, w_223_145, w_618_048);
  not1 I800_066(w_800_066, w_716_018);
  not1 I800_067(w_800_067, w_422_001);
  and2 I800_068(w_800_068, w_417_050, w_424_156);
  and2 I800_069(w_800_069, w_679_286, w_725_342);
  and2 I800_070(w_800_070, w_791_006, w_176_170);
  and2 I800_071(w_800_071, w_571_075, w_089_155);
  nand2 I800_072(w_800_072, w_313_397, w_689_227);
  nand2 I800_073(w_800_073, w_158_003, w_233_169);
  and2 I800_074(w_800_074, w_618_060, w_458_060);
  not1 I800_075(w_800_075, w_594_121);
  and2 I800_076(w_800_076, w_071_022, w_064_069);
  nand2 I800_077(w_800_077, w_240_109, w_623_364);
  not1 I800_078(w_800_078, w_265_327);
  or2  I800_079(w_800_079, w_578_724, w_342_103);
  and2 I800_080(w_800_080, w_052_006, w_797_003);
  or2  I800_081(w_800_081, w_615_033, w_744_058);
  or2  I800_082(w_800_082, w_090_531, w_641_058);
  not1 I800_083(w_800_083, w_258_481);
  or2  I800_084(w_800_084, w_498_120, w_213_414);
  not1 I800_085(w_800_085, w_478_335);
  nand2 I800_086(w_800_086, w_608_218, w_269_159);
  not1 I800_087(w_800_087, w_322_002);
  nand2 I800_088(w_800_088, w_507_016, w_147_050);
  and2 I800_089(w_800_089, w_557_111, w_155_288);
  and2 I800_090(w_800_090, w_669_261, w_638_350);
  and2 I800_091(w_800_091, w_689_226, w_549_047);
  and2 I800_092(w_800_092, w_227_597, w_539_387);
  nand2 I800_093(w_800_093, w_008_336, w_349_060);
  nand2 I800_094(w_800_094, w_680_105, w_484_379);
  nand2 I800_095(w_800_095, w_196_136, w_474_202);
  or2  I800_096(w_800_096, w_407_572, w_723_597);
  not1 I800_097(w_800_097, w_259_038);
  and2 I800_098(w_800_098, w_008_246, w_528_015);
  nand2 I800_099(w_800_099, w_267_216, w_762_253);
  nand2 I800_100(w_800_100, w_663_094, w_682_543);
  and2 I800_101(w_800_101, w_718_123, w_035_083);
  nand2 I800_102(w_800_102, w_062_370, w_140_021);
  nand2 I800_103(w_800_103, w_064_170, w_169_218);
  or2  I800_104(w_800_104, w_086_236, w_007_166);
  nand2 I800_105(w_800_105, w_402_114, w_102_364);
  not1 I800_106(w_800_106, w_517_227);
  and2 I800_107(w_800_107, w_751_322, w_424_222);
  or2  I800_108(w_800_108, w_012_338, w_609_050);
  nand2 I800_109(w_800_109, w_301_121, w_306_041);
  or2  I800_110(w_800_110, w_028_006, w_730_150);
  or2  I800_111(w_800_111, w_737_012, w_404_339);
  not1 I800_112(w_800_112, w_058_255);
  and2 I800_113(w_800_113, w_127_034, w_405_027);
  or2  I800_114(w_800_114, w_381_653, w_706_227);
  not1 I800_115(w_800_115, w_067_371);
  or2  I800_116(w_800_116, w_369_722, w_564_007);
  and2 I800_117(w_800_117, w_144_079, w_374_091);
  and2 I800_118(w_800_118, w_312_355, w_417_065);
  or2  I800_119(w_800_119, w_475_011, w_245_155);
  or2  I800_120(w_800_120, w_202_276, w_754_136);
  nand2 I800_121(w_800_121, w_661_018, w_533_110);
  or2  I800_122(w_800_122, w_790_297, w_727_106);
  and2 I800_123(w_800_123, w_371_000, w_215_206);
  and2 I800_124(w_800_124, w_676_258, w_407_293);
  or2  I800_125(w_800_125, w_572_131, w_024_017);
  nand2 I800_126(w_800_126, w_070_572, w_613_024);
  and2 I800_127(w_800_127, w_604_237, w_789_050);
  not1 I800_128(w_800_128, w_346_076);
  nand2 I800_129(w_800_129, w_626_338, w_599_032);
  or2  I800_130(w_800_130, w_015_143, w_553_027);
  or2  I800_131(w_800_131, w_512_088, w_767_284);
  and2 I800_132(w_800_132, w_791_006, w_788_095);
  not1 I800_133(w_800_133, w_601_123);
  not1 I800_134(w_800_134, w_758_227);
  nand2 I800_135(w_800_135, w_647_393, w_126_079);
  or2  I800_136(w_800_136, w_752_418, w_560_149);
  nand2 I800_137(w_800_137, w_575_053, w_664_018);
  not1 I800_138(w_800_138, w_377_013);
  or2  I800_139(w_800_139, w_213_419, w_557_419);
  nand2 I800_140(w_800_140, w_522_397, w_560_512);
  nand2 I800_141(w_800_141, w_518_010, w_063_366);
  or2  I800_142(w_800_142, w_189_445, w_198_062);
  nand2 I800_143(w_800_143, w_759_642, w_174_090);
  nand2 I800_144(w_800_144, w_391_105, w_382_033);
  nand2 I800_145(w_800_145, w_147_037, w_182_013);
  or2  I800_146(w_800_146, w_589_331, w_454_340);
  nand2 I800_147(w_800_147, w_290_106, w_687_198);
  not1 I800_148(w_800_148, w_125_446);
  and2 I800_149(w_800_149, w_323_139, w_751_282);
  or2  I800_150(w_800_150, w_126_175, w_117_057);
  not1 I800_151(w_800_151, w_051_037);
  or2  I800_152(w_800_152, w_550_122, w_324_029);
  nand2 I800_153(w_800_153, w_465_014, w_282_367);
  or2  I800_154(w_800_154, w_124_116, w_525_029);
  not1 I800_155(w_800_155, w_202_165);
  not1 I800_156(w_800_156, w_077_166);
  not1 I800_157(w_800_157, w_712_033);
  and2 I800_158(w_800_158, w_281_616, w_361_249);
  nand2 I800_159(w_800_159, w_750_448, w_770_072);
  and2 I800_160(w_800_160, w_681_252, w_790_123);
  not1 I800_161(w_800_161, w_357_408);
  not1 I800_162(w_800_162, w_697_033);
  nand2 I800_163(w_800_163, w_576_111, w_266_438);
  or2  I800_164(w_800_164, w_432_288, w_677_131);
  and2 I800_165(w_800_165, w_510_748, w_009_369);
  nand2 I800_166(w_800_166, w_311_369, w_489_384);
  not1 I800_167(w_800_167, w_370_084);
  and2 I800_168(w_800_168, w_493_093, w_145_039);
  and2 I800_169(w_800_169, w_043_043, w_275_619);
  nand2 I800_170(w_800_170, w_093_050, w_344_077);
  not1 I800_171(w_800_171, w_573_208);
  not1 I800_172(w_800_172, w_635_156);
  and2 I800_173(w_800_173, w_556_324, w_287_125);
  or2  I800_174(w_800_174, w_671_371, w_736_059);
  nand2 I800_175(w_800_175, w_429_115, w_305_083);
  or2  I800_176(w_800_176, w_348_213, w_196_254);
  not1 I800_177(w_800_177, w_641_072);
  not1 I800_178(w_800_178, w_718_646);
  nand2 I800_179(w_800_179, w_127_027, w_362_193);
  or2  I800_180(w_800_180, w_118_087, w_524_595);
  or2  I800_181(w_800_181, w_748_161, w_013_359);
  not1 I800_182(w_800_182, w_442_104);
  nand2 I800_183(w_800_183, w_078_166, w_083_008);
  nand2 I800_184(w_800_184, w_154_051, w_556_035);
  or2  I800_185(w_800_185, w_027_066, w_488_018);
  not1 I800_186(w_800_186, w_402_021);
  nand2 I800_187(w_800_187, w_520_053, w_360_315);
  not1 I800_188(w_800_188, w_308_034);
  nand2 I800_189(w_800_189, w_219_265, w_137_464);
  and2 I800_190(w_800_190, w_567_042, w_084_030);
  not1 I800_191(w_800_191, w_238_235);
  not1 I800_192(w_800_192, w_625_100);
  or2  I800_193(w_800_193, w_059_140, w_739_105);
  not1 I800_194(w_800_194, w_281_389);
  not1 I800_195(w_800_195, w_686_011);
  not1 I800_196(w_800_196, w_016_006);
  and2 I800_197(w_800_197, w_511_028, w_781_000);
  or2  I800_198(w_800_198, w_782_320, w_228_066);
  and2 I800_199(w_800_199, w_678_201, w_432_120);
  not1 I800_200(w_800_200, w_532_222);
  or2  I800_201(w_800_201, w_673_161, w_198_056);
  not1 I800_202(w_800_202, w_587_230);
  and2 I800_203(w_800_203, w_536_040, w_600_697);
  and2 I800_204(w_800_204, w_311_263, w_410_064);
  nand2 I800_205(w_800_205, w_392_185, w_199_048);
  and2 I800_206(w_800_206, w_429_096, w_564_065);
  and2 I800_207(w_800_207, w_649_026, w_793_014);
  or2  I800_208(w_800_208, w_192_041, w_347_331);
  nand2 I800_209(w_800_209, w_580_420, w_535_119);
  or2  I800_210(w_800_210, w_164_244, w_243_268);
  and2 I800_211(w_800_211, w_214_166, w_596_137);
  and2 I800_212(w_800_212, w_728_394, w_042_036);
  and2 I800_213(w_800_213, w_295_247, w_299_288);
  and2 I800_214(w_800_214, w_652_042, w_361_200);
  and2 I800_215(w_800_215, w_537_029, w_784_272);
  and2 I800_216(w_800_216, w_301_210, w_156_545);
  not1 I800_217(w_800_217, w_016_005);
  and2 I800_218(w_800_218, w_612_103, w_456_039);
  nand2 I800_219(w_800_219, w_051_171, w_235_056);
  and2 I800_220(w_800_220, w_087_186, w_352_314);
  nand2 I800_221(w_800_221, w_265_491, w_583_002);
  nand2 I800_222(w_800_222, w_567_040, w_288_068);
  nand2 I800_223(w_800_223, w_444_165, w_026_013);
  or2  I800_224(w_800_224, w_306_177, w_306_087);
  not1 I800_225(w_800_225, w_529_004);
  and2 I800_226(w_800_226, w_765_198, w_440_032);
  not1 I800_227(w_800_227, w_792_343);
  or2  I800_228(w_800_228, w_610_041, w_100_080);
  not1 I800_229(w_800_229, w_219_439);
  not1 I800_230(w_800_230, w_288_194);
  nand2 I800_231(w_800_231, w_005_281, w_260_201);
  nand2 I800_232(w_800_232, w_789_340, w_550_260);
  not1 I800_233(w_800_233, w_116_030);
  nand2 I800_234(w_800_234, w_028_074, w_343_479);
  or2  I800_235(w_800_235, w_686_102, w_015_625);
  or2  I800_236(w_800_236, w_180_020, w_668_171);
  not1 I800_237(w_800_237, w_508_074);
  or2  I800_238(w_800_238, w_514_170, w_545_117);
  nand2 I800_239(w_800_239, w_535_180, w_245_347);
  nand2 I800_240(w_800_240, w_714_009, w_450_052);
  and2 I800_241(w_800_241, w_793_053, w_186_231);
  not1 I800_242(w_800_242, w_201_057);
  nand2 I800_243(w_800_243, w_733_100, w_543_105);
  nand2 I800_244(w_800_244, w_252_103, w_169_318);
  nand2 I800_245(w_800_245, w_714_046, w_134_001);
  nand2 I800_246(w_800_246, w_731_103, w_122_005);
  and2 I800_247(w_800_247, w_572_140, w_448_117);
  or2  I800_248(w_800_248, w_634_295, w_787_032);
  not1 I800_249(w_800_249, w_662_321);
  nand2 I800_250(w_800_250, w_406_116, w_390_252);
  not1 I800_251(w_800_251, w_559_040);
  or2  I800_252(w_800_252, w_026_146, w_283_379);
  not1 I800_253(w_800_253, w_214_280);
  and2 I800_254(w_800_254, w_412_300, w_453_552);
  and2 I800_255(w_800_255, w_122_089, w_583_023);
  or2  I800_256(w_800_256, w_171_333, w_419_044);
  and2 I800_257(w_800_257, w_025_162, w_783_235);
  or2  I800_258(w_800_258, w_094_101, w_682_472);
  not1 I800_259(w_800_259, w_517_052);
  and2 I800_260(w_800_260, w_731_087, w_548_264);
  and2 I800_261(w_800_261, w_553_015, w_484_296);
  or2  I800_262(w_800_262, w_619_251, w_422_010);
  or2  I800_263(w_800_263, w_393_149, w_177_008);
  not1 I800_264(w_800_264, w_512_098);
  nand2 I800_265(w_800_265, w_607_016, w_025_279);
  and2 I800_266(w_800_266, w_542_331, w_052_025);
  nand2 I800_267(w_800_267, w_152_721, w_303_106);
  and2 I800_268(w_800_268, w_788_134, w_137_098);
  or2  I800_269(w_800_269, w_559_028, w_522_505);
  or2  I800_270(w_800_270, w_252_124, w_147_020);
  not1 I800_271(w_800_271, w_290_100);
  and2 I800_272(w_800_272, w_667_051, w_332_409);
  not1 I800_273(w_800_273, w_736_091);
  not1 I800_274(w_800_274, w_089_259);
  or2  I800_275(w_800_275, w_795_180, w_345_129);
  or2  I800_276(w_800_276, w_505_066, w_429_085);
  or2  I800_277(w_800_277, w_134_256, w_393_020);
  nand2 I800_278(w_800_278, w_357_588, w_733_045);
  or2  I800_279(w_800_279, w_600_084, w_173_017);
  not1 I800_280(w_800_280, w_462_547);
  and2 I800_281(w_800_281, w_551_007, w_334_098);
  nand2 I800_282(w_800_282, w_231_579, w_504_027);
  or2  I800_283(w_800_283, w_485_143, w_786_009);
  nand2 I800_284(w_800_284, w_731_077, w_178_076);
  not1 I800_285(w_800_285, w_463_119);
  nand2 I800_286(w_800_286, w_263_083, w_584_024);
  and2 I800_287(w_800_287, w_246_124, w_305_178);
  nand2 I800_288(w_800_288, w_191_076, w_222_422);
  not1 I800_289(w_800_289, w_278_045);
  and2 I800_290(w_800_290, w_764_054, w_410_027);
  not1 I800_291(w_800_291, w_342_213);
  and2 I800_292(w_800_292, w_535_000, w_336_057);
  not1 I800_293(w_800_293, w_151_367);
  not1 I800_294(w_800_294, w_528_039);
  or2  I800_295(w_800_295, w_652_041, w_774_008);
  nand2 I800_296(w_800_296, w_422_002, w_718_200);
  nand2 I800_297(w_800_297, w_629_624, w_351_235);
  nand2 I800_298(w_800_298, w_135_377, w_481_042);
  not1 I800_299(w_800_299, w_216_262);
  not1 I800_300(w_800_300, w_625_277);
  or2  I800_301(w_800_301, w_192_065, w_017_439);
  and2 I800_302(w_800_302, w_221_018, w_759_108);
  nand2 I800_303(w_800_303, w_733_108, w_757_133);
  or2  I800_304(w_800_304, w_138_310, w_156_374);
  or2  I800_305(w_800_305, w_643_303, w_578_543);
  or2  I800_306(w_800_306, w_794_102, w_595_130);
  nand2 I800_307(w_800_307, w_085_011, w_263_049);
  not1 I800_308(w_800_308, w_695_052);
  not1 I800_309(w_800_309, w_654_336);
  not1 I800_310(w_800_310, w_139_022);
  nand2 I800_311(w_800_311, w_273_093, w_586_125);
  nand2 I800_312(w_800_312, w_512_124, w_359_015);
  not1 I800_313(w_800_313, w_454_111);
  and2 I800_314(w_800_314, w_433_268, w_175_240);
  or2  I800_315(w_800_315, w_538_039, w_360_021);
  nand2 I800_316(w_800_316, w_588_111, w_157_124);
  or2  I800_317(w_800_317, w_297_116, w_072_122);
  or2  I800_318(w_800_318, w_210_107, w_305_103);
  or2  I800_319(w_800_319, w_216_290, w_499_222);
  nand2 I800_320(w_800_320, w_055_309, w_231_001);
  and2 I800_321(w_800_321, w_137_320, w_503_015);
  and2 I800_322(w_800_322, w_006_131, w_251_028);
  or2  I800_323(w_800_323, w_228_013, w_640_653);
  nand2 I800_324(w_800_324, w_429_130, w_744_072);
  not1 I800_325(w_800_325, w_433_054);
  and2 I800_326(w_800_326, w_484_277, w_495_096);
  and2 I800_327(w_800_327, w_726_165, w_132_415);
  or2  I800_328(w_800_328, w_636_112, w_157_135);
  or2  I800_329(w_800_329, w_761_018, w_263_001);
  nand2 I800_330(w_800_330, w_455_112, w_762_061);
  not1 I800_331(w_800_331, w_706_205);
  and2 I800_332(w_800_332, w_691_005, w_784_375);
  not1 I800_333(w_800_333, w_479_107);
  nand2 I800_334(w_800_334, w_405_137, w_423_021);
  and2 I800_335(w_800_335, w_611_485, w_242_006);
  nand2 I800_336(w_800_336, w_203_198, w_602_296);
  and2 I800_337(w_800_337, w_257_243, w_154_033);
  or2  I800_338(w_800_338, w_061_168, w_409_304);
  not1 I800_339(w_800_339, w_393_204);
  and2 I800_340(w_800_340, w_072_098, w_595_029);
  not1 I800_341(w_800_341, w_571_402);
  not1 I800_342(w_800_342, w_734_104);
  and2 I800_343(w_800_343, w_740_318, w_223_209);
  or2  I800_344(w_800_344, w_520_109, w_038_140);
  nand2 I800_345(w_800_345, w_283_131, w_168_452);
  or2  I800_346(w_800_346, w_473_502, w_122_065);
  not1 I800_347(w_800_347, w_546_086);
  not1 I800_348(w_800_348, w_127_043);
  or2  I800_349(w_800_349, w_082_027, w_211_036);
  and2 I800_350(w_800_350, w_504_053, w_512_157);
  not1 I800_351(w_800_351, w_584_666);
  and2 I800_352(w_800_352, w_547_045, w_059_667);
  not1 I800_353(w_800_353, w_511_396);
  nand2 I800_354(w_800_354, w_213_070, w_072_272);
  and2 I800_355(w_800_355, w_227_278, w_295_173);
  nand2 I800_356(w_800_356, w_377_066, w_670_024);
  or2  I800_357(w_800_357, w_374_056, w_697_187);
  not1 I800_358(w_800_358, w_481_057);
  not1 I800_359(w_800_359, w_580_031);
  not1 I800_360(w_800_360, w_447_173);
  or2  I800_361(w_800_361, w_043_004, w_355_113);
  and2 I800_362(w_800_362, w_479_281, w_191_309);
  or2  I800_363(w_800_363, w_716_029, w_506_261);
  not1 I800_364(w_800_364, w_510_447);
  or2  I800_365(w_800_365, w_118_060, w_404_361);
  not1 I800_366(w_800_366, w_462_379);
  not1 I800_367(w_800_367, w_493_095);
  not1 I800_368(w_800_368, w_218_599);
  or2  I800_369(w_800_369, w_558_122, w_219_522);
  or2  I800_370(w_800_370, w_052_030, w_398_074);
  not1 I800_371(w_800_371, w_014_240);
  nand2 I800_372(w_800_372, w_652_020, w_442_135);
  and2 I800_373(w_800_373, w_339_022, w_781_000);
  and2 I800_374(w_800_374, w_361_369, w_529_000);
  or2  I800_375(w_800_375, w_747_019, w_243_057);
  nand2 I800_376(w_800_376, w_014_282, w_316_066);
  and2 I800_377(w_800_377, w_714_000, w_130_280);
  and2 I800_378(w_800_378, w_126_133, w_790_120);
  not1 I800_379(w_800_379, w_410_011);
  and2 I800_380(w_800_380, w_392_081, w_160_753);
  and2 I800_381(w_800_381, w_241_059, w_653_188);
  or2  I800_382(w_800_382, w_448_245, w_528_046);
  and2 I800_383(w_800_383, w_397_081, w_325_005);
  or2  I800_384(w_800_384, w_455_144, w_369_133);
  or2  I800_385(w_800_385, w_711_004, w_731_122);
  or2  I800_386(w_800_386, w_056_713, w_098_043);
  not1 I800_387(w_800_387, w_262_010);
  not1 I800_388(w_800_388, w_467_181);
  nand2 I800_389(w_800_389, w_116_348, w_571_130);
  and2 I800_390(w_800_390, w_168_014, w_601_384);
  and2 I800_391(w_800_391, w_257_190, w_365_390);
  or2  I800_392(w_800_392, w_276_196, w_640_598);
  not1 I800_393(w_800_393, w_248_063);
  and2 I800_394(w_800_394, w_369_282, w_726_379);
  and2 I800_395(w_800_395, w_393_129, w_323_061);
  or2  I800_396(w_800_396, w_446_544, w_754_167);
  nand2 I800_397(w_800_397, w_107_125, w_304_178);
  nand2 I800_398(w_800_398, w_669_307, w_188_146);
  nand2 I800_399(w_800_399, w_380_296, w_069_181);
  nand2 I800_400(w_800_400, w_533_550, w_193_106);
  or2  I800_401(w_800_401, w_121_190, w_610_104);
  not1 I800_402(w_800_402, w_640_443);
  not1 I800_403(w_800_403, w_146_285);
  not1 I800_404(w_800_404, w_253_361);
  not1 I800_405(w_800_405, w_170_209);
  nand2 I800_406(w_800_406, w_029_026, w_293_084);
  and2 I800_407(w_800_407, w_589_154, w_493_139);
  nand2 I800_408(w_800_408, w_595_246, w_699_724);
  and2 I800_409(w_800_409, w_656_087, w_716_029);
  nand2 I800_410(w_800_410, w_359_021, w_073_169);
  nand2 I800_411(w_800_411, w_326_114, w_337_004);
  not1 I800_412(w_800_412, w_132_077);
  not1 I800_413(w_800_413, w_426_162);
  nand2 I800_414(w_800_414, w_567_010, w_212_162);
  nand2 I800_415(w_800_415, w_008_067, w_358_284);
  nand2 I800_416(w_800_416, w_214_371, w_255_089);
  not1 I800_417(w_800_417, w_615_078);
  nand2 I800_418(w_800_418, w_336_235, w_602_005);
  not1 I800_419(w_800_419, w_650_341);
  not1 I800_420(w_800_420, w_728_548);
  and2 I800_421(w_800_421, w_442_126, w_256_310);
  nand2 I800_422(w_800_422, w_076_277, w_039_495);
  and2 I800_423(w_800_423, w_676_185, w_094_599);
  not1 I800_424(w_800_424, w_535_189);
  or2  I800_425(w_800_425, w_613_089, w_441_023);
  nand2 I800_426(w_800_426, w_060_277, w_730_122);
  nand2 I800_427(w_800_427, w_658_054, w_079_044);
  or2  I800_428(w_800_428, w_335_162, w_704_043);
  nand2 I800_429(w_800_429, w_296_032, w_011_172);
  not1 I800_430(w_800_430, w_106_116);
  and2 I800_431(w_800_431, w_193_067, w_441_007);
  nand2 I800_432(w_800_432, w_082_213, w_330_201);
  not1 I800_433(w_800_433, w_260_001);
  or2  I800_434(w_800_434, w_470_407, w_468_154);
  and2 I800_435(w_800_435, w_004_484, w_184_052);
  and2 I800_436(w_800_436, w_480_107, w_179_204);
  or2  I800_437(w_800_437, w_637_242, w_361_031);
  or2  I800_438(w_800_438, w_002_390, w_304_437);
  nand2 I800_439(w_800_439, w_635_484, w_249_069);
  or2  I800_440(w_800_440, w_638_470, w_444_307);
  and2 I800_441(w_800_441, w_724_311, w_029_108);
  nand2 I800_442(w_800_442, w_197_141, w_514_191);
  or2  I800_443(w_800_443, w_540_118, w_777_101);
  or2  I800_444(w_800_444, w_031_456, w_091_144);
  or2  I800_445(w_800_445, w_246_074, w_577_496);
  not1 I800_446(w_800_446, w_614_334);
  and2 I800_447(w_800_447, w_258_193, w_184_132);
  and2 I800_448(w_800_448, w_213_194, w_239_000);
  nand2 I800_449(w_800_449, w_754_167, w_585_046);
  or2  I800_450(w_800_450, w_562_147, w_062_593);
  nand2 I800_451(w_800_451, w_505_236, w_248_111);
  nand2 I800_452(w_800_452, w_025_181, w_629_191);
  not1 I800_453(w_800_453, w_373_001);
  nand2 I800_454(w_800_454, w_558_151, w_136_063);
  not1 I800_455(w_800_455, w_375_071);
  or2  I800_456(w_800_456, w_681_081, w_402_087);
  not1 I800_457(w_800_457, w_165_105);
  and2 I800_458(w_800_458, w_310_582, w_561_343);
  nand2 I800_459(w_800_459, w_512_451, w_408_004);
  and2 I800_460(w_800_460, w_152_007, w_654_153);
  or2  I800_461(w_800_461, w_764_241, w_517_005);
  nand2 I800_462(w_800_462, w_445_029, w_788_008);
  not1 I800_463(w_800_463, w_743_021);
  and2 I800_464(w_800_464, w_460_233, w_608_359);
  nand2 I800_465(w_800_465, w_369_666, w_750_434);
  or2  I800_466(w_800_466, w_711_048, w_149_063);
  and2 I800_467(w_800_467, w_003_058, w_381_319);
  or2  I800_468(w_800_468, w_451_217, w_180_015);
  and2 I800_469(w_800_469, w_521_058, w_651_464);
  and2 I800_470(w_800_470, w_755_016, w_717_116);
  not1 I800_471(w_800_471, w_285_037);
  and2 I800_472(w_800_472, w_235_181, w_629_146);
  or2  I800_473(w_800_473, w_779_209, w_521_334);
  not1 I800_474(w_800_474, w_103_206);
  nand2 I800_475(w_800_475, w_106_096, w_520_202);
  or2  I800_476(w_800_476, w_241_000, w_660_001);
  or2  I800_477(w_800_477, w_168_381, w_578_284);
  nand2 I800_478(w_800_478, w_063_113, w_692_168);
  or2  I800_479(w_800_479, w_073_055, w_418_052);
  nand2 I800_480(w_800_480, w_492_275, w_089_291);
  or2  I800_481(w_800_481, w_780_023, w_414_151);
  nand2 I800_482(w_800_482, w_423_073, w_535_114);
  not1 I800_483(w_800_483, w_396_004);
  nand2 I800_484(w_800_484, w_527_061, w_063_142);
  or2  I800_485(w_800_485, w_307_305, w_410_102);
  nand2 I800_486(w_800_486, w_381_104, w_454_073);
  and2 I800_487(w_800_487, w_095_043, w_421_075);
  or2  I800_488(w_800_488, w_035_000, w_128_010);
  or2  I800_489(w_800_489, w_215_106, w_524_612);
  not1 I800_490(w_800_490, w_207_119);
  not1 I800_491(w_800_491, w_622_033);
  and2 I800_492(w_800_492, w_481_050, w_518_062);
  not1 I800_493(w_800_493, w_099_047);
  and2 I800_494(w_800_494, w_172_048, w_023_090);
  and2 I800_495(w_800_495, w_450_175, w_331_072);
  or2  I800_496(w_800_496, w_693_163, w_313_090);
  and2 I800_497(w_800_497, w_125_150, w_035_112);
  or2  I800_498(w_800_498, w_210_101, w_093_132);
  and2 I800_499(w_800_499, w_163_159, w_254_095);
  and2 I800_500(w_800_500, w_534_003, w_675_109);
  and2 I800_501(w_800_501, w_171_560, w_701_054);
  not1 I800_502(w_800_502, w_799_000);
  not1 I800_503(w_800_503, w_312_040);
  not1 I800_504(w_800_504, w_789_143);
  not1 I800_505(w_800_505, w_357_319);
  and2 I800_506(w_800_506, w_310_412, w_407_643);
  and2 I800_507(w_800_507, w_361_097, w_743_031);
  and2 I800_508(w_800_508, w_282_141, w_293_033);
  and2 I800_509(w_800_509, w_053_020, w_719_150);
  nand2 I800_510(w_800_510, w_219_738, w_683_259);
  or2  I800_511(w_800_511, w_224_241, w_163_133);
  or2  I800_512(w_800_512, w_679_443, w_077_286);
  not1 I800_513(w_800_513, w_205_199);
  and2 I800_514(w_800_514, w_148_017, w_120_042);
  not1 I800_515(w_800_515, w_413_015);
  not1 I800_516(w_800_516, w_019_002);
  or2  I800_517(w_800_517, w_315_140, w_064_253);
  nand2 I800_518(w_800_518, w_323_123, w_599_018);
  or2  I800_519(w_800_519, w_732_016, w_408_002);
  nand2 I800_520(w_800_520, w_247_142, w_065_098);
  not1 I800_521(w_800_521, w_213_015);
  not1 I800_522(w_800_522, w_196_173);
  and2 I800_523(w_800_523, w_298_100, w_159_065);
  or2  I800_524(w_800_524, w_026_112, w_010_631);
  nand2 I800_525(w_800_525, w_685_294, w_639_018);
  nand2 I800_526(w_800_526, w_123_584, w_432_051);
  and2 I800_527(w_800_527, w_679_618, w_509_075);
  and2 I800_528(w_800_528, w_274_171, w_399_023);
  not1 I800_529(w_800_529, w_539_321);
  not1 I800_530(w_800_530, w_250_292);
  and2 I800_531(w_800_531, w_276_296, w_378_107);
  and2 I800_532(w_800_532, w_263_078, w_635_170);
  or2  I800_533(w_800_533, w_310_061, w_761_022);
  not1 I800_534(w_800_534, w_640_532);
  nand2 I800_535(w_800_535, w_069_218, w_286_362);
  nand2 I800_536(w_800_536, w_309_352, w_094_182);
  nand2 I800_537(w_800_537, w_344_026, w_019_004);
  nand2 I800_538(w_800_538, w_397_048, w_779_213);
  or2  I800_539(w_800_539, w_166_056, w_114_020);
  or2  I800_540(w_800_540, w_075_076, w_640_267);
  not1 I800_541(w_800_541, w_651_337);
  nand2 I800_542(w_800_542, w_489_025, w_786_008);
  and2 I800_543(w_800_543, w_433_180, w_588_153);
  nand2 I800_544(w_800_544, w_159_030, w_542_061);
  not1 I800_545(w_800_545, w_521_322);
  nand2 I800_546(w_800_546, w_687_198, w_138_061);
  not1 I800_547(w_800_547, w_565_020);
  not1 I800_548(w_800_548, w_033_428);
  not1 I800_549(w_800_549, w_370_099);
  nand2 I800_550(w_800_550, w_573_020, w_230_038);
  nand2 I800_551(w_800_551, w_762_123, w_712_065);
  or2  I800_552(w_800_552, w_766_300, w_414_303);
  and2 I800_553(w_800_553, w_288_167, w_575_065);
  not1 I800_554(w_800_554, w_491_077);
  nand2 I800_555(w_800_555, w_349_230, w_516_329);
  and2 I800_556(w_800_556, w_438_253, w_556_212);
  nand2 I800_557(w_800_557, w_338_239, w_274_130);
  and2 I800_558(w_800_558, w_538_262, w_477_057);
  or2  I800_559(w_800_559, w_444_709, w_430_060);
  or2  I800_560(w_800_560, w_557_050, w_055_254);
  not1 I800_561(w_800_561, w_187_023);
  and2 I800_562(w_800_562, w_703_135, w_477_030);
  and2 I800_563(w_800_563, w_585_554, w_311_123);
  and2 I800_564(w_800_564, w_137_266, w_496_077);
  or2  I800_565(w_800_565, w_173_028, w_443_263);
  not1 I800_566(w_800_566, w_425_102);
  nand2 I800_567(w_800_567, w_182_013, w_739_093);
  not1 I800_568(w_800_568, w_478_078);
  not1 I800_569(w_800_569, w_381_163);
  nand2 I800_570(w_800_570, w_275_135, w_020_381);
  not1 I800_571(w_800_571, w_143_257);
  nand2 I800_572(w_800_572, w_471_074, w_363_372);
  nand2 I800_573(w_800_573, w_647_367, w_648_079);
  and2 I800_574(w_800_574, w_302_629, w_527_082);
  and2 I800_575(w_800_575, w_510_136, w_598_017);
  nand2 I800_576(w_800_576, w_179_710, w_578_007);
  or2  I800_577(w_800_577, w_151_388, w_044_646);
  not1 I800_578(w_800_578, w_531_317);
  nand2 I800_579(w_800_579, w_446_242, w_182_025);
  or2  I800_580(w_800_580, w_383_591, w_154_025);
  and2 I800_581(w_800_581, w_681_320, w_540_053);
  and2 I800_582(w_800_582, w_338_158, w_351_070);
  nand2 I800_583(w_800_583, w_482_077, w_797_003);
  or2  I800_584(w_800_584, w_393_003, w_663_060);
  or2  I800_585(w_800_585, w_367_123, w_591_101);
  or2  I800_586(w_800_586, w_400_024, w_560_106);
  not1 I800_587(w_800_587, w_533_169);
  not1 I800_588(w_800_588, w_273_065);
  not1 I800_589(w_800_589, w_612_076);
  not1 I800_590(w_800_590, w_682_371);
  and2 I800_591(w_800_591, w_759_047, w_021_226);
  or2  I800_592(w_800_592, w_500_274, w_790_401);
  nand2 I800_593(w_800_593, w_465_192, w_308_146);
  or2  I800_594(w_800_594, w_345_098, w_251_131);
  nand2 I800_595(w_800_595, w_239_000, w_457_099);
  nand2 I800_596(w_800_596, w_269_493, w_465_165);
  or2  I800_597(w_800_597, w_301_014, w_689_090);
  not1 I800_598(w_800_598, w_203_375);
  not1 I800_599(w_800_599, w_545_345);
  or2  I800_600(w_800_600, w_210_019, w_250_548);
  not1 I800_601(w_800_601, w_595_157);
  or2  I800_602(w_800_602, w_062_030, w_356_061);
  nand2 I800_603(w_800_603, w_430_114, w_308_155);
  and2 I800_604(w_800_604, w_011_444, w_753_377);
  not1 I800_605(w_800_605, w_276_367);
  or2  I800_606(w_800_606, w_203_032, w_634_179);
  nand2 I800_607(w_800_607, w_396_007, w_741_144);
  not1 I800_608(w_800_608, w_088_048);
  and2 I800_609(w_800_609, w_502_372, w_592_177);
  nand2 I800_610(w_800_610, w_574_164, w_719_250);
  and2 I800_611(w_800_611, w_282_246, w_121_211);
  and2 I800_612(w_800_612, w_749_131, w_669_152);
  or2  I800_613(w_800_613, w_503_202, w_724_451);
  and2 I800_614(w_800_614, w_218_595, w_703_306);
  not1 I800_615(w_800_615, w_587_009);
  not1 I800_616(w_800_616, w_731_186);
  not1 I800_617(w_800_617, w_506_071);
  or2  I800_618(w_800_618, w_756_070, w_132_202);
  and2 I800_619(w_800_619, w_343_335, w_493_026);
  and2 I800_620(w_800_620, w_646_003, w_260_082);
  and2 I800_621(w_800_621, w_711_018, w_402_027);
  or2  I800_622(w_800_622, w_708_064, w_708_269);
  nand2 I800_623(w_800_623, w_640_456, w_541_066);
  not1 I800_624(w_800_624, w_039_206);
  or2  I800_625(w_800_625, w_523_190, w_173_002);
  nand2 I800_626(w_800_626, w_666_445, w_500_064);
  and2 I800_627(w_800_627, w_312_146, w_088_076);
  or2  I800_628(w_800_628, w_042_282, w_038_303);
  nand2 I800_629(w_800_629, w_299_097, w_195_139);
  and2 I800_630(w_800_630, w_736_389, w_139_019);
  nand2 I800_631(w_800_631, w_120_402, w_555_293);
  or2  I800_632(w_800_632, w_051_096, w_466_103);
  and2 I800_633(w_800_633, w_722_415, w_626_011);
  not1 I800_634(w_800_634, w_191_034);
  or2  I800_635(w_800_635, w_582_708, w_056_081);
  or2  I800_636(w_800_636, w_251_028, w_261_000);
  or2  I800_637(w_800_637, w_400_051, w_756_072);
  not1 I800_638(w_800_638, w_511_186);
  nand2 I800_639(w_800_639, w_562_429, w_061_217);
  or2  I800_640(w_800_640, w_783_184, w_735_051);
  nand2 I800_641(w_800_641, w_479_034, w_048_001);
  and2 I800_642(w_800_642, w_104_342, w_693_319);
  not1 I800_643(w_800_643, w_155_000);
  nand2 I800_644(w_800_644, w_107_345, w_231_532);
  or2  I800_645(w_800_645, w_294_145, w_388_057);
  not1 I800_646(w_800_646, w_001_034);
  nand2 I800_647(w_800_647, w_785_011, w_475_057);
  not1 I800_648(w_800_648, w_154_055);
  not1 I800_649(w_800_649, w_415_072);
  not1 I800_650(w_800_650, w_309_264);
  not1 I800_651(w_800_651, w_423_022);
  not1 I800_652(w_800_652, w_250_012);
  not1 I800_653(w_800_653, w_481_215);
  nand2 I800_654(w_800_654, w_775_193, w_608_384);
  and2 I800_655(w_800_655, w_609_187, w_267_146);
  not1 I800_656(w_800_656, w_742_030);
  and2 I800_657(w_800_657, w_448_283, w_498_415);
  or2  I800_658(w_800_658, w_140_001, w_367_491);
  nand2 I800_659(w_800_659, w_719_393, w_149_027);
  nand2 I800_660(w_800_660, w_182_016, w_487_510);
  or2  I800_661(w_800_661, w_647_446, w_397_018);
  or2  I800_662(w_800_662, w_664_155, w_783_159);
  or2  I800_663(w_800_663, w_495_164, w_306_207);
  nand2 I800_664(w_800_664, w_028_099, w_051_395);
  or2  I800_665(w_800_665, w_751_314, w_322_017);
  not1 I800_666(w_800_666, w_142_187);
  or2  I800_667(w_800_667, w_181_153, w_494_028);
  nand2 I800_668(w_800_668, w_443_130, w_553_020);
  nand2 I800_669(w_800_669, w_088_019, w_728_136);
  not1 I800_670(w_800_670, w_235_101);
  or2  I800_671(w_800_671, w_263_119, w_357_658);
  and2 I800_672(w_800_672, w_660_000, w_371_000);
  not1 I800_673(w_800_673, w_513_499);
  and2 I800_674(w_800_674, w_246_107, w_290_117);
  and2 I800_675(w_800_675, w_734_086, w_749_176);
  not1 I800_676(w_800_676, w_389_150);
  not1 I800_677(w_800_677, w_525_029);
  or2  I800_678(w_800_678, w_759_649, w_480_078);
  not1 I800_679(w_800_679, w_690_025);
  not1 I800_680(w_800_680, w_415_050);
  not1 I800_681(w_800_681, w_737_115);
  not1 I800_682(w_800_682, w_533_361);
  not1 I800_683(w_800_683, w_024_055);
  not1 I800_684(w_800_684, w_310_145);
  nand2 I800_685(w_800_685, w_104_199, w_465_269);
  not1 I800_686(w_800_686, w_542_116);
  nand2 I800_687(w_800_687, w_501_013, w_080_132);
  nand2 I800_688(w_800_688, w_322_002, w_637_003);
  or2  I800_689(w_800_689, w_568_227, w_776_102);
  and2 I800_690(w_800_690, w_337_384, w_336_016);
  nand2 I800_691(w_800_691, w_646_013, w_586_073);
  or2  I800_692(w_800_692, w_603_123, w_603_163);
  and2 I800_693(w_800_693, w_202_089, w_301_182);
  nand2 I800_694(w_800_694, w_521_151, w_342_358);
  not1 I800_695(w_800_695, w_203_478);
  or2  I800_696(w_800_696, w_531_580, w_090_420);
  or2  I800_697(w_800_697, w_778_006, w_228_625);
  not1 I800_698(w_800_698, w_014_182);
  nand2 I800_699(w_800_699, w_170_172, w_494_241);
  nand2 I800_700(w_800_700, w_696_115, w_392_083);
  nand2 I800_701(w_800_701, w_113_231, w_541_024);
  not1 I800_702(w_800_702, w_297_054);
  and2 I800_703(w_800_703, w_028_187, w_010_449);
  and2 I800_704(w_800_704, w_788_145, w_132_165);
  nand2 I800_705(w_800_705, w_146_320, w_402_028);
  and2 I800_706(w_800_706, w_096_000, w_091_164);
  and2 I800_707(w_800_707, w_483_428, w_251_013);
  and2 I800_708(w_800_708, w_344_063, w_714_021);
  nand2 I800_709(w_800_709, w_634_264, w_318_015);
  nand2 I800_710(w_800_710, w_222_185, w_368_015);
  not1 I800_711(w_800_711, w_432_053);
  nand2 I800_712(w_800_712, w_386_146, w_547_035);
  not1 I800_713(w_800_713, w_638_380);
  not1 I800_714(w_800_714, w_674_360);
  or2  I800_715(w_800_715, w_023_132, w_057_100);
  not1 I800_716(w_800_716, w_699_231);
  or2  I800_717(w_800_717, w_121_120, w_077_344);

  initial begin
    $get_module_info();
  end
endmodule

// ****** Combined Logic Module Defination ******

// ****** TestBench Module Defination ******

/*
module tb();
  wire  w_000_000, w_000_001, w_000_002, w_000_003, w_000_004, w_000_005, w_000_006, w_000_007, w_000_008, w_000_009, w_000_010, w_000_011, w_000_012, w_000_013, w_000_014, w_000_015, w_000_016, w_000_017, w_000_018, w_000_019, w_000_020, w_000_021, w_000_022, w_000_023, w_000_024, w_000_025, w_000_026, w_000_027, w_000_028, w_000_029, w_000_030, w_000_031, w_000_032, w_000_033, w_000_034, w_000_035, w_000_036, w_000_037, w_000_038, w_000_039, w_000_040, w_000_041, w_000_042, w_000_043, w_000_044, w_000_045, w_000_046, w_000_047, w_000_048, w_000_049, w_000_050, w_000_051, w_000_052, w_000_053, w_000_054, w_000_055, w_000_056, w_000_057, w_000_058, w_000_059, w_000_060, w_000_061, w_000_062, w_000_063, w_000_064, w_000_065, w_000_066, w_000_067, w_000_068, w_000_069, w_000_070, w_000_071, w_000_072, w_000_073, w_000_074, w_000_075, w_000_076, w_000_077, w_000_078, w_000_079, w_000_080, w_000_081, w_000_082, w_000_083, w_000_084, w_000_085, w_000_086, w_000_087, w_000_088, w_000_089, w_000_090, w_000_091, w_000_092, w_000_093, w_000_094, w_000_095, w_000_096, w_000_097, w_000_098, w_000_099, w_000_100, w_000_101, w_000_102, w_000_103, w_000_104, w_000_105, w_000_106, w_000_107, w_000_108, w_000_109, w_000_110, w_000_111, w_000_112, w_000_113, w_000_114, w_000_115, w_000_116, w_000_117, w_000_118, w_000_119, w_000_120, w_000_121, w_000_122, w_000_123, w_000_124, w_000_125, w_000_126, w_000_127, w_000_128, w_000_129, w_000_130, w_000_131, w_000_132, w_000_133, w_000_134, w_000_135, w_000_136, w_000_137, w_000_138, w_000_139, w_000_140, w_000_141, w_000_142, w_000_143, w_000_144, w_000_145, w_000_146, w_000_147, w_000_148, w_000_149, w_000_150, w_000_151, w_000_152, w_000_153, w_000_154, w_000_155, w_000_156, w_000_157, w_000_158, w_000_159, w_000_160, w_000_161, w_000_162, w_000_163, w_000_164, w_000_165, w_000_166, w_000_167, w_000_169, w_000_170, w_000_171, w_000_172, w_000_173, w_000_174, w_000_175, w_000_176, w_000_177, w_000_178, w_000_179, w_000_180, w_000_181, w_000_182, w_000_183, w_000_184, w_000_185, w_000_186, w_000_187, w_000_188, w_000_189, w_000_190, w_000_191, w_000_192, w_000_193, w_000_194, w_000_195, w_000_196, w_000_197, w_000_198, w_000_199, w_000_200, w_000_202, w_000_203, w_000_204, w_000_205, w_000_206, w_000_207, w_000_208, w_000_209, w_000_210, w_000_211, w_000_212, w_000_213, w_000_214, w_000_215, w_000_216, w_000_217, w_000_218, w_000_219, w_000_220, w_000_221, w_000_222, w_000_223, w_000_224, w_000_225, w_000_226, w_000_227, w_000_228, w_000_229, w_000_230, w_000_231, w_000_232, w_000_233, w_000_234, w_000_235, w_000_236, w_000_237, w_000_238, w_000_239, w_000_240, w_000_241, w_000_242, w_000_243, w_000_244, w_000_245, w_000_246, w_000_247, w_000_248, w_000_249, w_000_250, w_000_251, w_000_252, w_000_253, w_000_254, w_000_255, w_000_256, w_000_257, w_000_258, w_000_259, w_000_260, w_000_261, w_000_262, w_000_263, w_000_264, w_000_265, w_000_266, w_000_267, w_000_268, w_000_269, w_000_270, w_000_271, w_000_272, w_000_273, w_000_274, w_000_275, w_000_276, w_000_277, w_000_278, w_000_279, w_000_280, w_000_281, w_000_282, w_000_283, w_000_284, w_000_285, w_000_286, w_000_287, w_000_288, w_000_289, w_000_290, w_000_291, w_000_292, w_000_293, w_000_294, w_000_295, w_000_296, w_000_297, w_000_298, w_000_299, w_000_300, w_000_301, w_000_302, w_000_303, w_000_304, w_000_305, w_000_306, w_000_307, w_000_308, w_000_309, w_000_310, w_000_311, w_000_312, w_000_313, w_000_314, w_000_315, w_000_316, w_000_317, w_000_318, w_000_319, w_000_320, w_000_321, w_000_322, w_000_323, w_000_324, w_000_325, w_000_326, w_000_327, w_000_328, w_000_329, w_000_330, w_000_331, w_000_332, w_000_333, w_000_334, w_000_335, w_000_336, w_000_337, w_000_338, w_000_339, w_000_340, w_000_341, w_000_342, w_000_343, w_000_344, w_000_345, w_000_346, w_000_347, w_000_348, w_000_349, w_000_350, w_000_351, w_000_352, w_000_353, w_000_354, w_000_355, w_000_356, w_000_357, w_000_358, w_000_359, w_000_360, w_000_361, w_000_362, w_000_363, w_000_364, w_000_365, w_000_366, w_000_367, w_000_368, w_000_370, w_000_371, w_000_372, w_000_373, w_000_374, w_000_375, w_000_376, w_000_377, w_000_378, w_000_379, w_000_380, w_000_381, w_000_382, w_000_383, w_000_384, w_000_385, w_000_386, w_000_387, w_000_388, w_000_389, w_000_390, w_000_391, w_000_392, w_000_393, w_000_394, w_000_395, w_000_396, w_000_397, w_000_398, w_000_399, w_000_400, w_000_401, w_000_402, w_000_403, w_000_404, w_000_405, w_000_406, w_000_408, w_000_409, w_000_410, w_000_411, w_000_412, w_000_413, w_000_414, w_000_415, w_000_416, w_000_417, w_000_418, w_000_419, w_000_420, w_000_421, w_000_422, w_000_423, w_000_424, w_000_425, w_000_426, w_000_427, w_000_428, w_000_429, w_000_430, w_000_431, w_000_432, w_000_433, w_000_434, w_000_435, w_000_436, w_000_437, w_000_438, w_000_439, w_000_440, w_000_441, w_000_442, w_000_443, w_000_444, w_000_445, w_000_446, w_000_447, w_000_448, w_000_449, w_000_450, w_000_451, w_000_452, w_000_453, w_000_454, w_000_455, w_000_456, w_000_457, w_000_458, w_000_459, w_000_460, w_000_461, w_000_462, w_000_463, w_000_464, w_000_465, w_000_466, w_000_467, w_000_468, w_000_469, w_000_470, w_000_471, w_000_472, w_000_473, w_000_474, w_000_475, w_000_476, w_000_477, w_000_478, w_000_479, w_000_480, w_000_481, w_000_482, w_000_483, w_000_484, w_000_485, w_000_486, w_000_487, w_000_488, w_000_489, w_000_490, w_000_491, w_000_492, w_000_493, w_000_494, w_000_495, w_000_496, w_000_497, w_000_498, w_000_499, w_000_500, w_000_501, w_000_502, w_000_503, w_000_504, w_000_505, w_000_506, w_000_507, w_000_508, w_000_510, w_000_511, w_000_512, w_000_513, w_000_514, w_000_515, w_000_516, w_000_517, w_000_518, w_000_519, w_000_520, w_000_521, w_000_522, w_000_523, w_000_524, w_000_525, w_000_526, w_000_527, w_000_528, w_000_529, w_000_530, w_000_531, w_000_532, w_000_533, w_000_534, w_000_535, w_000_536, w_000_537, w_000_538, w_000_540, w_000_541, w_000_542, w_000_543, w_000_544, w_000_545, w_000_546, w_000_547, w_000_548, w_000_549, w_000_550, w_000_551, w_000_552, w_000_553, w_000_554, w_000_555, w_000_556, w_000_557, w_000_558, w_000_559, w_000_560, w_000_561, w_000_563, w_000_564, w_000_565, w_000_566, w_000_567, w_000_568, w_000_569, w_000_570, w_000_571, w_000_572, w_000_573, w_000_574, w_000_575, w_000_576, w_000_577, w_000_578, w_000_579, w_000_580, w_000_581, w_000_582, w_000_583, w_000_584, w_000_585, w_000_586, w_000_587, w_000_588, w_000_589, w_000_590, w_000_591, w_000_592, w_000_593, w_000_594, w_000_595, w_000_596, w_000_597, w_000_598, w_000_599, w_000_600, w_000_601, w_000_602, w_000_603, w_000_604, w_000_605, w_000_606, w_000_607, w_000_608, w_000_609, w_000_610, w_000_611, w_000_612, w_000_613, w_000_614, w_000_615, w_000_616, w_000_617, w_000_618, w_000_619, w_000_620, w_000_621, w_000_622, w_000_623, w_000_624, w_000_625, w_000_626, w_000_627, w_000_628, w_000_629, w_000_630, w_000_632, w_000_634, w_000_635, w_000_636, w_000_637, w_000_638, w_000_639, w_000_640, w_000_641, w_000_642, w_000_643, w_000_644, w_000_645, w_000_646, w_000_647, w_000_648, w_000_649, w_000_650, w_000_651, w_000_652, w_000_653, w_000_654, w_000_655, w_000_656, w_000_657, w_000_658, w_000_659, w_000_660, w_000_661, w_000_662, w_000_663, w_000_664, w_000_665, w_000_666, w_000_667, w_000_668, w_000_671, w_000_674, w_000_675, w_000_676, w_000_679, w_000_680, w_000_681, w_000_682, w_000_683, w_000_684, w_000_685, w_000_687, w_000_688, w_000_689, w_000_690, w_000_691, w_000_692, w_000_693, w_000_694, w_000_695, w_000_696, w_000_697, w_000_698, w_000_699, w_000_701, w_000_702, w_000_703, w_000_704, w_000_705, w_000_706, w_000_707, w_000_708, w_000_709, w_000_710, w_000_711, w_000_712, w_000_713, w_000_714, w_000_715, w_000_716, w_000_717, w_000_718, w_000_720, w_000_722, w_000_724, w_000_725, w_000_726, w_000_727, w_000_728, w_000_731, w_000_732, w_000_733, w_000_734, w_000_735, w_000_736, w_000_738, w_000_739, w_000_740, w_000_741, w_000_743, w_000_744, w_000_745, w_000_747, w_000_748, w_000_749, w_000_751, w_000_754, w_000_756, w_000_757, w_000_758, w_000_759, w_000_762, w_000_763, w_000_768, w_000_770, w_000_772, w_000_776, w_000_777, w_000_780, w_000_783, w_800_000, w_800_001, w_800_002, w_800_003, w_800_004, w_800_005, w_800_006, w_800_007, w_800_008, w_800_009, w_800_010, w_800_011, w_800_012, w_800_013, w_800_014, w_800_015, w_800_016, w_800_017, w_800_018, w_800_019, w_800_020, w_800_021, w_800_022, w_800_023, w_800_024, w_800_025, w_800_026, w_800_027, w_800_028, w_800_029, w_800_030, w_800_031, w_800_032, w_800_033, w_800_034, w_800_035, w_800_036, w_800_037, w_800_038, w_800_039, w_800_040, w_800_041, w_800_042, w_800_043, w_800_044, w_800_045, w_800_046, w_800_047, w_800_048, w_800_049, w_800_050, w_800_051, w_800_052, w_800_053, w_800_054, w_800_055, w_800_056, w_800_057, w_800_058, w_800_059, w_800_060, w_800_061, w_800_062, w_800_063, w_800_064, w_800_065, w_800_066, w_800_067, w_800_068, w_800_069, w_800_070, w_800_071, w_800_072, w_800_073, w_800_074, w_800_075, w_800_076, w_800_077, w_800_078, w_800_079, w_800_080, w_800_081, w_800_082, w_800_083, w_800_084, w_800_085, w_800_086, w_800_087, w_800_088, w_800_089, w_800_090, w_800_091, w_800_092, w_800_093, w_800_094, w_800_095, w_800_096, w_800_097, w_800_098, w_800_099, w_800_100, w_800_101, w_800_102, w_800_103, w_800_104, w_800_105, w_800_106, w_800_107, w_800_108, w_800_109, w_800_110, w_800_111, w_800_112, w_800_113, w_800_114, w_800_115, w_800_116, w_800_117, w_800_118, w_800_119, w_800_120, w_800_121, w_800_122, w_800_123, w_800_124, w_800_125, w_800_126, w_800_127, w_800_128, w_800_129, w_800_130, w_800_131, w_800_132, w_800_133, w_800_134, w_800_135, w_800_136, w_800_137, w_800_138, w_800_139, w_800_140, w_800_141, w_800_142, w_800_143, w_800_144, w_800_145, w_800_146, w_800_147, w_800_148, w_800_149, w_800_150, w_800_151, w_800_152, w_800_153, w_800_154, w_800_155, w_800_156, w_800_157, w_800_158, w_800_159, w_800_160, w_800_161, w_800_162, w_800_163, w_800_164, w_800_165, w_800_166, w_800_167, w_800_168, w_800_169, w_800_170, w_800_171, w_800_172, w_800_173, w_800_174, w_800_175, w_800_176, w_800_177, w_800_178, w_800_179, w_800_180, w_800_181, w_800_182, w_800_183, w_800_184, w_800_185, w_800_186, w_800_187, w_800_188, w_800_189, w_800_190, w_800_191, w_800_192, w_800_193, w_800_194, w_800_195, w_800_196, w_800_197, w_800_198, w_800_199, w_800_200, w_800_201, w_800_202, w_800_203, w_800_204, w_800_205, w_800_206, w_800_207, w_800_208, w_800_209, w_800_210, w_800_211, w_800_212, w_800_213, w_800_214, w_800_215, w_800_216, w_800_217, w_800_218, w_800_219, w_800_220, w_800_221, w_800_222, w_800_223, w_800_224, w_800_225, w_800_226, w_800_227, w_800_228, w_800_229, w_800_230, w_800_231, w_800_232, w_800_233, w_800_234, w_800_235, w_800_236, w_800_237, w_800_238, w_800_239, w_800_240, w_800_241, w_800_242, w_800_243, w_800_244, w_800_245, w_800_246, w_800_247, w_800_248, w_800_249, w_800_250, w_800_251, w_800_252, w_800_253, w_800_254, w_800_255, w_800_256, w_800_257, w_800_258, w_800_259, w_800_260, w_800_261, w_800_262, w_800_263, w_800_264, w_800_265, w_800_266, w_800_267, w_800_268, w_800_269, w_800_270, w_800_271, w_800_272, w_800_273, w_800_274, w_800_275, w_800_276, w_800_277, w_800_278, w_800_279, w_800_280, w_800_281, w_800_282, w_800_283, w_800_284, w_800_285, w_800_286, w_800_287, w_800_288, w_800_289, w_800_290, w_800_291, w_800_292, w_800_293, w_800_294, w_800_295, w_800_296, w_800_297, w_800_298, w_800_299, w_800_300, w_800_301, w_800_302, w_800_303, w_800_304, w_800_305, w_800_306, w_800_307, w_800_308, w_800_309, w_800_310, w_800_311, w_800_312, w_800_313, w_800_314, w_800_315, w_800_316, w_800_317, w_800_318, w_800_319, w_800_320, w_800_321, w_800_322, w_800_323, w_800_324, w_800_325, w_800_326, w_800_327, w_800_328, w_800_329, w_800_330, w_800_331, w_800_332, w_800_333, w_800_334, w_800_335, w_800_336, w_800_337, w_800_338, w_800_339, w_800_340, w_800_341, w_800_342, w_800_343, w_800_344, w_800_345, w_800_346, w_800_347, w_800_348, w_800_349, w_800_350, w_800_351, w_800_352, w_800_353, w_800_354, w_800_355, w_800_356, w_800_357, w_800_358, w_800_359, w_800_360, w_800_361, w_800_362, w_800_363, w_800_364, w_800_365, w_800_366, w_800_367, w_800_368, w_800_369, w_800_370, w_800_371, w_800_372, w_800_373, w_800_374, w_800_375, w_800_376, w_800_377, w_800_378, w_800_379, w_800_380, w_800_381, w_800_382, w_800_383, w_800_384, w_800_385, w_800_386, w_800_387, w_800_388, w_800_389, w_800_390, w_800_391, w_800_392, w_800_393, w_800_394, w_800_395, w_800_396, w_800_397, w_800_398, w_800_399, w_800_400, w_800_401, w_800_402, w_800_403, w_800_404, w_800_405, w_800_406, w_800_407, w_800_408, w_800_409, w_800_410, w_800_411, w_800_412, w_800_413, w_800_414, w_800_415, w_800_416, w_800_417, w_800_418, w_800_419, w_800_420, w_800_421, w_800_422, w_800_423, w_800_424, w_800_425, w_800_426, w_800_427, w_800_428, w_800_429, w_800_430, w_800_431, w_800_432, w_800_433, w_800_434, w_800_435, w_800_436, w_800_437, w_800_438, w_800_439, w_800_440, w_800_441, w_800_442, w_800_443, w_800_444, w_800_445, w_800_446, w_800_447, w_800_448, w_800_449, w_800_450, w_800_451, w_800_452, w_800_453, w_800_454, w_800_455, w_800_456, w_800_457, w_800_458, w_800_459, w_800_460, w_800_461, w_800_462, w_800_463, w_800_464, w_800_465, w_800_466, w_800_467, w_800_468, w_800_469, w_800_470, w_800_471, w_800_472, w_800_473, w_800_474, w_800_475, w_800_476, w_800_477, w_800_478, w_800_479, w_800_480, w_800_481, w_800_482, w_800_483, w_800_484, w_800_485, w_800_486, w_800_487, w_800_488, w_800_489, w_800_490, w_800_491, w_800_492, w_800_493, w_800_494, w_800_495, w_800_496, w_800_497, w_800_498, w_800_499, w_800_500, w_800_501, w_800_502, w_800_503, w_800_504, w_800_505, w_800_506, w_800_507, w_800_508, w_800_509, w_800_510, w_800_511, w_800_512, w_800_513, w_800_514, w_800_515, w_800_516, w_800_517, w_800_518, w_800_519, w_800_520, w_800_521, w_800_522, w_800_523, w_800_524, w_800_525, w_800_526, w_800_527, w_800_528, w_800_529, w_800_530, w_800_531, w_800_532, w_800_533, w_800_534, w_800_535, w_800_536, w_800_537, w_800_538, w_800_539, w_800_540, w_800_541, w_800_542, w_800_543, w_800_544, w_800_545, w_800_546, w_800_547, w_800_548, w_800_549, w_800_550, w_800_551, w_800_552, w_800_553, w_800_554, w_800_555, w_800_556, w_800_557, w_800_558, w_800_559, w_800_560, w_800_561, w_800_562, w_800_563, w_800_564, w_800_565, w_800_566, w_800_567, w_800_568, w_800_569, w_800_570, w_800_571, w_800_572, w_800_573, w_800_574, w_800_575, w_800_576, w_800_577, w_800_578, w_800_579, w_800_580, w_800_581, w_800_582, w_800_583, w_800_584, w_800_585, w_800_586, w_800_587, w_800_588, w_800_589, w_800_590, w_800_591, w_800_592, w_800_593, w_800_594, w_800_595, w_800_596, w_800_597, w_800_598, w_800_599, w_800_600, w_800_601, w_800_602, w_800_603, w_800_604, w_800_605, w_800_606, w_800_607, w_800_608, w_800_609, w_800_610, w_800_611, w_800_612, w_800_613, w_800_614, w_800_615, w_800_616, w_800_617, w_800_618, w_800_619, w_800_620, w_800_621, w_800_622, w_800_623, w_800_624, w_800_625, w_800_626, w_800_627, w_800_628, w_800_629, w_800_630, w_800_631, w_800_632, w_800_633, w_800_634, w_800_635, w_800_636, w_800_637, w_800_638, w_800_639, w_800_640, w_800_641, w_800_642, w_800_643, w_800_644, w_800_645, w_800_646, w_800_647, w_800_648, w_800_649, w_800_650, w_800_651, w_800_652, w_800_653, w_800_654, w_800_655, w_800_656, w_800_657, w_800_658, w_800_659, w_800_660, w_800_661, w_800_662, w_800_663, w_800_664, w_800_665, w_800_666, w_800_667, w_800_668, w_800_669, w_800_670, w_800_671, w_800_672, w_800_673, w_800_674, w_800_675, w_800_676, w_800_677, w_800_678, w_800_679, w_800_680, w_800_681, w_800_682, w_800_683, w_800_684, w_800_685, w_800_686, w_800_687, w_800_688, w_800_689, w_800_690, w_800_691, w_800_692, w_800_693, w_800_694, w_800_695, w_800_696, w_800_697, w_800_698, w_800_699, w_800_700, w_800_701, w_800_702, w_800_703, w_800_704, w_800_705, w_800_706, w_800_707, w_800_708, w_800_709, w_800_710, w_800_711, w_800_712, w_800_713, w_800_714, w_800_715, w_800_716, w_800_717 ;
  combLogic I0(  w_000_000, w_000_001, w_000_002, w_000_003, w_000_004, w_000_005, w_000_006, w_000_007, w_000_008, w_000_009, w_000_010, w_000_011, w_000_012, w_000_013, w_000_014, w_000_015, w_000_016, w_000_017, w_000_018, w_000_019, w_000_020, w_000_021, w_000_022, w_000_023, w_000_024, w_000_025, w_000_026, w_000_027, w_000_028, w_000_029, w_000_030, w_000_031, w_000_032, w_000_033, w_000_034, w_000_035, w_000_036, w_000_037, w_000_038, w_000_039, w_000_040, w_000_041, w_000_042, w_000_043, w_000_044, w_000_045, w_000_046, w_000_047, w_000_048, w_000_049, w_000_050, w_000_051, w_000_052, w_000_053, w_000_054, w_000_055, w_000_056, w_000_057, w_000_058, w_000_059, w_000_060, w_000_061, w_000_062, w_000_063, w_000_064, w_000_065, w_000_066, w_000_067, w_000_068, w_000_069, w_000_070, w_000_071, w_000_072, w_000_073, w_000_074, w_000_075, w_000_076, w_000_077, w_000_078, w_000_079, w_000_080, w_000_081, w_000_082, w_000_083, w_000_084, w_000_085, w_000_086, w_000_087, w_000_088, w_000_089, w_000_090, w_000_091, w_000_092, w_000_093, w_000_094, w_000_095, w_000_096, w_000_097, w_000_098, w_000_099, w_000_100, w_000_101, w_000_102, w_000_103, w_000_104, w_000_105, w_000_106, w_000_107, w_000_108, w_000_109, w_000_110, w_000_111, w_000_112, w_000_113, w_000_114, w_000_115, w_000_116, w_000_117, w_000_118, w_000_119, w_000_120, w_000_121, w_000_122, w_000_123, w_000_124, w_000_125, w_000_126, w_000_127, w_000_128, w_000_129, w_000_130, w_000_131, w_000_132, w_000_133, w_000_134, w_000_135, w_000_136, w_000_137, w_000_138, w_000_139, w_000_140, w_000_141, w_000_142, w_000_143, w_000_144, w_000_145, w_000_146, w_000_147, w_000_148, w_000_149, w_000_150, w_000_151, w_000_152, w_000_153, w_000_154, w_000_155, w_000_156, w_000_157, w_000_158, w_000_159, w_000_160, w_000_161, w_000_162, w_000_163, w_000_164, w_000_165, w_000_166, w_000_167, w_000_169, w_000_170, w_000_171, w_000_172, w_000_173, w_000_174, w_000_175, w_000_176, w_000_177, w_000_178, w_000_179, w_000_180, w_000_181, w_000_182, w_000_183, w_000_184, w_000_185, w_000_186, w_000_187, w_000_188, w_000_189, w_000_190, w_000_191, w_000_192, w_000_193, w_000_194, w_000_195, w_000_196, w_000_197, w_000_198, w_000_199, w_000_200, w_000_202, w_000_203, w_000_204, w_000_205, w_000_206, w_000_207, w_000_208, w_000_209, w_000_210, w_000_211, w_000_212, w_000_213, w_000_214, w_000_215, w_000_216, w_000_217, w_000_218, w_000_219, w_000_220, w_000_221, w_000_222, w_000_223, w_000_224, w_000_225, w_000_226, w_000_227, w_000_228, w_000_229, w_000_230, w_000_231, w_000_232, w_000_233, w_000_234, w_000_235, w_000_236, w_000_237, w_000_238, w_000_239, w_000_240, w_000_241, w_000_242, w_000_243, w_000_244, w_000_245, w_000_246, w_000_247, w_000_248, w_000_249, w_000_250, w_000_251, w_000_252, w_000_253, w_000_254, w_000_255, w_000_256, w_000_257, w_000_258, w_000_259, w_000_260, w_000_261, w_000_262, w_000_263, w_000_264, w_000_265, w_000_266, w_000_267, w_000_268, w_000_269, w_000_270, w_000_271, w_000_272, w_000_273, w_000_274, w_000_275, w_000_276, w_000_277, w_000_278, w_000_279, w_000_280, w_000_281, w_000_282, w_000_283, w_000_284, w_000_285, w_000_286, w_000_287, w_000_288, w_000_289, w_000_290, w_000_291, w_000_292, w_000_293, w_000_294, w_000_295, w_000_296, w_000_297, w_000_298, w_000_299, w_000_300, w_000_301, w_000_302, w_000_303, w_000_304, w_000_305, w_000_306, w_000_307, w_000_308, w_000_309, w_000_310, w_000_311, w_000_312, w_000_313, w_000_314, w_000_315, w_000_316, w_000_317, w_000_318, w_000_319, w_000_320, w_000_321, w_000_322, w_000_323, w_000_324, w_000_325, w_000_326, w_000_327, w_000_328, w_000_329, w_000_330, w_000_331, w_000_332, w_000_333, w_000_334, w_000_335, w_000_336, w_000_337, w_000_338, w_000_339, w_000_340, w_000_341, w_000_342, w_000_343, w_000_344, w_000_345, w_000_346, w_000_347, w_000_348, w_000_349, w_000_350, w_000_351, w_000_352, w_000_353, w_000_354, w_000_355, w_000_356, w_000_357, w_000_358, w_000_359, w_000_360, w_000_361, w_000_362, w_000_363, w_000_364, w_000_365, w_000_366, w_000_367, w_000_368, w_000_370, w_000_371, w_000_372, w_000_373, w_000_374, w_000_375, w_000_376, w_000_377, w_000_378, w_000_379, w_000_380, w_000_381, w_000_382, w_000_383, w_000_384, w_000_385, w_000_386, w_000_387, w_000_388, w_000_389, w_000_390, w_000_391, w_000_392, w_000_393, w_000_394, w_000_395, w_000_396, w_000_397, w_000_398, w_000_399, w_000_400, w_000_401, w_000_402, w_000_403, w_000_404, w_000_405, w_000_406, w_000_408, w_000_409, w_000_410, w_000_411, w_000_412, w_000_413, w_000_414, w_000_415, w_000_416, w_000_417, w_000_418, w_000_419, w_000_420, w_000_421, w_000_422, w_000_423, w_000_424, w_000_425, w_000_426, w_000_427, w_000_428, w_000_429, w_000_430, w_000_431, w_000_432, w_000_433, w_000_434, w_000_435, w_000_436, w_000_437, w_000_438, w_000_439, w_000_440, w_000_441, w_000_442, w_000_443, w_000_444, w_000_445, w_000_446, w_000_447, w_000_448, w_000_449, w_000_450, w_000_451, w_000_452, w_000_453, w_000_454, w_000_455, w_000_456, w_000_457, w_000_458, w_000_459, w_000_460, w_000_461, w_000_462, w_000_463, w_000_464, w_000_465, w_000_466, w_000_467, w_000_468, w_000_469, w_000_470, w_000_471, w_000_472, w_000_473, w_000_474, w_000_475, w_000_476, w_000_477, w_000_478, w_000_479, w_000_480, w_000_481, w_000_482, w_000_483, w_000_484, w_000_485, w_000_486, w_000_487, w_000_488, w_000_489, w_000_490, w_000_491, w_000_492, w_000_493, w_000_494, w_000_495, w_000_496, w_000_497, w_000_498, w_000_499, w_000_500, w_000_501, w_000_502, w_000_503, w_000_504, w_000_505, w_000_506, w_000_507, w_000_508, w_000_510, w_000_511, w_000_512, w_000_513, w_000_514, w_000_515, w_000_516, w_000_517, w_000_518, w_000_519, w_000_520, w_000_521, w_000_522, w_000_523, w_000_524, w_000_525, w_000_526, w_000_527, w_000_528, w_000_529, w_000_530, w_000_531, w_000_532, w_000_533, w_000_534, w_000_535, w_000_536, w_000_537, w_000_538, w_000_540, w_000_541, w_000_542, w_000_543, w_000_544, w_000_545, w_000_546, w_000_547, w_000_548, w_000_549, w_000_550, w_000_551, w_000_552, w_000_553, w_000_554, w_000_555, w_000_556, w_000_557, w_000_558, w_000_559, w_000_560, w_000_561, w_000_563, w_000_564, w_000_565, w_000_566, w_000_567, w_000_568, w_000_569, w_000_570, w_000_571, w_000_572, w_000_573, w_000_574, w_000_575, w_000_576, w_000_577, w_000_578, w_000_579, w_000_580, w_000_581, w_000_582, w_000_583, w_000_584, w_000_585, w_000_586, w_000_587, w_000_588, w_000_589, w_000_590, w_000_591, w_000_592, w_000_593, w_000_594, w_000_595, w_000_596, w_000_597, w_000_598, w_000_599, w_000_600, w_000_601, w_000_602, w_000_603, w_000_604, w_000_605, w_000_606, w_000_607, w_000_608, w_000_609, w_000_610, w_000_611, w_000_612, w_000_613, w_000_614, w_000_615, w_000_616, w_000_617, w_000_618, w_000_619, w_000_620, w_000_621, w_000_622, w_000_623, w_000_624, w_000_625, w_000_626, w_000_627, w_000_628, w_000_629, w_000_630, w_000_632, w_000_634, w_000_635, w_000_636, w_000_637, w_000_638, w_000_639, w_000_640, w_000_641, w_000_642, w_000_643, w_000_644, w_000_645, w_000_646, w_000_647, w_000_648, w_000_649, w_000_650, w_000_651, w_000_652, w_000_653, w_000_654, w_000_655, w_000_656, w_000_657, w_000_658, w_000_659, w_000_660, w_000_661, w_000_662, w_000_663, w_000_664, w_000_665, w_000_666, w_000_667, w_000_668, w_000_671, w_000_674, w_000_675, w_000_676, w_000_679, w_000_680, w_000_681, w_000_682, w_000_683, w_000_684, w_000_685, w_000_687, w_000_688, w_000_689, w_000_690, w_000_691, w_000_692, w_000_693, w_000_694, w_000_695, w_000_696, w_000_697, w_000_698, w_000_699, w_000_701, w_000_702, w_000_703, w_000_704, w_000_705, w_000_706, w_000_707, w_000_708, w_000_709, w_000_710, w_000_711, w_000_712, w_000_713, w_000_714, w_000_715, w_000_716, w_000_717, w_000_718, w_000_720, w_000_722, w_000_724, w_000_725, w_000_726, w_000_727, w_000_728, w_000_731, w_000_732, w_000_733, w_000_734, w_000_735, w_000_736, w_000_738, w_000_739, w_000_740, w_000_741, w_000_743, w_000_744, w_000_745, w_000_747, w_000_748, w_000_749, w_000_751, w_000_754, w_000_756, w_000_757, w_000_758, w_000_759, w_000_762, w_000_763, w_000_768, w_000_770, w_000_772, w_000_776, w_000_777, w_000_780, w_000_783, w_800_000, w_800_001, w_800_002, w_800_003, w_800_004, w_800_005, w_800_006, w_800_007, w_800_008, w_800_009, w_800_010, w_800_011, w_800_012, w_800_013, w_800_014, w_800_015, w_800_016, w_800_017, w_800_018, w_800_019, w_800_020, w_800_021, w_800_022, w_800_023, w_800_024, w_800_025, w_800_026, w_800_027, w_800_028, w_800_029, w_800_030, w_800_031, w_800_032, w_800_033, w_800_034, w_800_035, w_800_036, w_800_037, w_800_038, w_800_039, w_800_040, w_800_041, w_800_042, w_800_043, w_800_044, w_800_045, w_800_046, w_800_047, w_800_048, w_800_049, w_800_050, w_800_051, w_800_052, w_800_053, w_800_054, w_800_055, w_800_056, w_800_057, w_800_058, w_800_059, w_800_060, w_800_061, w_800_062, w_800_063, w_800_064, w_800_065, w_800_066, w_800_067, w_800_068, w_800_069, w_800_070, w_800_071, w_800_072, w_800_073, w_800_074, w_800_075, w_800_076, w_800_077, w_800_078, w_800_079, w_800_080, w_800_081, w_800_082, w_800_083, w_800_084, w_800_085, w_800_086, w_800_087, w_800_088, w_800_089, w_800_090, w_800_091, w_800_092, w_800_093, w_800_094, w_800_095, w_800_096, w_800_097, w_800_098, w_800_099, w_800_100, w_800_101, w_800_102, w_800_103, w_800_104, w_800_105, w_800_106, w_800_107, w_800_108, w_800_109, w_800_110, w_800_111, w_800_112, w_800_113, w_800_114, w_800_115, w_800_116, w_800_117, w_800_118, w_800_119, w_800_120, w_800_121, w_800_122, w_800_123, w_800_124, w_800_125, w_800_126, w_800_127, w_800_128, w_800_129, w_800_130, w_800_131, w_800_132, w_800_133, w_800_134, w_800_135, w_800_136, w_800_137, w_800_138, w_800_139, w_800_140, w_800_141, w_800_142, w_800_143, w_800_144, w_800_145, w_800_146, w_800_147, w_800_148, w_800_149, w_800_150, w_800_151, w_800_152, w_800_153, w_800_154, w_800_155, w_800_156, w_800_157, w_800_158, w_800_159, w_800_160, w_800_161, w_800_162, w_800_163, w_800_164, w_800_165, w_800_166, w_800_167, w_800_168, w_800_169, w_800_170, w_800_171, w_800_172, w_800_173, w_800_174, w_800_175, w_800_176, w_800_177, w_800_178, w_800_179, w_800_180, w_800_181, w_800_182, w_800_183, w_800_184, w_800_185, w_800_186, w_800_187, w_800_188, w_800_189, w_800_190, w_800_191, w_800_192, w_800_193, w_800_194, w_800_195, w_800_196, w_800_197, w_800_198, w_800_199, w_800_200, w_800_201, w_800_202, w_800_203, w_800_204, w_800_205, w_800_206, w_800_207, w_800_208, w_800_209, w_800_210, w_800_211, w_800_212, w_800_213, w_800_214, w_800_215, w_800_216, w_800_217, w_800_218, w_800_219, w_800_220, w_800_221, w_800_222, w_800_223, w_800_224, w_800_225, w_800_226, w_800_227, w_800_228, w_800_229, w_800_230, w_800_231, w_800_232, w_800_233, w_800_234, w_800_235, w_800_236, w_800_237, w_800_238, w_800_239, w_800_240, w_800_241, w_800_242, w_800_243, w_800_244, w_800_245, w_800_246, w_800_247, w_800_248, w_800_249, w_800_250, w_800_251, w_800_252, w_800_253, w_800_254, w_800_255, w_800_256, w_800_257, w_800_258, w_800_259, w_800_260, w_800_261, w_800_262, w_800_263, w_800_264, w_800_265, w_800_266, w_800_267, w_800_268, w_800_269, w_800_270, w_800_271, w_800_272, w_800_273, w_800_274, w_800_275, w_800_276, w_800_277, w_800_278, w_800_279, w_800_280, w_800_281, w_800_282, w_800_283, w_800_284, w_800_285, w_800_286, w_800_287, w_800_288, w_800_289, w_800_290, w_800_291, w_800_292, w_800_293, w_800_294, w_800_295, w_800_296, w_800_297, w_800_298, w_800_299, w_800_300, w_800_301, w_800_302, w_800_303, w_800_304, w_800_305, w_800_306, w_800_307, w_800_308, w_800_309, w_800_310, w_800_311, w_800_312, w_800_313, w_800_314, w_800_315, w_800_316, w_800_317, w_800_318, w_800_319, w_800_320, w_800_321, w_800_322, w_800_323, w_800_324, w_800_325, w_800_326, w_800_327, w_800_328, w_800_329, w_800_330, w_800_331, w_800_332, w_800_333, w_800_334, w_800_335, w_800_336, w_800_337, w_800_338, w_800_339, w_800_340, w_800_341, w_800_342, w_800_343, w_800_344, w_800_345, w_800_346, w_800_347, w_800_348, w_800_349, w_800_350, w_800_351, w_800_352, w_800_353, w_800_354, w_800_355, w_800_356, w_800_357, w_800_358, w_800_359, w_800_360, w_800_361, w_800_362, w_800_363, w_800_364, w_800_365, w_800_366, w_800_367, w_800_368, w_800_369, w_800_370, w_800_371, w_800_372, w_800_373, w_800_374, w_800_375, w_800_376, w_800_377, w_800_378, w_800_379, w_800_380, w_800_381, w_800_382, w_800_383, w_800_384, w_800_385, w_800_386, w_800_387, w_800_388, w_800_389, w_800_390, w_800_391, w_800_392, w_800_393, w_800_394, w_800_395, w_800_396, w_800_397, w_800_398, w_800_399, w_800_400, w_800_401, w_800_402, w_800_403, w_800_404, w_800_405, w_800_406, w_800_407, w_800_408, w_800_409, w_800_410, w_800_411, w_800_412, w_800_413, w_800_414, w_800_415, w_800_416, w_800_417, w_800_418, w_800_419, w_800_420, w_800_421, w_800_422, w_800_423, w_800_424, w_800_425, w_800_426, w_800_427, w_800_428, w_800_429, w_800_430, w_800_431, w_800_432, w_800_433, w_800_434, w_800_435, w_800_436, w_800_437, w_800_438, w_800_439, w_800_440, w_800_441, w_800_442, w_800_443, w_800_444, w_800_445, w_800_446, w_800_447, w_800_448, w_800_449, w_800_450, w_800_451, w_800_452, w_800_453, w_800_454, w_800_455, w_800_456, w_800_457, w_800_458, w_800_459, w_800_460, w_800_461, w_800_462, w_800_463, w_800_464, w_800_465, w_800_466, w_800_467, w_800_468, w_800_469, w_800_470, w_800_471, w_800_472, w_800_473, w_800_474, w_800_475, w_800_476, w_800_477, w_800_478, w_800_479, w_800_480, w_800_481, w_800_482, w_800_483, w_800_484, w_800_485, w_800_486, w_800_487, w_800_488, w_800_489, w_800_490, w_800_491, w_800_492, w_800_493, w_800_494, w_800_495, w_800_496, w_800_497, w_800_498, w_800_499, w_800_500, w_800_501, w_800_502, w_800_503, w_800_504, w_800_505, w_800_506, w_800_507, w_800_508, w_800_509, w_800_510, w_800_511, w_800_512, w_800_513, w_800_514, w_800_515, w_800_516, w_800_517, w_800_518, w_800_519, w_800_520, w_800_521, w_800_522, w_800_523, w_800_524, w_800_525, w_800_526, w_800_527, w_800_528, w_800_529, w_800_530, w_800_531, w_800_532, w_800_533, w_800_534, w_800_535, w_800_536, w_800_537, w_800_538, w_800_539, w_800_540, w_800_541, w_800_542, w_800_543, w_800_544, w_800_545, w_800_546, w_800_547, w_800_548, w_800_549, w_800_550, w_800_551, w_800_552, w_800_553, w_800_554, w_800_555, w_800_556, w_800_557, w_800_558, w_800_559, w_800_560, w_800_561, w_800_562, w_800_563, w_800_564, w_800_565, w_800_566, w_800_567, w_800_568, w_800_569, w_800_570, w_800_571, w_800_572, w_800_573, w_800_574, w_800_575, w_800_576, w_800_577, w_800_578, w_800_579, w_800_580, w_800_581, w_800_582, w_800_583, w_800_584, w_800_585, w_800_586, w_800_587, w_800_588, w_800_589, w_800_590, w_800_591, w_800_592, w_800_593, w_800_594, w_800_595, w_800_596, w_800_597, w_800_598, w_800_599, w_800_600, w_800_601, w_800_602, w_800_603, w_800_604, w_800_605, w_800_606, w_800_607, w_800_608, w_800_609, w_800_610, w_800_611, w_800_612, w_800_613, w_800_614, w_800_615, w_800_616, w_800_617, w_800_618, w_800_619, w_800_620, w_800_621, w_800_622, w_800_623, w_800_624, w_800_625, w_800_626, w_800_627, w_800_628, w_800_629, w_800_630, w_800_631, w_800_632, w_800_633, w_800_634, w_800_635, w_800_636, w_800_637, w_800_638, w_800_639, w_800_640, w_800_641, w_800_642, w_800_643, w_800_644, w_800_645, w_800_646, w_800_647, w_800_648, w_800_649, w_800_650, w_800_651, w_800_652, w_800_653, w_800_654, w_800_655, w_800_656, w_800_657, w_800_658, w_800_659, w_800_660, w_800_661, w_800_662, w_800_663, w_800_664, w_800_665, w_800_666, w_800_667, w_800_668, w_800_669, w_800_670, w_800_671, w_800_672, w_800_673, w_800_674, w_800_675, w_800_676, w_800_677, w_800_678, w_800_679, w_800_680, w_800_681, w_800_682, w_800_683, w_800_684, w_800_685, w_800_686, w_800_687, w_800_688, w_800_689, w_800_690, w_800_691, w_800_692, w_800_693, w_800_694, w_800_695, w_800_696, w_800_697, w_800_698, w_800_699, w_800_700, w_800_701, w_800_702, w_800_703, w_800_704, w_800_705, w_800_706, w_800_707, w_800_708, w_800_709, w_800_710, w_800_711, w_800_712, w_800_713, w_800_714, w_800_715, w_800_716, w_800_717  );

  reg r0, r1, r2, r3, r4, r5, r6, r7, r8, r9, r10, r11, r12, r13, r14, r15, r16, r17, r18, r19, r20, r21, r22, r23, r24, r25, r26, r27, r28, r29, r30, r31, r32, r33, r34, r35, r36, r37, r38, r39, r40, r41, r42, r43, r44, r45, r46, r47, r48, r49, r50, r51, r52, r53, r54, r55, r56, r57, r58, r59, r60, r61, r62, r63, r64, r65, r66, r67, r68, r69, r70, r71, r72, r73, r74, r75, r76, r77, r78, r79, r80, r81, r82, r83, r84, r85, r86, r87, r88, r89, r90, r91, r92, r93, r94, r95, r96, r97, r98, r99, r100, r101, r102, r103, r104, r105, r106, r107, r108, r109, r110, r111, r112, r113, r114, r115, r116, r117, r118, r119, r120, r121, r122, r123, r124, r125, r126, r127, r128, r129, r130, r131, r132, r133, r134, r135, r136, r137, r138, r139, r140, r141, r142, r143, r144, r145, r146, r147, r148, r149, r150, r151, r152, r153, r154, r155, r156, r157, r158, r159, r160, r161, r162, r163, r164, r165, r166, r167, r168, r169, r170, r171, r172, r173, r174, r175, r176, r177, r178, r179, r180, r181, r182, r183, r184, r185, r186, r187, r188, r189, r190, r191, r192, r193, r194, r195, r196, r197, r198, r199, r200, r201, r202, r203, r204, r205, r206, r207, r208, r209, r210, r211, r212, r213, r214, r215, r216, r217, r218, r219, r220, r221, r222, r223, r224, r225, r226, r227, r228, r229, r230, r231, r232, r233, r234, r235, r236, r237, r238, r239, r240, r241, r242, r243, r244, r245, r246, r247, r248, r249, r250, r251, r252, r253, r254, r255, r256, r257, r258, r259, r260, r261, r262, r263, r264, r265, r266, r267, r268, r269, r270, r271, r272, r273, r274, r275, r276, r277, r278, r279, r280, r281, r282, r283, r284, r285, r286, r287, r288, r289, r290, r291, r292, r293, r294, r295, r296, r297, r298, r299, r300, r301, r302, r303, r304, r305, r306, r307, r308, r309, r310, r311, r312, r313, r314, r315, r316, r317, r318, r319, r320, r321, r322, r323, r324, r325, r326, r327, r328, r329, r330, r331, r332, r333, r334, r335, r336, r337, r338, r339, r340, r341, r342, r343, r344, r345, r346, r347, r348, r349, r350, r351, r352, r353, r354, r355, r356, r357, r358, r359, r360, r361, r362, r363, r364, r365, r366, r367, r368, r369, r370, r371, r372, r373, r374, r375, r376, r377, r378, r379, r380, r381, r382, r383, r384, r385, r386, r387, r388, r389, r390, r391, r392, r393, r394, r395, r396, r397, r398, r399, r400, r401, r402, r403, r404, r405, r406, r407, r408, r409, r410, r411, r412, r413, r414, r415, r416, r417, r418, r419, r420, r421, r422, r423, r424, r425, r426, r427, r428, r429, r430, r431, r432, r433, r434, r435, r436, r437, r438, r439, r440, r441, r442, r443, r444, r445, r446, r447, r448, r449, r450, r451, r452, r453, r454, r455, r456, r457, r458, r459, r460, r461, r462, r463, r464, r465, r466, r467, r468, r469, r470, r471, r472, r473, r474, r475, r476, r477, r478, r479, r480, r481, r482, r483, r484, r485, r486, r487, r488, r489, r490, r491, r492, r493, r494, r495, r496, r497, r498, r499, r500, r501, r502, r503, r504, r505, r506, r507, r508, r509, r510, r511, r512, r513, r514, r515, r516, r517, r518, r519, r520, r521, r522, r523, r524, r525, r526, r527, r528, r529, r530, r531, r532, r533, r534, r535, r536, r537, r538, r539, r540, r541, r542, r543, r544, r545, r546, r547, r548, r549, r550, r551, r552, r553, r554, r555, r556, r557, r558, r559, r560, r561, r562, r563, r564, r565, r566, r567, r568, r569, r570, r571, r572, r573, r574, r575, r576, r577, r578, r579, r580, r581, r582, r583, r584, r585, r586, r587, r588, r589, r590, r591, r592, r593, r594, r595, r596, r597, r598, r599, r600, r601, r602, r603, r604, r605, r606, r607, r608, r609, r610, r611, r612, r613, r614, r615, r616, r617, r618, r619, r620, r621, r622, r623, r624, r625, r626, r627, r628, r629, r630, r631, r632, r633, r634, r635, r636, r637, r638, r639, r640, r641, r642, r643, r644, r645, r646, r647, r648, r649, r650, r651, r652, r653, r654, r655, r656, r657, r658, r659, r660, r661, r662, r663, r664, r665, r666, r667, r668, r669, r670, r671, r672, r673, r674, r675, r676, r677, r678, r679, r680, r681, r682, r683, r684, r685, r686, r687, r688, r689, r690, r691, r692, r693, r694, r695, r696, r697, r698, r699, r700, r701, r702, r703, r704, r705, r706, r707, r708, r709, r710, r711, r712, r713, r714, r715, r716, r717, r718, r719, r720, r721, r722, r723, r724, r725, r726, r727, r728, r729, r730, r731, r732, r733, r734, r735, r736, r737, r738, r739, r740, r741, r742, r743, r744, r745, r746, r747, r748, r749, r750, r751, r752, r753, r754, r755, r756, r757, r758, r759, r760, r761, r762, r763, r764, r765, r766, r767, r768, r769, r770, r771, r772, r773, r774, r775, r776, r777, r778, r779, r780, r781, r782, r783, r784, r785, r786, r787, r788, r789, r790, r791, r792, r793, r794, r795, r796, r797, rEnd; 

  assign w_000_000 = r0;
  assign w_000_001 = r1;
  assign w_000_002 = r2;
  assign w_000_003 = r3;
  assign w_000_004 = r4;
  assign w_000_005 = r5;
  assign w_000_006 = r6;
  assign w_000_007 = r7;
  assign w_000_008 = r8;
  assign w_000_009 = r9;
  assign w_000_010 = r10;
  assign w_000_011 = r11;
  assign w_000_012 = r12;
  assign w_000_013 = r13;
  assign w_000_014 = r14;
  assign w_000_015 = r15;
  assign w_000_016 = r16;
  assign w_000_017 = r17;
  assign w_000_018 = r18;
  assign w_000_019 = r19;
  assign w_000_020 = r20;
  assign w_000_021 = r21;
  assign w_000_022 = r22;
  assign w_000_023 = r23;
  assign w_000_024 = r24;
  assign w_000_025 = r25;
  assign w_000_026 = r26;
  assign w_000_027 = r27;
  assign w_000_028 = r28;
  assign w_000_029 = r29;
  assign w_000_030 = r30;
  assign w_000_031 = r31;
  assign w_000_032 = r32;
  assign w_000_033 = r33;
  assign w_000_034 = r34;
  assign w_000_035 = r35;
  assign w_000_036 = r36;
  assign w_000_037 = r37;
  assign w_000_038 = r38;
  assign w_000_039 = r39;
  assign w_000_040 = r40;
  assign w_000_041 = r41;
  assign w_000_042 = r42;
  assign w_000_043 = r43;
  assign w_000_044 = r44;
  assign w_000_045 = r45;
  assign w_000_046 = r46;
  assign w_000_047 = r47;
  assign w_000_048 = r48;
  assign w_000_049 = r49;
  assign w_000_050 = r50;
  assign w_000_051 = r51;
  assign w_000_052 = r52;
  assign w_000_053 = r53;
  assign w_000_054 = r54;
  assign w_000_055 = r55;
  assign w_000_056 = r56;
  assign w_000_057 = r57;
  assign w_000_058 = r58;
  assign w_000_059 = r59;
  assign w_000_060 = r60;
  assign w_000_061 = r61;
  assign w_000_062 = r62;
  assign w_000_063 = r63;
  assign w_000_064 = r64;
  assign w_000_065 = r65;
  assign w_000_066 = r66;
  assign w_000_067 = r67;
  assign w_000_068 = r68;
  assign w_000_069 = r69;
  assign w_000_070 = r70;
  assign w_000_071 = r71;
  assign w_000_072 = r72;
  assign w_000_073 = r73;
  assign w_000_074 = r74;
  assign w_000_075 = r75;
  assign w_000_076 = r76;
  assign w_000_077 = r77;
  assign w_000_078 = r78;
  assign w_000_079 = r79;
  assign w_000_080 = r80;
  assign w_000_081 = r81;
  assign w_000_082 = r82;
  assign w_000_083 = r83;
  assign w_000_084 = r84;
  assign w_000_085 = r85;
  assign w_000_086 = r86;
  assign w_000_087 = r87;
  assign w_000_088 = r88;
  assign w_000_089 = r89;
  assign w_000_090 = r90;
  assign w_000_091 = r91;
  assign w_000_092 = r92;
  assign w_000_093 = r93;
  assign w_000_094 = r94;
  assign w_000_095 = r95;
  assign w_000_096 = r96;
  assign w_000_097 = r97;
  assign w_000_098 = r98;
  assign w_000_099 = r99;
  assign w_000_100 = r100;
  assign w_000_101 = r101;
  assign w_000_102 = r102;
  assign w_000_103 = r103;
  assign w_000_104 = r104;
  assign w_000_105 = r105;
  assign w_000_106 = r106;
  assign w_000_107 = r107;
  assign w_000_108 = r108;
  assign w_000_109 = r109;
  assign w_000_110 = r110;
  assign w_000_111 = r111;
  assign w_000_112 = r112;
  assign w_000_113 = r113;
  assign w_000_114 = r114;
  assign w_000_115 = r115;
  assign w_000_116 = r116;
  assign w_000_117 = r117;
  assign w_000_118 = r118;
  assign w_000_119 = r119;
  assign w_000_120 = r120;
  assign w_000_121 = r121;
  assign w_000_122 = r122;
  assign w_000_123 = r123;
  assign w_000_124 = r124;
  assign w_000_125 = r125;
  assign w_000_126 = r126;
  assign w_000_127 = r127;
  assign w_000_128 = r128;
  assign w_000_129 = r129;
  assign w_000_130 = r130;
  assign w_000_131 = r131;
  assign w_000_132 = r132;
  assign w_000_133 = r133;
  assign w_000_134 = r134;
  assign w_000_135 = r135;
  assign w_000_136 = r136;
  assign w_000_137 = r137;
  assign w_000_138 = r138;
  assign w_000_139 = r139;
  assign w_000_140 = r140;
  assign w_000_141 = r141;
  assign w_000_142 = r142;
  assign w_000_143 = r143;
  assign w_000_144 = r144;
  assign w_000_145 = r145;
  assign w_000_146 = r146;
  assign w_000_147 = r147;
  assign w_000_148 = r148;
  assign w_000_149 = r149;
  assign w_000_150 = r150;
  assign w_000_151 = r151;
  assign w_000_152 = r152;
  assign w_000_153 = r153;
  assign w_000_154 = r154;
  assign w_000_155 = r155;
  assign w_000_156 = r156;
  assign w_000_157 = r157;
  assign w_000_158 = r158;
  assign w_000_159 = r159;
  assign w_000_160 = r160;
  assign w_000_161 = r161;
  assign w_000_162 = r162;
  assign w_000_163 = r163;
  assign w_000_164 = r164;
  assign w_000_165 = r165;
  assign w_000_166 = r166;
  assign w_000_167 = r167;
  assign w_000_168 = r168;
  assign w_000_169 = r169;
  assign w_000_170 = r170;
  assign w_000_171 = r171;
  assign w_000_172 = r172;
  assign w_000_173 = r173;
  assign w_000_174 = r174;
  assign w_000_175 = r175;
  assign w_000_176 = r176;
  assign w_000_177 = r177;
  assign w_000_178 = r178;
  assign w_000_179 = r179;
  assign w_000_180 = r180;
  assign w_000_181 = r181;
  assign w_000_182 = r182;
  assign w_000_183 = r183;
  assign w_000_184 = r184;
  assign w_000_185 = r185;
  assign w_000_186 = r186;
  assign w_000_187 = r187;
  assign w_000_188 = r188;
  assign w_000_189 = r189;
  assign w_000_190 = r190;
  assign w_000_191 = r191;
  assign w_000_192 = r192;
  assign w_000_193 = r193;
  assign w_000_194 = r194;
  assign w_000_195 = r195;
  assign w_000_196 = r196;
  assign w_000_197 = r197;
  assign w_000_198 = r198;
  assign w_000_199 = r199;
  assign w_000_200 = r200;
  assign w_000_201 = r201;
  assign w_000_202 = r202;
  assign w_000_203 = r203;
  assign w_000_204 = r204;
  assign w_000_205 = r205;
  assign w_000_206 = r206;
  assign w_000_207 = r207;
  assign w_000_208 = r208;
  assign w_000_209 = r209;
  assign w_000_210 = r210;
  assign w_000_211 = r211;
  assign w_000_212 = r212;
  assign w_000_213 = r213;
  assign w_000_214 = r214;
  assign w_000_215 = r215;
  assign w_000_216 = r216;
  assign w_000_217 = r217;
  assign w_000_218 = r218;
  assign w_000_219 = r219;
  assign w_000_220 = r220;
  assign w_000_221 = r221;
  assign w_000_222 = r222;
  assign w_000_223 = r223;
  assign w_000_224 = r224;
  assign w_000_225 = r225;
  assign w_000_226 = r226;
  assign w_000_227 = r227;
  assign w_000_228 = r228;
  assign w_000_229 = r229;
  assign w_000_230 = r230;
  assign w_000_231 = r231;
  assign w_000_232 = r232;
  assign w_000_233 = r233;
  assign w_000_234 = r234;
  assign w_000_235 = r235;
  assign w_000_236 = r236;
  assign w_000_237 = r237;
  assign w_000_238 = r238;
  assign w_000_239 = r239;
  assign w_000_240 = r240;
  assign w_000_241 = r241;
  assign w_000_242 = r242;
  assign w_000_243 = r243;
  assign w_000_244 = r244;
  assign w_000_245 = r245;
  assign w_000_246 = r246;
  assign w_000_247 = r247;
  assign w_000_248 = r248;
  assign w_000_249 = r249;
  assign w_000_250 = r250;
  assign w_000_251 = r251;
  assign w_000_252 = r252;
  assign w_000_253 = r253;
  assign w_000_254 = r254;
  assign w_000_255 = r255;
  assign w_000_256 = r256;
  assign w_000_257 = r257;
  assign w_000_258 = r258;
  assign w_000_259 = r259;
  assign w_000_260 = r260;
  assign w_000_261 = r261;
  assign w_000_262 = r262;
  assign w_000_263 = r263;
  assign w_000_264 = r264;
  assign w_000_265 = r265;
  assign w_000_266 = r266;
  assign w_000_267 = r267;
  assign w_000_268 = r268;
  assign w_000_269 = r269;
  assign w_000_270 = r270;
  assign w_000_271 = r271;
  assign w_000_272 = r272;
  assign w_000_273 = r273;
  assign w_000_274 = r274;
  assign w_000_275 = r275;
  assign w_000_276 = r276;
  assign w_000_277 = r277;
  assign w_000_278 = r278;
  assign w_000_279 = r279;
  assign w_000_280 = r280;
  assign w_000_281 = r281;
  assign w_000_282 = r282;
  assign w_000_283 = r283;
  assign w_000_284 = r284;
  assign w_000_285 = r285;
  assign w_000_286 = r286;
  assign w_000_287 = r287;
  assign w_000_288 = r288;
  assign w_000_289 = r289;
  assign w_000_290 = r290;
  assign w_000_291 = r291;
  assign w_000_292 = r292;
  assign w_000_293 = r293;
  assign w_000_294 = r294;
  assign w_000_295 = r295;
  assign w_000_296 = r296;
  assign w_000_297 = r297;
  assign w_000_298 = r298;
  assign w_000_299 = r299;
  assign w_000_300 = r300;
  assign w_000_301 = r301;
  assign w_000_302 = r302;
  assign w_000_303 = r303;
  assign w_000_304 = r304;
  assign w_000_305 = r305;
  assign w_000_306 = r306;
  assign w_000_307 = r307;
  assign w_000_308 = r308;
  assign w_000_309 = r309;
  assign w_000_310 = r310;
  assign w_000_311 = r311;
  assign w_000_312 = r312;
  assign w_000_313 = r313;
  assign w_000_314 = r314;
  assign w_000_315 = r315;
  assign w_000_316 = r316;
  assign w_000_317 = r317;
  assign w_000_318 = r318;
  assign w_000_319 = r319;
  assign w_000_320 = r320;
  assign w_000_321 = r321;
  assign w_000_322 = r322;
  assign w_000_323 = r323;
  assign w_000_324 = r324;
  assign w_000_325 = r325;
  assign w_000_326 = r326;
  assign w_000_327 = r327;
  assign w_000_328 = r328;
  assign w_000_329 = r329;
  assign w_000_330 = r330;
  assign w_000_331 = r331;
  assign w_000_332 = r332;
  assign w_000_333 = r333;
  assign w_000_334 = r334;
  assign w_000_335 = r335;
  assign w_000_336 = r336;
  assign w_000_337 = r337;
  assign w_000_338 = r338;
  assign w_000_339 = r339;
  assign w_000_340 = r340;
  assign w_000_341 = r341;
  assign w_000_342 = r342;
  assign w_000_343 = r343;
  assign w_000_344 = r344;
  assign w_000_345 = r345;
  assign w_000_346 = r346;
  assign w_000_347 = r347;
  assign w_000_348 = r348;
  assign w_000_349 = r349;
  assign w_000_350 = r350;
  assign w_000_351 = r351;
  assign w_000_352 = r352;
  assign w_000_353 = r353;
  assign w_000_354 = r354;
  assign w_000_355 = r355;
  assign w_000_356 = r356;
  assign w_000_357 = r357;
  assign w_000_358 = r358;
  assign w_000_359 = r359;
  assign w_000_360 = r360;
  assign w_000_361 = r361;
  assign w_000_362 = r362;
  assign w_000_363 = r363;
  assign w_000_364 = r364;
  assign w_000_365 = r365;
  assign w_000_366 = r366;
  assign w_000_367 = r367;
  assign w_000_368 = r368;
  assign w_000_369 = r369;
  assign w_000_370 = r370;
  assign w_000_371 = r371;
  assign w_000_372 = r372;
  assign w_000_373 = r373;
  assign w_000_374 = r374;
  assign w_000_375 = r375;
  assign w_000_376 = r376;
  assign w_000_377 = r377;
  assign w_000_378 = r378;
  assign w_000_379 = r379;
  assign w_000_380 = r380;
  assign w_000_381 = r381;
  assign w_000_382 = r382;
  assign w_000_383 = r383;
  assign w_000_384 = r384;
  assign w_000_385 = r385;
  assign w_000_386 = r386;
  assign w_000_387 = r387;
  assign w_000_388 = r388;
  assign w_000_389 = r389;
  assign w_000_390 = r390;
  assign w_000_391 = r391;
  assign w_000_392 = r392;
  assign w_000_393 = r393;
  assign w_000_394 = r394;
  assign w_000_395 = r395;
  assign w_000_396 = r396;
  assign w_000_397 = r397;
  assign w_000_398 = r398;
  assign w_000_399 = r399;
  assign w_000_400 = r400;
  assign w_000_401 = r401;
  assign w_000_402 = r402;
  assign w_000_403 = r403;
  assign w_000_404 = r404;
  assign w_000_405 = r405;
  assign w_000_406 = r406;
  assign w_000_407 = r407;
  assign w_000_408 = r408;
  assign w_000_409 = r409;
  assign w_000_410 = r410;
  assign w_000_411 = r411;
  assign w_000_412 = r412;
  assign w_000_413 = r413;
  assign w_000_414 = r414;
  assign w_000_415 = r415;
  assign w_000_416 = r416;
  assign w_000_417 = r417;
  assign w_000_418 = r418;
  assign w_000_419 = r419;
  assign w_000_420 = r420;
  assign w_000_421 = r421;
  assign w_000_422 = r422;
  assign w_000_423 = r423;
  assign w_000_424 = r424;
  assign w_000_425 = r425;
  assign w_000_426 = r426;
  assign w_000_427 = r427;
  assign w_000_428 = r428;
  assign w_000_429 = r429;
  assign w_000_430 = r430;
  assign w_000_431 = r431;
  assign w_000_432 = r432;
  assign w_000_433 = r433;
  assign w_000_434 = r434;
  assign w_000_435 = r435;
  assign w_000_436 = r436;
  assign w_000_437 = r437;
  assign w_000_438 = r438;
  assign w_000_439 = r439;
  assign w_000_440 = r440;
  assign w_000_441 = r441;
  assign w_000_442 = r442;
  assign w_000_443 = r443;
  assign w_000_444 = r444;
  assign w_000_445 = r445;
  assign w_000_446 = r446;
  assign w_000_447 = r447;
  assign w_000_448 = r448;
  assign w_000_449 = r449;
  assign w_000_450 = r450;
  assign w_000_451 = r451;
  assign w_000_452 = r452;
  assign w_000_453 = r453;
  assign w_000_454 = r454;
  assign w_000_455 = r455;
  assign w_000_456 = r456;
  assign w_000_457 = r457;
  assign w_000_458 = r458;
  assign w_000_459 = r459;
  assign w_000_460 = r460;
  assign w_000_461 = r461;
  assign w_000_462 = r462;
  assign w_000_463 = r463;
  assign w_000_464 = r464;
  assign w_000_465 = r465;
  assign w_000_466 = r466;
  assign w_000_467 = r467;
  assign w_000_468 = r468;
  assign w_000_469 = r469;
  assign w_000_470 = r470;
  assign w_000_471 = r471;
  assign w_000_472 = r472;
  assign w_000_473 = r473;
  assign w_000_474 = r474;
  assign w_000_475 = r475;
  assign w_000_476 = r476;
  assign w_000_477 = r477;
  assign w_000_478 = r478;
  assign w_000_479 = r479;
  assign w_000_480 = r480;
  assign w_000_481 = r481;
  assign w_000_482 = r482;
  assign w_000_483 = r483;
  assign w_000_484 = r484;
  assign w_000_485 = r485;
  assign w_000_486 = r486;
  assign w_000_487 = r487;
  assign w_000_488 = r488;
  assign w_000_489 = r489;
  assign w_000_490 = r490;
  assign w_000_491 = r491;
  assign w_000_492 = r492;
  assign w_000_493 = r493;
  assign w_000_494 = r494;
  assign w_000_495 = r495;
  assign w_000_496 = r496;
  assign w_000_497 = r497;
  assign w_000_498 = r498;
  assign w_000_499 = r499;
  assign w_000_500 = r500;
  assign w_000_501 = r501;
  assign w_000_502 = r502;
  assign w_000_503 = r503;
  assign w_000_504 = r504;
  assign w_000_505 = r505;
  assign w_000_506 = r506;
  assign w_000_507 = r507;
  assign w_000_508 = r508;
  assign w_000_509 = r509;
  assign w_000_510 = r510;
  assign w_000_511 = r511;
  assign w_000_512 = r512;
  assign w_000_513 = r513;
  assign w_000_514 = r514;
  assign w_000_515 = r515;
  assign w_000_516 = r516;
  assign w_000_517 = r517;
  assign w_000_518 = r518;
  assign w_000_519 = r519;
  assign w_000_520 = r520;
  assign w_000_521 = r521;
  assign w_000_522 = r522;
  assign w_000_523 = r523;
  assign w_000_524 = r524;
  assign w_000_525 = r525;
  assign w_000_526 = r526;
  assign w_000_527 = r527;
  assign w_000_528 = r528;
  assign w_000_529 = r529;
  assign w_000_530 = r530;
  assign w_000_531 = r531;
  assign w_000_532 = r532;
  assign w_000_533 = r533;
  assign w_000_534 = r534;
  assign w_000_535 = r535;
  assign w_000_536 = r536;
  assign w_000_537 = r537;
  assign w_000_538 = r538;
  assign w_000_539 = r539;
  assign w_000_540 = r540;
  assign w_000_541 = r541;
  assign w_000_542 = r542;
  assign w_000_543 = r543;
  assign w_000_544 = r544;
  assign w_000_545 = r545;
  assign w_000_546 = r546;
  assign w_000_547 = r547;
  assign w_000_548 = r548;
  assign w_000_549 = r549;
  assign w_000_550 = r550;
  assign w_000_551 = r551;
  assign w_000_552 = r552;
  assign w_000_553 = r553;
  assign w_000_554 = r554;
  assign w_000_555 = r555;
  assign w_000_556 = r556;
  assign w_000_557 = r557;
  assign w_000_558 = r558;
  assign w_000_559 = r559;
  assign w_000_560 = r560;
  assign w_000_561 = r561;
  assign w_000_562 = r562;
  assign w_000_563 = r563;
  assign w_000_564 = r564;
  assign w_000_565 = r565;
  assign w_000_566 = r566;
  assign w_000_567 = r567;
  assign w_000_568 = r568;
  assign w_000_569 = r569;
  assign w_000_570 = r570;
  assign w_000_571 = r571;
  assign w_000_572 = r572;
  assign w_000_573 = r573;
  assign w_000_574 = r574;
  assign w_000_575 = r575;
  assign w_000_576 = r576;
  assign w_000_577 = r577;
  assign w_000_578 = r578;
  assign w_000_579 = r579;
  assign w_000_580 = r580;
  assign w_000_581 = r581;
  assign w_000_582 = r582;
  assign w_000_583 = r583;
  assign w_000_584 = r584;
  assign w_000_585 = r585;
  assign w_000_586 = r586;
  assign w_000_587 = r587;
  assign w_000_588 = r588;
  assign w_000_589 = r589;
  assign w_000_590 = r590;
  assign w_000_591 = r591;
  assign w_000_592 = r592;
  assign w_000_593 = r593;
  assign w_000_594 = r594;
  assign w_000_595 = r595;
  assign w_000_596 = r596;
  assign w_000_597 = r597;
  assign w_000_598 = r598;
  assign w_000_599 = r599;
  assign w_000_600 = r600;
  assign w_000_601 = r601;
  assign w_000_602 = r602;
  assign w_000_603 = r603;
  assign w_000_604 = r604;
  assign w_000_605 = r605;
  assign w_000_606 = r606;
  assign w_000_607 = r607;
  assign w_000_608 = r608;
  assign w_000_609 = r609;
  assign w_000_610 = r610;
  assign w_000_611 = r611;
  assign w_000_612 = r612;
  assign w_000_613 = r613;
  assign w_000_614 = r614;
  assign w_000_615 = r615;
  assign w_000_616 = r616;
  assign w_000_617 = r617;
  assign w_000_618 = r618;
  assign w_000_619 = r619;
  assign w_000_620 = r620;
  assign w_000_621 = r621;
  assign w_000_622 = r622;
  assign w_000_623 = r623;
  assign w_000_624 = r624;
  assign w_000_625 = r625;
  assign w_000_626 = r626;
  assign w_000_627 = r627;
  assign w_000_628 = r628;
  assign w_000_629 = r629;
  assign w_000_630 = r630;
  assign w_000_631 = r631;
  assign w_000_632 = r632;
  assign w_000_633 = r633;
  assign w_000_634 = r634;
  assign w_000_635 = r635;
  assign w_000_636 = r636;
  assign w_000_637 = r637;
  assign w_000_638 = r638;
  assign w_000_639 = r639;
  assign w_000_640 = r640;
  assign w_000_641 = r641;
  assign w_000_642 = r642;
  assign w_000_643 = r643;
  assign w_000_644 = r644;
  assign w_000_645 = r645;
  assign w_000_646 = r646;
  assign w_000_647 = r647;
  assign w_000_648 = r648;
  assign w_000_649 = r649;
  assign w_000_650 = r650;
  assign w_000_651 = r651;
  assign w_000_652 = r652;
  assign w_000_653 = r653;
  assign w_000_654 = r654;
  assign w_000_655 = r655;
  assign w_000_656 = r656;
  assign w_000_657 = r657;
  assign w_000_658 = r658;
  assign w_000_659 = r659;
  assign w_000_660 = r660;
  assign w_000_661 = r661;
  assign w_000_662 = r662;
  assign w_000_663 = r663;
  assign w_000_664 = r664;
  assign w_000_665 = r665;
  assign w_000_666 = r666;
  assign w_000_667 = r667;
  assign w_000_668 = r668;
  assign w_000_669 = r669;
  assign w_000_670 = r670;
  assign w_000_671 = r671;
  assign w_000_672 = r672;
  assign w_000_673 = r673;
  assign w_000_674 = r674;
  assign w_000_675 = r675;
  assign w_000_676 = r676;
  assign w_000_677 = r677;
  assign w_000_678 = r678;
  assign w_000_679 = r679;
  assign w_000_680 = r680;
  assign w_000_681 = r681;
  assign w_000_682 = r682;
  assign w_000_683 = r683;
  assign w_000_684 = r684;
  assign w_000_685 = r685;
  assign w_000_686 = r686;
  assign w_000_687 = r687;
  assign w_000_688 = r688;
  assign w_000_689 = r689;
  assign w_000_690 = r690;
  assign w_000_691 = r691;
  assign w_000_692 = r692;
  assign w_000_693 = r693;
  assign w_000_694 = r694;
  assign w_000_695 = r695;
  assign w_000_696 = r696;
  assign w_000_697 = r697;
  assign w_000_698 = r698;
  assign w_000_699 = r699;
  assign w_000_700 = r700;
  assign w_000_701 = r701;
  assign w_000_702 = r702;
  assign w_000_703 = r703;
  assign w_000_704 = r704;
  assign w_000_705 = r705;
  assign w_000_706 = r706;
  assign w_000_707 = r707;
  assign w_000_708 = r708;
  assign w_000_709 = r709;
  assign w_000_710 = r710;
  assign w_000_711 = r711;
  assign w_000_712 = r712;
  assign w_000_713 = r713;
  assign w_000_714 = r714;
  assign w_000_715 = r715;
  assign w_000_716 = r716;
  assign w_000_717 = r717;
  assign w_000_718 = r718;
  assign w_000_719 = r719;
  assign w_000_720 = r720;
  assign w_000_721 = r721;
  assign w_000_722 = r722;
  assign w_000_723 = r723;
  assign w_000_724 = r724;
  assign w_000_725 = r725;
  assign w_000_726 = r726;
  assign w_000_727 = r727;
  assign w_000_728 = r728;
  assign w_000_729 = r729;
  assign w_000_730 = r730;
  assign w_000_731 = r731;
  assign w_000_732 = r732;
  assign w_000_733 = r733;
  assign w_000_734 = r734;
  assign w_000_735 = r735;
  assign w_000_736 = r736;
  assign w_000_737 = r737;
  assign w_000_738 = r738;
  assign w_000_739 = r739;
  assign w_000_740 = r740;
  assign w_000_741 = r741;
  assign w_000_742 = r742;
  assign w_000_743 = r743;
  assign w_000_744 = r744;
  assign w_000_745 = r745;
  assign w_000_746 = r746;
  assign w_000_747 = r747;
  assign w_000_748 = r748;
  assign w_000_749 = r749;
  assign w_000_750 = r750;
  assign w_000_751 = r751;
  assign w_000_752 = r752;
  assign w_000_753 = r753;
  assign w_000_754 = r754;
  assign w_000_755 = r755;
  assign w_000_756 = r756;
  assign w_000_757 = r757;
  assign w_000_758 = r758;
  assign w_000_759 = r759;
  assign w_000_760 = r760;
  assign w_000_761 = r761;
  assign w_000_762 = r762;
  assign w_000_763 = r763;
  assign w_000_764 = r764;
  assign w_000_765 = r765;
  assign w_000_766 = r766;
  assign w_000_767 = r767;
  assign w_000_768 = r768;
  assign w_000_769 = r769;
  assign w_000_770 = r770;
  assign w_000_771 = r771;
  assign w_000_772 = r772;
  assign w_000_773 = r773;
  assign w_000_774 = r774;
  assign w_000_775 = r775;
  assign w_000_776 = r776;
  assign w_000_777 = r777;
  assign w_000_778 = r778;
  assign w_000_779 = r779;
  assign w_000_780 = r780;
  assign w_000_781 = r781;
  assign w_000_782 = r782;
  assign w_000_783 = r783;
  assign w_000_784 = r784;
  assign w_000_785 = r785;
  assign w_000_786 = r786;
  assign w_000_787 = r787;
  assign w_000_788 = r788;
  assign w_000_789 = r789;
  assign w_000_790 = r790;
  assign w_000_791 = r791;
  assign w_000_792 = r792;
  assign w_000_793 = r793;
  assign w_000_794 = r794;
  assign w_000_795 = r795;
  assign w_000_796 = r796;
  assign w_000_797 = r797;

  initial begin 
    r0 = 1'b0; 
    r1 = 1'b0; 
    r2 = 1'b0; 
    r3 = 1'b0; 
    r4 = 1'b0; 
    r5 = 1'b0; 
    r6 = 1'b0; 
    r7 = 1'b0; 
    r8 = 1'b0; 
    r9 = 1'b0; 
    r10 = 1'b0; 
    r11 = 1'b0; 
    r12 = 1'b0; 
    r13 = 1'b0; 
    r14 = 1'b0; 
    r15 = 1'b0; 
    r16 = 1'b0; 
    r17 = 1'b0; 
    r18 = 1'b0; 
    r19 = 1'b0; 
    r20 = 1'b0; 
    r21 = 1'b0; 
    r22 = 1'b0; 
    r23 = 1'b0; 
    r24 = 1'b0; 
    r25 = 1'b0; 
    r26 = 1'b0; 
    r27 = 1'b0; 
    r28 = 1'b0; 
    r29 = 1'b0; 
    r30 = 1'b0; 
    r31 = 1'b0; 
    r32 = 1'b0; 
    r33 = 1'b0; 
    r34 = 1'b0; 
    r35 = 1'b0; 
    r36 = 1'b0; 
    r37 = 1'b0; 
    r38 = 1'b0; 
    r39 = 1'b0; 
    r40 = 1'b0; 
    r41 = 1'b0; 
    r42 = 1'b0; 
    r43 = 1'b0; 
    r44 = 1'b0; 
    r45 = 1'b0; 
    r46 = 1'b0; 
    r47 = 1'b0; 
    r48 = 1'b0; 
    r49 = 1'b0; 
    r50 = 1'b0; 
    r51 = 1'b0; 
    r52 = 1'b0; 
    r53 = 1'b0; 
    r54 = 1'b0; 
    r55 = 1'b0; 
    r56 = 1'b0; 
    r57 = 1'b0; 
    r58 = 1'b0; 
    r59 = 1'b0; 
    r60 = 1'b0; 
    r61 = 1'b0; 
    r62 = 1'b0; 
    r63 = 1'b0; 
    r64 = 1'b0; 
    r65 = 1'b0; 
    r66 = 1'b0; 
    r67 = 1'b0; 
    r68 = 1'b0; 
    r69 = 1'b0; 
    r70 = 1'b0; 
    r71 = 1'b0; 
    r72 = 1'b0; 
    r73 = 1'b0; 
    r74 = 1'b0; 
    r75 = 1'b0; 
    r76 = 1'b0; 
    r77 = 1'b0; 
    r78 = 1'b0; 
    r79 = 1'b0; 
    r80 = 1'b0; 
    r81 = 1'b0; 
    r82 = 1'b0; 
    r83 = 1'b0; 
    r84 = 1'b0; 
    r85 = 1'b0; 
    r86 = 1'b0; 
    r87 = 1'b0; 
    r88 = 1'b0; 
    r89 = 1'b0; 
    r90 = 1'b0; 
    r91 = 1'b0; 
    r92 = 1'b0; 
    r93 = 1'b0; 
    r94 = 1'b0; 
    r95 = 1'b0; 
    r96 = 1'b0; 
    r97 = 1'b0; 
    r98 = 1'b0; 
    r99 = 1'b0; 
    r100 = 1'b0; 
    r101 = 1'b0; 
    r102 = 1'b0; 
    r103 = 1'b0; 
    r104 = 1'b0; 
    r105 = 1'b0; 
    r106 = 1'b0; 
    r107 = 1'b0; 
    r108 = 1'b0; 
    r109 = 1'b0; 
    r110 = 1'b0; 
    r111 = 1'b0; 
    r112 = 1'b0; 
    r113 = 1'b0; 
    r114 = 1'b0; 
    r115 = 1'b0; 
    r116 = 1'b0; 
    r117 = 1'b0; 
    r118 = 1'b0; 
    r119 = 1'b0; 
    r120 = 1'b0; 
    r121 = 1'b0; 
    r122 = 1'b0; 
    r123 = 1'b0; 
    r124 = 1'b0; 
    r125 = 1'b0; 
    r126 = 1'b0; 
    r127 = 1'b0; 
    r128 = 1'b0; 
    r129 = 1'b0; 
    r130 = 1'b0; 
    r131 = 1'b0; 
    r132 = 1'b0; 
    r133 = 1'b0; 
    r134 = 1'b0; 
    r135 = 1'b0; 
    r136 = 1'b0; 
    r137 = 1'b0; 
    r138 = 1'b0; 
    r139 = 1'b0; 
    r140 = 1'b0; 
    r141 = 1'b0; 
    r142 = 1'b0; 
    r143 = 1'b0; 
    r144 = 1'b0; 
    r145 = 1'b0; 
    r146 = 1'b0; 
    r147 = 1'b0; 
    r148 = 1'b0; 
    r149 = 1'b0; 
    r150 = 1'b0; 
    r151 = 1'b0; 
    r152 = 1'b0; 
    r153 = 1'b0; 
    r154 = 1'b0; 
    r155 = 1'b0; 
    r156 = 1'b0; 
    r157 = 1'b0; 
    r158 = 1'b0; 
    r159 = 1'b0; 
    r160 = 1'b0; 
    r161 = 1'b0; 
    r162 = 1'b0; 
    r163 = 1'b0; 
    r164 = 1'b0; 
    r165 = 1'b0; 
    r166 = 1'b0; 
    r167 = 1'b0; 
    r168 = 1'b0; 
    r169 = 1'b0; 
    r170 = 1'b0; 
    r171 = 1'b0; 
    r172 = 1'b0; 
    r173 = 1'b0; 
    r174 = 1'b0; 
    r175 = 1'b0; 
    r176 = 1'b0; 
    r177 = 1'b0; 
    r178 = 1'b0; 
    r179 = 1'b0; 
    r180 = 1'b0; 
    r181 = 1'b0; 
    r182 = 1'b0; 
    r183 = 1'b0; 
    r184 = 1'b0; 
    r185 = 1'b0; 
    r186 = 1'b0; 
    r187 = 1'b0; 
    r188 = 1'b0; 
    r189 = 1'b0; 
    r190 = 1'b0; 
    r191 = 1'b0; 
    r192 = 1'b0; 
    r193 = 1'b0; 
    r194 = 1'b0; 
    r195 = 1'b0; 
    r196 = 1'b0; 
    r197 = 1'b0; 
    r198 = 1'b0; 
    r199 = 1'b0; 
    r200 = 1'b0; 
    r201 = 1'b0; 
    r202 = 1'b0; 
    r203 = 1'b0; 
    r204 = 1'b0; 
    r205 = 1'b0; 
    r206 = 1'b0; 
    r207 = 1'b0; 
    r208 = 1'b0; 
    r209 = 1'b0; 
    r210 = 1'b0; 
    r211 = 1'b0; 
    r212 = 1'b0; 
    r213 = 1'b0; 
    r214 = 1'b0; 
    r215 = 1'b0; 
    r216 = 1'b0; 
    r217 = 1'b0; 
    r218 = 1'b0; 
    r219 = 1'b0; 
    r220 = 1'b0; 
    r221 = 1'b0; 
    r222 = 1'b0; 
    r223 = 1'b0; 
    r224 = 1'b0; 
    r225 = 1'b0; 
    r226 = 1'b0; 
    r227 = 1'b0; 
    r228 = 1'b0; 
    r229 = 1'b0; 
    r230 = 1'b0; 
    r231 = 1'b0; 
    r232 = 1'b0; 
    r233 = 1'b0; 
    r234 = 1'b0; 
    r235 = 1'b0; 
    r236 = 1'b0; 
    r237 = 1'b0; 
    r238 = 1'b0; 
    r239 = 1'b0; 
    r240 = 1'b0; 
    r241 = 1'b0; 
    r242 = 1'b0; 
    r243 = 1'b0; 
    r244 = 1'b0; 
    r245 = 1'b0; 
    r246 = 1'b0; 
    r247 = 1'b0; 
    r248 = 1'b0; 
    r249 = 1'b0; 
    r250 = 1'b0; 
    r251 = 1'b0; 
    r252 = 1'b0; 
    r253 = 1'b0; 
    r254 = 1'b0; 
    r255 = 1'b0; 
    r256 = 1'b0; 
    r257 = 1'b0; 
    r258 = 1'b0; 
    r259 = 1'b0; 
    r260 = 1'b0; 
    r261 = 1'b0; 
    r262 = 1'b0; 
    r263 = 1'b0; 
    r264 = 1'b0; 
    r265 = 1'b0; 
    r266 = 1'b0; 
    r267 = 1'b0; 
    r268 = 1'b0; 
    r269 = 1'b0; 
    r270 = 1'b0; 
    r271 = 1'b0; 
    r272 = 1'b0; 
    r273 = 1'b0; 
    r274 = 1'b0; 
    r275 = 1'b0; 
    r276 = 1'b0; 
    r277 = 1'b0; 
    r278 = 1'b0; 
    r279 = 1'b0; 
    r280 = 1'b0; 
    r281 = 1'b0; 
    r282 = 1'b0; 
    r283 = 1'b0; 
    r284 = 1'b0; 
    r285 = 1'b0; 
    r286 = 1'b0; 
    r287 = 1'b0; 
    r288 = 1'b0; 
    r289 = 1'b0; 
    r290 = 1'b0; 
    r291 = 1'b0; 
    r292 = 1'b0; 
    r293 = 1'b0; 
    r294 = 1'b0; 
    r295 = 1'b0; 
    r296 = 1'b0; 
    r297 = 1'b0; 
    r298 = 1'b0; 
    r299 = 1'b0; 
    r300 = 1'b0; 
    r301 = 1'b0; 
    r302 = 1'b0; 
    r303 = 1'b0; 
    r304 = 1'b0; 
    r305 = 1'b0; 
    r306 = 1'b0; 
    r307 = 1'b0; 
    r308 = 1'b0; 
    r309 = 1'b0; 
    r310 = 1'b0; 
    r311 = 1'b0; 
    r312 = 1'b0; 
    r313 = 1'b0; 
    r314 = 1'b0; 
    r315 = 1'b0; 
    r316 = 1'b0; 
    r317 = 1'b0; 
    r318 = 1'b0; 
    r319 = 1'b0; 
    r320 = 1'b0; 
    r321 = 1'b0; 
    r322 = 1'b0; 
    r323 = 1'b0; 
    r324 = 1'b0; 
    r325 = 1'b0; 
    r326 = 1'b0; 
    r327 = 1'b0; 
    r328 = 1'b0; 
    r329 = 1'b0; 
    r330 = 1'b0; 
    r331 = 1'b0; 
    r332 = 1'b0; 
    r333 = 1'b0; 
    r334 = 1'b0; 
    r335 = 1'b0; 
    r336 = 1'b0; 
    r337 = 1'b0; 
    r338 = 1'b0; 
    r339 = 1'b0; 
    r340 = 1'b0; 
    r341 = 1'b0; 
    r342 = 1'b0; 
    r343 = 1'b0; 
    r344 = 1'b0; 
    r345 = 1'b0; 
    r346 = 1'b0; 
    r347 = 1'b0; 
    r348 = 1'b0; 
    r349 = 1'b0; 
    r350 = 1'b0; 
    r351 = 1'b0; 
    r352 = 1'b0; 
    r353 = 1'b0; 
    r354 = 1'b0; 
    r355 = 1'b0; 
    r356 = 1'b0; 
    r357 = 1'b0; 
    r358 = 1'b0; 
    r359 = 1'b0; 
    r360 = 1'b0; 
    r361 = 1'b0; 
    r362 = 1'b0; 
    r363 = 1'b0; 
    r364 = 1'b0; 
    r365 = 1'b0; 
    r366 = 1'b0; 
    r367 = 1'b0; 
    r368 = 1'b0; 
    r369 = 1'b0; 
    r370 = 1'b0; 
    r371 = 1'b0; 
    r372 = 1'b0; 
    r373 = 1'b0; 
    r374 = 1'b0; 
    r375 = 1'b0; 
    r376 = 1'b0; 
    r377 = 1'b0; 
    r378 = 1'b0; 
    r379 = 1'b0; 
    r380 = 1'b0; 
    r381 = 1'b0; 
    r382 = 1'b0; 
    r383 = 1'b0; 
    r384 = 1'b0; 
    r385 = 1'b0; 
    r386 = 1'b0; 
    r387 = 1'b0; 
    r388 = 1'b0; 
    r389 = 1'b0; 
    r390 = 1'b0; 
    r391 = 1'b0; 
    r392 = 1'b0; 
    r393 = 1'b0; 
    r394 = 1'b0; 
    r395 = 1'b0; 
    r396 = 1'b0; 
    r397 = 1'b0; 
    r398 = 1'b0; 
    r399 = 1'b0; 
    r400 = 1'b0; 
    r401 = 1'b0; 
    r402 = 1'b0; 
    r403 = 1'b0; 
    r404 = 1'b0; 
    r405 = 1'b0; 
    r406 = 1'b0; 
    r407 = 1'b0; 
    r408 = 1'b0; 
    r409 = 1'b0; 
    r410 = 1'b0; 
    r411 = 1'b0; 
    r412 = 1'b0; 
    r413 = 1'b0; 
    r414 = 1'b0; 
    r415 = 1'b0; 
    r416 = 1'b0; 
    r417 = 1'b0; 
    r418 = 1'b0; 
    r419 = 1'b0; 
    r420 = 1'b0; 
    r421 = 1'b0; 
    r422 = 1'b0; 
    r423 = 1'b0; 
    r424 = 1'b0; 
    r425 = 1'b0; 
    r426 = 1'b0; 
    r427 = 1'b0; 
    r428 = 1'b0; 
    r429 = 1'b0; 
    r430 = 1'b0; 
    r431 = 1'b0; 
    r432 = 1'b0; 
    r433 = 1'b0; 
    r434 = 1'b0; 
    r435 = 1'b0; 
    r436 = 1'b0; 
    r437 = 1'b0; 
    r438 = 1'b0; 
    r439 = 1'b0; 
    r440 = 1'b0; 
    r441 = 1'b0; 
    r442 = 1'b0; 
    r443 = 1'b0; 
    r444 = 1'b0; 
    r445 = 1'b0; 
    r446 = 1'b0; 
    r447 = 1'b0; 
    r448 = 1'b0; 
    r449 = 1'b0; 
    r450 = 1'b0; 
    r451 = 1'b0; 
    r452 = 1'b0; 
    r453 = 1'b0; 
    r454 = 1'b0; 
    r455 = 1'b0; 
    r456 = 1'b0; 
    r457 = 1'b0; 
    r458 = 1'b0; 
    r459 = 1'b0; 
    r460 = 1'b0; 
    r461 = 1'b0; 
    r462 = 1'b0; 
    r463 = 1'b0; 
    r464 = 1'b0; 
    r465 = 1'b0; 
    r466 = 1'b0; 
    r467 = 1'b0; 
    r468 = 1'b0; 
    r469 = 1'b0; 
    r470 = 1'b0; 
    r471 = 1'b0; 
    r472 = 1'b0; 
    r473 = 1'b0; 
    r474 = 1'b0; 
    r475 = 1'b0; 
    r476 = 1'b0; 
    r477 = 1'b0; 
    r478 = 1'b0; 
    r479 = 1'b0; 
    r480 = 1'b0; 
    r481 = 1'b0; 
    r482 = 1'b0; 
    r483 = 1'b0; 
    r484 = 1'b0; 
    r485 = 1'b0; 
    r486 = 1'b0; 
    r487 = 1'b0; 
    r488 = 1'b0; 
    r489 = 1'b0; 
    r490 = 1'b0; 
    r491 = 1'b0; 
    r492 = 1'b0; 
    r493 = 1'b0; 
    r494 = 1'b0; 
    r495 = 1'b0; 
    r496 = 1'b0; 
    r497 = 1'b0; 
    r498 = 1'b0; 
    r499 = 1'b0; 
    r500 = 1'b0; 
    r501 = 1'b0; 
    r502 = 1'b0; 
    r503 = 1'b0; 
    r504 = 1'b0; 
    r505 = 1'b0; 
    r506 = 1'b0; 
    r507 = 1'b0; 
    r508 = 1'b0; 
    r509 = 1'b0; 
    r510 = 1'b0; 
    r511 = 1'b0; 
    r512 = 1'b0; 
    r513 = 1'b0; 
    r514 = 1'b0; 
    r515 = 1'b0; 
    r516 = 1'b0; 
    r517 = 1'b0; 
    r518 = 1'b0; 
    r519 = 1'b0; 
    r520 = 1'b0; 
    r521 = 1'b0; 
    r522 = 1'b0; 
    r523 = 1'b0; 
    r524 = 1'b0; 
    r525 = 1'b0; 
    r526 = 1'b0; 
    r527 = 1'b0; 
    r528 = 1'b0; 
    r529 = 1'b0; 
    r530 = 1'b0; 
    r531 = 1'b0; 
    r532 = 1'b0; 
    r533 = 1'b0; 
    r534 = 1'b0; 
    r535 = 1'b0; 
    r536 = 1'b0; 
    r537 = 1'b0; 
    r538 = 1'b0; 
    r539 = 1'b0; 
    r540 = 1'b0; 
    r541 = 1'b0; 
    r542 = 1'b0; 
    r543 = 1'b0; 
    r544 = 1'b0; 
    r545 = 1'b0; 
    r546 = 1'b0; 
    r547 = 1'b0; 
    r548 = 1'b0; 
    r549 = 1'b0; 
    r550 = 1'b0; 
    r551 = 1'b0; 
    r552 = 1'b0; 
    r553 = 1'b0; 
    r554 = 1'b0; 
    r555 = 1'b0; 
    r556 = 1'b0; 
    r557 = 1'b0; 
    r558 = 1'b0; 
    r559 = 1'b0; 
    r560 = 1'b0; 
    r561 = 1'b0; 
    r562 = 1'b0; 
    r563 = 1'b0; 
    r564 = 1'b0; 
    r565 = 1'b0; 
    r566 = 1'b0; 
    r567 = 1'b0; 
    r568 = 1'b0; 
    r569 = 1'b0; 
    r570 = 1'b0; 
    r571 = 1'b0; 
    r572 = 1'b0; 
    r573 = 1'b0; 
    r574 = 1'b0; 
    r575 = 1'b0; 
    r576 = 1'b0; 
    r577 = 1'b0; 
    r578 = 1'b0; 
    r579 = 1'b0; 
    r580 = 1'b0; 
    r581 = 1'b0; 
    r582 = 1'b0; 
    r583 = 1'b0; 
    r584 = 1'b0; 
    r585 = 1'b0; 
    r586 = 1'b0; 
    r587 = 1'b0; 
    r588 = 1'b0; 
    r589 = 1'b0; 
    r590 = 1'b0; 
    r591 = 1'b0; 
    r592 = 1'b0; 
    r593 = 1'b0; 
    r594 = 1'b0; 
    r595 = 1'b0; 
    r596 = 1'b0; 
    r597 = 1'b0; 
    r598 = 1'b0; 
    r599 = 1'b0; 
    r600 = 1'b0; 
    r601 = 1'b0; 
    r602 = 1'b0; 
    r603 = 1'b0; 
    r604 = 1'b0; 
    r605 = 1'b0; 
    r606 = 1'b0; 
    r607 = 1'b0; 
    r608 = 1'b0; 
    r609 = 1'b0; 
    r610 = 1'b0; 
    r611 = 1'b0; 
    r612 = 1'b0; 
    r613 = 1'b0; 
    r614 = 1'b0; 
    r615 = 1'b0; 
    r616 = 1'b0; 
    r617 = 1'b0; 
    r618 = 1'b0; 
    r619 = 1'b0; 
    r620 = 1'b0; 
    r621 = 1'b0; 
    r622 = 1'b0; 
    r623 = 1'b0; 
    r624 = 1'b0; 
    r625 = 1'b0; 
    r626 = 1'b0; 
    r627 = 1'b0; 
    r628 = 1'b0; 
    r629 = 1'b0; 
    r630 = 1'b0; 
    r631 = 1'b0; 
    r632 = 1'b0; 
    r633 = 1'b0; 
    r634 = 1'b0; 
    r635 = 1'b0; 
    r636 = 1'b0; 
    r637 = 1'b0; 
    r638 = 1'b0; 
    r639 = 1'b0; 
    r640 = 1'b0; 
    r641 = 1'b0; 
    r642 = 1'b0; 
    r643 = 1'b0; 
    r644 = 1'b0; 
    r645 = 1'b0; 
    r646 = 1'b0; 
    r647 = 1'b0; 
    r648 = 1'b0; 
    r649 = 1'b0; 
    r650 = 1'b0; 
    r651 = 1'b0; 
    r652 = 1'b0; 
    r653 = 1'b0; 
    r654 = 1'b0; 
    r655 = 1'b0; 
    r656 = 1'b0; 
    r657 = 1'b0; 
    r658 = 1'b0; 
    r659 = 1'b0; 
    r660 = 1'b0; 
    r661 = 1'b0; 
    r662 = 1'b0; 
    r663 = 1'b0; 
    r664 = 1'b0; 
    r665 = 1'b0; 
    r666 = 1'b0; 
    r667 = 1'b0; 
    r668 = 1'b0; 
    r669 = 1'b0; 
    r670 = 1'b0; 
    r671 = 1'b0; 
    r672 = 1'b0; 
    r673 = 1'b0; 
    r674 = 1'b0; 
    r675 = 1'b0; 
    r676 = 1'b0; 
    r677 = 1'b0; 
    r678 = 1'b0; 
    r679 = 1'b0; 
    r680 = 1'b0; 
    r681 = 1'b0; 
    r682 = 1'b0; 
    r683 = 1'b0; 
    r684 = 1'b0; 
    r685 = 1'b0; 
    r686 = 1'b0; 
    r687 = 1'b0; 
    r688 = 1'b0; 
    r689 = 1'b0; 
    r690 = 1'b0; 
    r691 = 1'b0; 
    r692 = 1'b0; 
    r693 = 1'b0; 
    r694 = 1'b0; 
    r695 = 1'b0; 
    r696 = 1'b0; 
    r697 = 1'b0; 
    r698 = 1'b0; 
    r699 = 1'b0; 
    r700 = 1'b0; 
    r701 = 1'b0; 
    r702 = 1'b0; 
    r703 = 1'b0; 
    r704 = 1'b0; 
    r705 = 1'b0; 
    r706 = 1'b0; 
    r707 = 1'b0; 
    r708 = 1'b0; 
    r709 = 1'b0; 
    r710 = 1'b0; 
    r711 = 1'b0; 
    r712 = 1'b0; 
    r713 = 1'b0; 
    r714 = 1'b0; 
    r715 = 1'b0; 
    r716 = 1'b0; 
    r717 = 1'b0; 
    r718 = 1'b0; 
    r719 = 1'b0; 
    r720 = 1'b0; 
    r721 = 1'b0; 
    r722 = 1'b0; 
    r723 = 1'b0; 
    r724 = 1'b0; 
    r725 = 1'b0; 
    r726 = 1'b0; 
    r727 = 1'b0; 
    r728 = 1'b0; 
    r729 = 1'b0; 
    r730 = 1'b0; 
    r731 = 1'b0; 
    r732 = 1'b0; 
    r733 = 1'b0; 
    r734 = 1'b0; 
    r735 = 1'b0; 
    r736 = 1'b0; 
    r737 = 1'b0; 
    r738 = 1'b0; 
    r739 = 1'b0; 
    r740 = 1'b0; 
    r741 = 1'b0; 
    r742 = 1'b0; 
    r743 = 1'b0; 
    r744 = 1'b0; 
    r745 = 1'b0; 
    r746 = 1'b0; 
    r747 = 1'b0; 
    r748 = 1'b0; 
    r749 = 1'b0; 
    r750 = 1'b0; 
    r751 = 1'b0; 
    r752 = 1'b0; 
    r753 = 1'b0; 
    r754 = 1'b0; 
    r755 = 1'b0; 
    r756 = 1'b0; 
    r757 = 1'b0; 
    r758 = 1'b0; 
    r759 = 1'b0; 
    r760 = 1'b0; 
    r761 = 1'b0; 
    r762 = 1'b0; 
    r763 = 1'b0; 
    r764 = 1'b0; 
    r765 = 1'b0; 
    r766 = 1'b0; 
    r767 = 1'b0; 
    r768 = 1'b0; 
    r769 = 1'b0; 
    r770 = 1'b0; 
    r771 = 1'b0; 
    r772 = 1'b0; 
    r773 = 1'b0; 
    r774 = 1'b0; 
    r775 = 1'b0; 
    r776 = 1'b0; 
    r777 = 1'b0; 
    r778 = 1'b0; 
    r779 = 1'b0; 
    r780 = 1'b0; 
    r781 = 1'b0; 
    r782 = 1'b0; 
    r783 = 1'b0; 
    r784 = 1'b0; 
    r785 = 1'b0; 
    r786 = 1'b0; 
    r787 = 1'b0; 
    r788 = 1'b0; 
    r789 = 1'b0; 
    r790 = 1'b0; 
    r791 = 1'b0; 
    r792 = 1'b0; 
    r793 = 1'b0; 
    r794 = 1'b0; 
    r795 = 1'b0; 
    r796 = 1'b0; 
    r797 = 1'b0; 
    $monitor("%t %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b  ", $time, w_000_000, w_000_001, w_000_002, w_000_003, w_000_004, w_000_005, w_000_006, w_000_007, w_000_008, w_000_009, w_000_010, w_000_011, w_000_012, w_000_013, w_000_014, w_000_015, w_000_016, w_000_017, w_000_018, w_000_019, w_000_020, w_000_021, w_000_022, w_000_023, w_000_024, w_000_025, w_000_026, w_000_027, w_000_028, w_000_029, w_000_030, w_000_031, w_000_032, w_000_033, w_000_034, w_000_035, w_000_036, w_000_037, w_000_038, w_000_039, w_000_040, w_000_041, w_000_042, w_000_043, w_000_044, w_000_045, w_000_046, w_000_047, w_000_048, w_000_049, w_000_050, w_000_051, w_000_052, w_000_053, w_000_054, w_000_055, w_000_056, w_000_057, w_000_058, w_000_059, w_000_060, w_000_061, w_000_062, w_000_063, w_000_064, w_000_065, w_000_066, w_000_067, w_000_068, w_000_069, w_000_070, w_000_071, w_000_072, w_000_073, w_000_074, w_000_075, w_000_076, w_000_077, w_000_078, w_000_079, w_000_080, w_000_081, w_000_082, w_000_083, w_000_084, w_000_085, w_000_086, w_000_087, w_000_088, w_000_089, w_000_090, w_000_091, w_000_092, w_000_093, w_000_094, w_000_095, w_000_096, w_000_097, w_000_098, w_000_099, w_000_100, w_000_101, w_000_102, w_000_103, w_000_104, w_000_105, w_000_106, w_000_107, w_000_108, w_000_109, w_000_110, w_000_111, w_000_112, w_000_113, w_000_114, w_000_115, w_000_116, w_000_117, w_000_118, w_000_119, w_000_120, w_000_121, w_000_122, w_000_123, w_000_124, w_000_125, w_000_126, w_000_127, w_000_128, w_000_129, w_000_130, w_000_131, w_000_132, w_000_133, w_000_134, w_000_135, w_000_136, w_000_137, w_000_138, w_000_139, w_000_140, w_000_141, w_000_142, w_000_143, w_000_144, w_000_145, w_000_146, w_000_147, w_000_148, w_000_149, w_000_150, w_000_151, w_000_152, w_000_153, w_000_154, w_000_155, w_000_156, w_000_157, w_000_158, w_000_159, w_000_160, w_000_161, w_000_162, w_000_163, w_000_164, w_000_165, w_000_166, w_000_167, w_000_168, w_000_169, w_000_170, w_000_171, w_000_172, w_000_173, w_000_174, w_000_175, w_000_176, w_000_177, w_000_178, w_000_179, w_000_180, w_000_181, w_000_182, w_000_183, w_000_184, w_000_185, w_000_186, w_000_187, w_000_188, w_000_189, w_000_190, w_000_191, w_000_192, w_000_193, w_000_194, w_000_195, w_000_196, w_000_197, w_000_198, w_000_199, w_000_200, w_000_201, w_000_202, w_000_203, w_000_204, w_000_205, w_000_206, w_000_207, w_000_208, w_000_209, w_000_210, w_000_211, w_000_212, w_000_213, w_000_214, w_000_215, w_000_216, w_000_217, w_000_218, w_000_219, w_000_220, w_000_221, w_000_222, w_000_223, w_000_224, w_000_225, w_000_226, w_000_227, w_000_228, w_000_229, w_000_230, w_000_231, w_000_232, w_000_233, w_000_234, w_000_235, w_000_236, w_000_237, w_000_238, w_000_239, w_000_240, w_000_241, w_000_242, w_000_243, w_000_244, w_000_245, w_000_246, w_000_247, w_000_248, w_000_249, w_000_250, w_000_251, w_000_252, w_000_253, w_000_254, w_000_255, w_000_256, w_000_257, w_000_258, w_000_259, w_000_260, w_000_261, w_000_262, w_000_263, w_000_264, w_000_265, w_000_266, w_000_267, w_000_268, w_000_269, w_000_270, w_000_271, w_000_272, w_000_273, w_000_274, w_000_275, w_000_276, w_000_277, w_000_278, w_000_279, w_000_280, w_000_281, w_000_282, w_000_283, w_000_284, w_000_285, w_000_286, w_000_287, w_000_288, w_000_289, w_000_290, w_000_291, w_000_292, w_000_293, w_000_294, w_000_295, w_000_296, w_000_297, w_000_298, w_000_299, w_000_300, w_000_301, w_000_302, w_000_303, w_000_304, w_000_305, w_000_306, w_000_307, w_000_308, w_000_309, w_000_310, w_000_311, w_000_312, w_000_313, w_000_314, w_000_315, w_000_316, w_000_317, w_000_318, w_000_319, w_000_320, w_000_321, w_000_322, w_000_323, w_000_324, w_000_325, w_000_326, w_000_327, w_000_328, w_000_329, w_000_330, w_000_331, w_000_332, w_000_333, w_000_334, w_000_335, w_000_336, w_000_337, w_000_338, w_000_339, w_000_340, w_000_341, w_000_342, w_000_343, w_000_344, w_000_345, w_000_346, w_000_347, w_000_348, w_000_349, w_000_350, w_000_351, w_000_352, w_000_353, w_000_354, w_000_355, w_000_356, w_000_357, w_000_358, w_000_359, w_000_360, w_000_361, w_000_362, w_000_363, w_000_364, w_000_365, w_000_366, w_000_367, w_000_368, w_000_369, w_000_370, w_000_371, w_000_372, w_000_373, w_000_374, w_000_375, w_000_376, w_000_377, w_000_378, w_000_379, w_000_380, w_000_381, w_000_382, w_000_383, w_000_384, w_000_385, w_000_386, w_000_387, w_000_388, w_000_389, w_000_390, w_000_391, w_000_392, w_000_393, w_000_394, w_000_395, w_000_396, w_000_397, w_000_398, w_000_399, w_000_400, w_000_401, w_000_402, w_000_403, w_000_404, w_000_405, w_000_406, w_000_407, w_000_408, w_000_409, w_000_410, w_000_411, w_000_412, w_000_413, w_000_414, w_000_415, w_000_416, w_000_417, w_000_418, w_000_419, w_000_420, w_000_421, w_000_422, w_000_423, w_000_424, w_000_425, w_000_426, w_000_427, w_000_428, w_000_429, w_000_430, w_000_431, w_000_432, w_000_433, w_000_434, w_000_435, w_000_436, w_000_437, w_000_438, w_000_439, w_000_440, w_000_441, w_000_442, w_000_443, w_000_444, w_000_445, w_000_446, w_000_447, w_000_448, w_000_449, w_000_450, w_000_451, w_000_452, w_000_453, w_000_454, w_000_455, w_000_456, w_000_457, w_000_458, w_000_459, w_000_460, w_000_461, w_000_462, w_000_463, w_000_464, w_000_465, w_000_466, w_000_467, w_000_468, w_000_469, w_000_470, w_000_471, w_000_472, w_000_473, w_000_474, w_000_475, w_000_476, w_000_477, w_000_478, w_000_479, w_000_480, w_000_481, w_000_482, w_000_483, w_000_484, w_000_485, w_000_486, w_000_487, w_000_488, w_000_489, w_000_490, w_000_491, w_000_492, w_000_493, w_000_494, w_000_495, w_000_496, w_000_497, w_000_498, w_000_499, w_000_500, w_000_501, w_000_502, w_000_503, w_000_504, w_000_505, w_000_506, w_000_507, w_000_508, w_000_509, w_000_510, w_000_511, w_000_512, w_000_513, w_000_514, w_000_515, w_000_516, w_000_517, w_000_518, w_000_519, w_000_520, w_000_521, w_000_522, w_000_523, w_000_524, w_000_525, w_000_526, w_000_527, w_000_528, w_000_529, w_000_530, w_000_531, w_000_532, w_000_533, w_000_534, w_000_535, w_000_536, w_000_537, w_000_538, w_000_539, w_000_540, w_000_541, w_000_542, w_000_543, w_000_544, w_000_545, w_000_546, w_000_547, w_000_548, w_000_549, w_000_550, w_000_551, w_000_552, w_000_553, w_000_554, w_000_555, w_000_556, w_000_557, w_000_558, w_000_559, w_000_560, w_000_561, w_000_562, w_000_563, w_000_564, w_000_565, w_000_566, w_000_567, w_000_568, w_000_569, w_000_570, w_000_571, w_000_572, w_000_573, w_000_574, w_000_575, w_000_576, w_000_577, w_000_578, w_000_579, w_000_580, w_000_581, w_000_582, w_000_583, w_000_584, w_000_585, w_000_586, w_000_587, w_000_588, w_000_589, w_000_590, w_000_591, w_000_592, w_000_593, w_000_594, w_000_595, w_000_596, w_000_597, w_000_598, w_000_599, w_000_600, w_000_601, w_000_602, w_000_603, w_000_604, w_000_605, w_000_606, w_000_607, w_000_608, w_000_609, w_000_610, w_000_611, w_000_612, w_000_613, w_000_614, w_000_615, w_000_616, w_000_617, w_000_618, w_000_619, w_000_620, w_000_621, w_000_622, w_000_623, w_000_624, w_000_625, w_000_626, w_000_627, w_000_628, w_000_629, w_000_630, w_000_631, w_000_632, w_000_633, w_000_634, w_000_635, w_000_636, w_000_637, w_000_638, w_000_639, w_000_640, w_000_641, w_000_642, w_000_643, w_000_644, w_000_645, w_000_646, w_000_647, w_000_648, w_000_649, w_000_650, w_000_651, w_000_652, w_000_653, w_000_654, w_000_655, w_000_656, w_000_657, w_000_658, w_000_659, w_000_660, w_000_661, w_000_662, w_000_663, w_000_664, w_000_665, w_000_666, w_000_667, w_000_668, w_000_669, w_000_670, w_000_671, w_000_672, w_000_673, w_000_674, w_000_675, w_000_676, w_000_677, w_000_678, w_000_679, w_000_680, w_000_681, w_000_682, w_000_683, w_000_684, w_000_685, w_000_686, w_000_687, w_000_688, w_000_689, w_000_690, w_000_691, w_000_692, w_000_693, w_000_694, w_000_695, w_000_696, w_000_697, w_000_698, w_000_699, w_000_700, w_000_701, w_000_702, w_000_703, w_000_704, w_000_705, w_000_706, w_000_707, w_000_708, w_000_709, w_000_710, w_000_711, w_000_712, w_000_713, w_000_714, w_000_715, w_000_716, w_000_717, w_000_718, w_000_719, w_000_720, w_000_721, w_000_722, w_000_723, w_000_724, w_000_725, w_000_726, w_000_727, w_000_728, w_000_729, w_000_730, w_000_731, w_000_732, w_000_733, w_000_734, w_000_735, w_000_736, w_000_737, w_000_738, w_000_739, w_000_740, w_000_741, w_000_742, w_000_743, w_000_744, w_000_745, w_000_746, w_000_747, w_000_748, w_000_749, w_000_750, w_000_751, w_000_752, w_000_753, w_000_754, w_000_755, w_000_756, w_000_757, w_000_758, w_000_759, w_000_760, w_000_761, w_000_762, w_000_763, w_000_764, w_000_765, w_000_766, w_000_767, w_000_768, w_000_769, w_000_770, w_000_771, w_000_772, w_000_773, w_000_774, w_000_775, w_000_776, w_000_777, w_000_778, w_000_779, w_000_780, w_000_781, w_000_782, w_000_783, w_000_784, w_000_785, w_000_786, w_000_787, w_000_788, w_000_789, w_000_790, w_000_791, w_000_792, w_000_793, w_000_794, w_000_795, w_000_796, w_000_797, w_800_000, w_800_001, w_800_002, w_800_003, w_800_004, w_800_005, w_800_006, w_800_007, w_800_008, w_800_009, w_800_010, w_800_011, w_800_012, w_800_013, w_800_014, w_800_015, w_800_016, w_800_017, w_800_018, w_800_019, w_800_020, w_800_021, w_800_022, w_800_023, w_800_024, w_800_025, w_800_026, w_800_027, w_800_028, w_800_029, w_800_030, w_800_031, w_800_032, w_800_033, w_800_034, w_800_035, w_800_036, w_800_037, w_800_038, w_800_039, w_800_040, w_800_041, w_800_042, w_800_043, w_800_044, w_800_045, w_800_046, w_800_047, w_800_048, w_800_049, w_800_050, w_800_051, w_800_052, w_800_053, w_800_054, w_800_055, w_800_056, w_800_057, w_800_058, w_800_059, w_800_060, w_800_061, w_800_062, w_800_063, w_800_064, w_800_065, w_800_066, w_800_067, w_800_068, w_800_069, w_800_070, w_800_071, w_800_072, w_800_073, w_800_074, w_800_075, w_800_076, w_800_077, w_800_078, w_800_079, w_800_080, w_800_081, w_800_082, w_800_083, w_800_084, w_800_085, w_800_086, w_800_087, w_800_088, w_800_089, w_800_090, w_800_091, w_800_092, w_800_093, w_800_094, w_800_095, w_800_096, w_800_097, w_800_098, w_800_099, w_800_100, w_800_101, w_800_102, w_800_103, w_800_104, w_800_105, w_800_106, w_800_107, w_800_108, w_800_109, w_800_110, w_800_111, w_800_112, w_800_113, w_800_114, w_800_115, w_800_116, w_800_117, w_800_118, w_800_119, w_800_120, w_800_121, w_800_122, w_800_123, w_800_124, w_800_125, w_800_126, w_800_127, w_800_128, w_800_129, w_800_130, w_800_131, w_800_132, w_800_133, w_800_134, w_800_135, w_800_136, w_800_137, w_800_138, w_800_139, w_800_140, w_800_141, w_800_142, w_800_143, w_800_144, w_800_145, w_800_146, w_800_147, w_800_148, w_800_149, w_800_150, w_800_151, w_800_152, w_800_153, w_800_154, w_800_155, w_800_156, w_800_157, w_800_158, w_800_159, w_800_160, w_800_161, w_800_162, w_800_163, w_800_164, w_800_165, w_800_166, w_800_167, w_800_168, w_800_169, w_800_170, w_800_171, w_800_172, w_800_173, w_800_174, w_800_175, w_800_176, w_800_177, w_800_178, w_800_179, w_800_180, w_800_181, w_800_182, w_800_183, w_800_184, w_800_185, w_800_186, w_800_187, w_800_188, w_800_189, w_800_190, w_800_191, w_800_192, w_800_193, w_800_194, w_800_195, w_800_196, w_800_197, w_800_198, w_800_199, w_800_200, w_800_201, w_800_202, w_800_203, w_800_204, w_800_205, w_800_206, w_800_207, w_800_208, w_800_209, w_800_210, w_800_211, w_800_212, w_800_213, w_800_214, w_800_215, w_800_216, w_800_217, w_800_218, w_800_219, w_800_220, w_800_221, w_800_222, w_800_223, w_800_224, w_800_225, w_800_226, w_800_227, w_800_228, w_800_229, w_800_230, w_800_231, w_800_232, w_800_233, w_800_234, w_800_235, w_800_236, w_800_237, w_800_238, w_800_239, w_800_240, w_800_241, w_800_242, w_800_243, w_800_244, w_800_245, w_800_246, w_800_247, w_800_248, w_800_249, w_800_250, w_800_251, w_800_252, w_800_253, w_800_254, w_800_255, w_800_256, w_800_257, w_800_258, w_800_259, w_800_260, w_800_261, w_800_262, w_800_263, w_800_264, w_800_265, w_800_266, w_800_267, w_800_268, w_800_269, w_800_270, w_800_271, w_800_272, w_800_273, w_800_274, w_800_275, w_800_276, w_800_277, w_800_278, w_800_279, w_800_280, w_800_281, w_800_282, w_800_283, w_800_284, w_800_285, w_800_286, w_800_287, w_800_288, w_800_289, w_800_290, w_800_291, w_800_292, w_800_293, w_800_294, w_800_295, w_800_296, w_800_297, w_800_298, w_800_299, w_800_300, w_800_301, w_800_302, w_800_303, w_800_304, w_800_305, w_800_306, w_800_307, w_800_308, w_800_309, w_800_310, w_800_311, w_800_312, w_800_313, w_800_314, w_800_315, w_800_316, w_800_317, w_800_318, w_800_319, w_800_320, w_800_321, w_800_322, w_800_323, w_800_324, w_800_325, w_800_326, w_800_327, w_800_328, w_800_329, w_800_330, w_800_331, w_800_332, w_800_333, w_800_334, w_800_335, w_800_336, w_800_337, w_800_338, w_800_339, w_800_340, w_800_341, w_800_342, w_800_343, w_800_344, w_800_345, w_800_346, w_800_347, w_800_348, w_800_349, w_800_350, w_800_351, w_800_352, w_800_353, w_800_354, w_800_355, w_800_356, w_800_357, w_800_358, w_800_359, w_800_360, w_800_361, w_800_362, w_800_363, w_800_364, w_800_365, w_800_366, w_800_367, w_800_368, w_800_369, w_800_370, w_800_371, w_800_372, w_800_373, w_800_374, w_800_375, w_800_376, w_800_377, w_800_378, w_800_379, w_800_380, w_800_381, w_800_382, w_800_383, w_800_384, w_800_385, w_800_386, w_800_387, w_800_388, w_800_389, w_800_390, w_800_391, w_800_392, w_800_393, w_800_394, w_800_395, w_800_396, w_800_397, w_800_398, w_800_399, w_800_400, w_800_401, w_800_402, w_800_403, w_800_404, w_800_405, w_800_406, w_800_407, w_800_408, w_800_409, w_800_410, w_800_411, w_800_412, w_800_413, w_800_414, w_800_415, w_800_416, w_800_417, w_800_418, w_800_419, w_800_420, w_800_421, w_800_422, w_800_423, w_800_424, w_800_425, w_800_426, w_800_427, w_800_428, w_800_429, w_800_430, w_800_431, w_800_432, w_800_433, w_800_434, w_800_435, w_800_436, w_800_437, w_800_438, w_800_439, w_800_440, w_800_441, w_800_442, w_800_443, w_800_444, w_800_445, w_800_446, w_800_447, w_800_448, w_800_449, w_800_450, w_800_451, w_800_452, w_800_453, w_800_454, w_800_455, w_800_456, w_800_457, w_800_458, w_800_459, w_800_460, w_800_461, w_800_462, w_800_463, w_800_464, w_800_465, w_800_466, w_800_467, w_800_468, w_800_469, w_800_470, w_800_471, w_800_472, w_800_473, w_800_474, w_800_475, w_800_476, w_800_477, w_800_478, w_800_479, w_800_480, w_800_481, w_800_482, w_800_483, w_800_484, w_800_485, w_800_486, w_800_487, w_800_488, w_800_489, w_800_490, w_800_491, w_800_492, w_800_493, w_800_494, w_800_495, w_800_496, w_800_497, w_800_498, w_800_499, w_800_500, w_800_501, w_800_502, w_800_503, w_800_504, w_800_505, w_800_506, w_800_507, w_800_508, w_800_509, w_800_510, w_800_511, w_800_512, w_800_513, w_800_514, w_800_515, w_800_516, w_800_517, w_800_518, w_800_519, w_800_520, w_800_521, w_800_522, w_800_523, w_800_524, w_800_525, w_800_526, w_800_527, w_800_528, w_800_529, w_800_530, w_800_531, w_800_532, w_800_533, w_800_534, w_800_535, w_800_536, w_800_537, w_800_538, w_800_539, w_800_540, w_800_541, w_800_542, w_800_543, w_800_544, w_800_545, w_800_546, w_800_547, w_800_548, w_800_549, w_800_550, w_800_551, w_800_552, w_800_553, w_800_554, w_800_555, w_800_556, w_800_557, w_800_558, w_800_559, w_800_560, w_800_561, w_800_562, w_800_563, w_800_564, w_800_565, w_800_566, w_800_567, w_800_568, w_800_569, w_800_570, w_800_571, w_800_572, w_800_573, w_800_574, w_800_575, w_800_576, w_800_577, w_800_578, w_800_579, w_800_580, w_800_581, w_800_582, w_800_583, w_800_584, w_800_585, w_800_586, w_800_587, w_800_588, w_800_589, w_800_590, w_800_591, w_800_592, w_800_593, w_800_594, w_800_595, w_800_596, w_800_597, w_800_598, w_800_599, w_800_600, w_800_601, w_800_602, w_800_603, w_800_604, w_800_605, w_800_606, w_800_607, w_800_608, w_800_609, w_800_610, w_800_611, w_800_612, w_800_613, w_800_614, w_800_615, w_800_616, w_800_617, w_800_618, w_800_619, w_800_620, w_800_621, w_800_622, w_800_623, w_800_624, w_800_625, w_800_626, w_800_627, w_800_628, w_800_629, w_800_630, w_800_631, w_800_632, w_800_633, w_800_634, w_800_635, w_800_636, w_800_637, w_800_638, w_800_639, w_800_640, w_800_641, w_800_642, w_800_643, w_800_644, w_800_645, w_800_646, w_800_647, w_800_648, w_800_649, w_800_650, w_800_651, w_800_652, w_800_653, w_800_654, w_800_655, w_800_656, w_800_657, w_800_658, w_800_659, w_800_660, w_800_661, w_800_662, w_800_663, w_800_664, w_800_665, w_800_666, w_800_667, w_800_668, w_800_669, w_800_670, w_800_671, w_800_672, w_800_673, w_800_674, w_800_675, w_800_676, w_800_677, w_800_678, w_800_679, w_800_680, w_800_681, w_800_682, w_800_683, w_800_684, w_800_685, w_800_686, w_800_687, w_800_688, w_800_689, w_800_690, w_800_691, w_800_692, w_800_693, w_800_694, w_800_695, w_800_696, w_800_697, w_800_698, w_800_699, w_800_700, w_800_701, w_800_702, w_800_703, w_800_704, w_800_705, w_800_706, w_800_707, w_800_708, w_800_709, w_800_710, w_800_711, w_800_712, w_800_713, w_800_714, w_800_715, w_800_716, w_800_717);
    #100;
    $finish;
  end
  always #1 r0 = ~r0;
  always #2 r1 = ~r1;
  always #4 r2 = ~r2;
  always #8 r3 = ~r3;
  always #16 r4 = ~r4;
  always #32 r5 = ~r5;
  always #64 r6 = ~r6;
  always #128 r7 = ~r7;
  always #256 r8 = ~r8;
  always #512 r9 = ~r9;
  always #1024 r10 = ~r10;
  always #2048 r11 = ~r11;
  always #4096 r12 = ~r12;
  always #8192 r13 = ~r13;
  always #16384 r14 = ~r14;
  always #32768 r15 = ~r15;
  always #65536 r16 = ~r16;
  always #131072 r17 = ~r17;
  always #262144 r18 = ~r18;
  always #524288 r19 = ~r19;
  always #1048576 r20 = ~r20;
  always #2097152 r21 = ~r21;
  always #4194304 r22 = ~r22;
  always #8388608 r23 = ~r23;
  always #16777216 r24 = ~r24;
  always #33554432 r25 = ~r25;
  always #67108864 r26 = ~r26;
  always #134217728 r27 = ~r27;
  always #268435456 r28 = ~r28;
  always #536870912 r29 = ~r29;
  always #1073741824 r30 = ~r30;
  always #2147483648 r31 = ~r31;
  always #4294967296 r32 = ~r32;
  always #8589934592 r33 = ~r33;
  always #17179869184 r34 = ~r34;
  always #34359738368 r35 = ~r35;
  always #68719476736 r36 = ~r36;
  always #137438953472 r37 = ~r37;
  always #274877906944 r38 = ~r38;
  always #549755813888 r39 = ~r39;
  always #1099511627776 r40 = ~r40;
  always #2199023255552 r41 = ~r41;
  always #4398046511104 r42 = ~r42;
  always #8796093022208 r43 = ~r43;
  always #17592186044416 r44 = ~r44;
  always #35184372088832 r45 = ~r45;
  always #70368744177664 r46 = ~r46;
  always #140737488355328 r47 = ~r47;
  always #281474976710656 r48 = ~r48;
  always #562949953421312 r49 = ~r49;
  always #1125899906842624 r50 = ~r50;
  always #2251799813685248 r51 = ~r51;
  always #4503599627370496 r52 = ~r52;
  always #9007199254740992 r53 = ~r53;
  always #18014398509481984 r54 = ~r54;
  always #36028797018963968 r55 = ~r55;
  always #72057594037927936 r56 = ~r56;
  always #144115188075855872 r57 = ~r57;
  always #288230376151711744 r58 = ~r58;
  always #576460752303423488 r59 = ~r59;
  always #1152921504606846976 r60 = ~r60;
  always #2305843009213693952 r61 = ~r61;
  always #4611686018427387904 r62 = ~r62;
  always #9223372036854775808 r63 = ~r63;
  always #1 r64 = ~r64;
  always #2 r65 = ~r65;
  always #4 r66 = ~r66;
  always #8 r67 = ~r67;
  always #16 r68 = ~r68;
  always #32 r69 = ~r69;
  always #64 r70 = ~r70;
  always #128 r71 = ~r71;
  always #256 r72 = ~r72;
  always #512 r73 = ~r73;
  always #1024 r74 = ~r74;
  always #2048 r75 = ~r75;
  always #4096 r76 = ~r76;
  always #8192 r77 = ~r77;
  always #16384 r78 = ~r78;
  always #32768 r79 = ~r79;
  always #65536 r80 = ~r80;
  always #131072 r81 = ~r81;
  always #262144 r82 = ~r82;
  always #524288 r83 = ~r83;
  always #1048576 r84 = ~r84;
  always #2097152 r85 = ~r85;
  always #4194304 r86 = ~r86;
  always #8388608 r87 = ~r87;
  always #16777216 r88 = ~r88;
  always #33554432 r89 = ~r89;
  always #67108864 r90 = ~r90;
  always #134217728 r91 = ~r91;
  always #268435456 r92 = ~r92;
  always #536870912 r93 = ~r93;
  always #1073741824 r94 = ~r94;
  always #2147483648 r95 = ~r95;
  always #4294967296 r96 = ~r96;
  always #8589934592 r97 = ~r97;
  always #17179869184 r98 = ~r98;
  always #34359738368 r99 = ~r99;
  always #68719476736 r100 = ~r100;
  always #137438953472 r101 = ~r101;
  always #274877906944 r102 = ~r102;
  always #549755813888 r103 = ~r103;
  always #1099511627776 r104 = ~r104;
  always #2199023255552 r105 = ~r105;
  always #4398046511104 r106 = ~r106;
  always #8796093022208 r107 = ~r107;
  always #17592186044416 r108 = ~r108;
  always #35184372088832 r109 = ~r109;
  always #70368744177664 r110 = ~r110;
  always #140737488355328 r111 = ~r111;
  always #281474976710656 r112 = ~r112;
  always #562949953421312 r113 = ~r113;
  always #1125899906842624 r114 = ~r114;
  always #2251799813685248 r115 = ~r115;
  always #4503599627370496 r116 = ~r116;
  always #9007199254740992 r117 = ~r117;
  always #18014398509481984 r118 = ~r118;
  always #36028797018963968 r119 = ~r119;
  always #72057594037927936 r120 = ~r120;
  always #144115188075855872 r121 = ~r121;
  always #288230376151711744 r122 = ~r122;
  always #576460752303423488 r123 = ~r123;
  always #1152921504606846976 r124 = ~r124;
  always #2305843009213693952 r125 = ~r125;
  always #4611686018427387904 r126 = ~r126;
  always #9223372036854775808 r127 = ~r127;
  always #1 r128 = ~r128;
  always #2 r129 = ~r129;
  always #4 r130 = ~r130;
  always #8 r131 = ~r131;
  always #16 r132 = ~r132;
  always #32 r133 = ~r133;
  always #64 r134 = ~r134;
  always #128 r135 = ~r135;
  always #256 r136 = ~r136;
  always #512 r137 = ~r137;
  always #1024 r138 = ~r138;
  always #2048 r139 = ~r139;
  always #4096 r140 = ~r140;
  always #8192 r141 = ~r141;
  always #16384 r142 = ~r142;
  always #32768 r143 = ~r143;
  always #65536 r144 = ~r144;
  always #131072 r145 = ~r145;
  always #262144 r146 = ~r146;
  always #524288 r147 = ~r147;
  always #1048576 r148 = ~r148;
  always #2097152 r149 = ~r149;
  always #4194304 r150 = ~r150;
  always #8388608 r151 = ~r151;
  always #16777216 r152 = ~r152;
  always #33554432 r153 = ~r153;
  always #67108864 r154 = ~r154;
  always #134217728 r155 = ~r155;
  always #268435456 r156 = ~r156;
  always #536870912 r157 = ~r157;
  always #1073741824 r158 = ~r158;
  always #2147483648 r159 = ~r159;
  always #4294967296 r160 = ~r160;
  always #8589934592 r161 = ~r161;
  always #17179869184 r162 = ~r162;
  always #34359738368 r163 = ~r163;
  always #68719476736 r164 = ~r164;
  always #137438953472 r165 = ~r165;
  always #274877906944 r166 = ~r166;
  always #549755813888 r167 = ~r167;
  always #1099511627776 r168 = ~r168;
  always #2199023255552 r169 = ~r169;
  always #4398046511104 r170 = ~r170;
  always #8796093022208 r171 = ~r171;
  always #17592186044416 r172 = ~r172;
  always #35184372088832 r173 = ~r173;
  always #70368744177664 r174 = ~r174;
  always #140737488355328 r175 = ~r175;
  always #281474976710656 r176 = ~r176;
  always #562949953421312 r177 = ~r177;
  always #1125899906842624 r178 = ~r178;
  always #2251799813685248 r179 = ~r179;
  always #4503599627370496 r180 = ~r180;
  always #9007199254740992 r181 = ~r181;
  always #18014398509481984 r182 = ~r182;
  always #36028797018963968 r183 = ~r183;
  always #72057594037927936 r184 = ~r184;
  always #144115188075855872 r185 = ~r185;
  always #288230376151711744 r186 = ~r186;
  always #576460752303423488 r187 = ~r187;
  always #1152921504606846976 r188 = ~r188;
  always #2305843009213693952 r189 = ~r189;
  always #4611686018427387904 r190 = ~r190;
  always #9223372036854775808 r191 = ~r191;
  always #1 r192 = ~r192;
  always #2 r193 = ~r193;
  always #4 r194 = ~r194;
  always #8 r195 = ~r195;
  always #16 r196 = ~r196;
  always #32 r197 = ~r197;
  always #64 r198 = ~r198;
  always #128 r199 = ~r199;
  always #256 r200 = ~r200;
  always #512 r201 = ~r201;
  always #1024 r202 = ~r202;
  always #2048 r203 = ~r203;
  always #4096 r204 = ~r204;
  always #8192 r205 = ~r205;
  always #16384 r206 = ~r206;
  always #32768 r207 = ~r207;
  always #65536 r208 = ~r208;
  always #131072 r209 = ~r209;
  always #262144 r210 = ~r210;
  always #524288 r211 = ~r211;
  always #1048576 r212 = ~r212;
  always #2097152 r213 = ~r213;
  always #4194304 r214 = ~r214;
  always #8388608 r215 = ~r215;
  always #16777216 r216 = ~r216;
  always #33554432 r217 = ~r217;
  always #67108864 r218 = ~r218;
  always #134217728 r219 = ~r219;
  always #268435456 r220 = ~r220;
  always #536870912 r221 = ~r221;
  always #1073741824 r222 = ~r222;
  always #2147483648 r223 = ~r223;
  always #4294967296 r224 = ~r224;
  always #8589934592 r225 = ~r225;
  always #17179869184 r226 = ~r226;
  always #34359738368 r227 = ~r227;
  always #68719476736 r228 = ~r228;
  always #137438953472 r229 = ~r229;
  always #274877906944 r230 = ~r230;
  always #549755813888 r231 = ~r231;
  always #1099511627776 r232 = ~r232;
  always #2199023255552 r233 = ~r233;
  always #4398046511104 r234 = ~r234;
  always #8796093022208 r235 = ~r235;
  always #17592186044416 r236 = ~r236;
  always #35184372088832 r237 = ~r237;
  always #70368744177664 r238 = ~r238;
  always #140737488355328 r239 = ~r239;
  always #281474976710656 r240 = ~r240;
  always #562949953421312 r241 = ~r241;
  always #1125899906842624 r242 = ~r242;
  always #2251799813685248 r243 = ~r243;
  always #4503599627370496 r244 = ~r244;
  always #9007199254740992 r245 = ~r245;
  always #18014398509481984 r246 = ~r246;
  always #36028797018963968 r247 = ~r247;
  always #72057594037927936 r248 = ~r248;
  always #144115188075855872 r249 = ~r249;
  always #288230376151711744 r250 = ~r250;
  always #576460752303423488 r251 = ~r251;
  always #1152921504606846976 r252 = ~r252;
  always #2305843009213693952 r253 = ~r253;
  always #4611686018427387904 r254 = ~r254;
  always #9223372036854775808 r255 = ~r255;
  always #1 r256 = ~r256;
  always #2 r257 = ~r257;
  always #4 r258 = ~r258;
  always #8 r259 = ~r259;
  always #16 r260 = ~r260;
  always #32 r261 = ~r261;
  always #64 r262 = ~r262;
  always #128 r263 = ~r263;
  always #256 r264 = ~r264;
  always #512 r265 = ~r265;
  always #1024 r266 = ~r266;
  always #2048 r267 = ~r267;
  always #4096 r268 = ~r268;
  always #8192 r269 = ~r269;
  always #16384 r270 = ~r270;
  always #32768 r271 = ~r271;
  always #65536 r272 = ~r272;
  always #131072 r273 = ~r273;
  always #262144 r274 = ~r274;
  always #524288 r275 = ~r275;
  always #1048576 r276 = ~r276;
  always #2097152 r277 = ~r277;
  always #4194304 r278 = ~r278;
  always #8388608 r279 = ~r279;
  always #16777216 r280 = ~r280;
  always #33554432 r281 = ~r281;
  always #67108864 r282 = ~r282;
  always #134217728 r283 = ~r283;
  always #268435456 r284 = ~r284;
  always #536870912 r285 = ~r285;
  always #1073741824 r286 = ~r286;
  always #2147483648 r287 = ~r287;
  always #4294967296 r288 = ~r288;
  always #8589934592 r289 = ~r289;
  always #17179869184 r290 = ~r290;
  always #34359738368 r291 = ~r291;
  always #68719476736 r292 = ~r292;
  always #137438953472 r293 = ~r293;
  always #274877906944 r294 = ~r294;
  always #549755813888 r295 = ~r295;
  always #1099511627776 r296 = ~r296;
  always #2199023255552 r297 = ~r297;
  always #4398046511104 r298 = ~r298;
  always #8796093022208 r299 = ~r299;
  always #17592186044416 r300 = ~r300;
  always #35184372088832 r301 = ~r301;
  always #70368744177664 r302 = ~r302;
  always #140737488355328 r303 = ~r303;
  always #281474976710656 r304 = ~r304;
  always #562949953421312 r305 = ~r305;
  always #1125899906842624 r306 = ~r306;
  always #2251799813685248 r307 = ~r307;
  always #4503599627370496 r308 = ~r308;
  always #9007199254740992 r309 = ~r309;
  always #18014398509481984 r310 = ~r310;
  always #36028797018963968 r311 = ~r311;
  always #72057594037927936 r312 = ~r312;
  always #144115188075855872 r313 = ~r313;
  always #288230376151711744 r314 = ~r314;
  always #576460752303423488 r315 = ~r315;
  always #1152921504606846976 r316 = ~r316;
  always #2305843009213693952 r317 = ~r317;
  always #4611686018427387904 r318 = ~r318;
  always #9223372036854775808 r319 = ~r319;
  always #1 r320 = ~r320;
  always #2 r321 = ~r321;
  always #4 r322 = ~r322;
  always #8 r323 = ~r323;
  always #16 r324 = ~r324;
  always #32 r325 = ~r325;
  always #64 r326 = ~r326;
  always #128 r327 = ~r327;
  always #256 r328 = ~r328;
  always #512 r329 = ~r329;
  always #1024 r330 = ~r330;
  always #2048 r331 = ~r331;
  always #4096 r332 = ~r332;
  always #8192 r333 = ~r333;
  always #16384 r334 = ~r334;
  always #32768 r335 = ~r335;
  always #65536 r336 = ~r336;
  always #131072 r337 = ~r337;
  always #262144 r338 = ~r338;
  always #524288 r339 = ~r339;
  always #1048576 r340 = ~r340;
  always #2097152 r341 = ~r341;
  always #4194304 r342 = ~r342;
  always #8388608 r343 = ~r343;
  always #16777216 r344 = ~r344;
  always #33554432 r345 = ~r345;
  always #67108864 r346 = ~r346;
  always #134217728 r347 = ~r347;
  always #268435456 r348 = ~r348;
  always #536870912 r349 = ~r349;
  always #1073741824 r350 = ~r350;
  always #2147483648 r351 = ~r351;
  always #4294967296 r352 = ~r352;
  always #8589934592 r353 = ~r353;
  always #17179869184 r354 = ~r354;
  always #34359738368 r355 = ~r355;
  always #68719476736 r356 = ~r356;
  always #137438953472 r357 = ~r357;
  always #274877906944 r358 = ~r358;
  always #549755813888 r359 = ~r359;
  always #1099511627776 r360 = ~r360;
  always #2199023255552 r361 = ~r361;
  always #4398046511104 r362 = ~r362;
  always #8796093022208 r363 = ~r363;
  always #17592186044416 r364 = ~r364;
  always #35184372088832 r365 = ~r365;
  always #70368744177664 r366 = ~r366;
  always #140737488355328 r367 = ~r367;
  always #281474976710656 r368 = ~r368;
  always #562949953421312 r369 = ~r369;
  always #1125899906842624 r370 = ~r370;
  always #2251799813685248 r371 = ~r371;
  always #4503599627370496 r372 = ~r372;
  always #9007199254740992 r373 = ~r373;
  always #18014398509481984 r374 = ~r374;
  always #36028797018963968 r375 = ~r375;
  always #72057594037927936 r376 = ~r376;
  always #144115188075855872 r377 = ~r377;
  always #288230376151711744 r378 = ~r378;
  always #576460752303423488 r379 = ~r379;
  always #1152921504606846976 r380 = ~r380;
  always #2305843009213693952 r381 = ~r381;
  always #4611686018427387904 r382 = ~r382;
  always #9223372036854775808 r383 = ~r383;
  always #1 r384 = ~r384;
  always #2 r385 = ~r385;
  always #4 r386 = ~r386;
  always #8 r387 = ~r387;
  always #16 r388 = ~r388;
  always #32 r389 = ~r389;
  always #64 r390 = ~r390;
  always #128 r391 = ~r391;
  always #256 r392 = ~r392;
  always #512 r393 = ~r393;
  always #1024 r394 = ~r394;
  always #2048 r395 = ~r395;
  always #4096 r396 = ~r396;
  always #8192 r397 = ~r397;
  always #16384 r398 = ~r398;
  always #32768 r399 = ~r399;
  always #65536 r400 = ~r400;
  always #131072 r401 = ~r401;
  always #262144 r402 = ~r402;
  always #524288 r403 = ~r403;
  always #1048576 r404 = ~r404;
  always #2097152 r405 = ~r405;
  always #4194304 r406 = ~r406;
  always #8388608 r407 = ~r407;
  always #16777216 r408 = ~r408;
  always #33554432 r409 = ~r409;
  always #67108864 r410 = ~r410;
  always #134217728 r411 = ~r411;
  always #268435456 r412 = ~r412;
  always #536870912 r413 = ~r413;
  always #1073741824 r414 = ~r414;
  always #2147483648 r415 = ~r415;
  always #4294967296 r416 = ~r416;
  always #8589934592 r417 = ~r417;
  always #17179869184 r418 = ~r418;
  always #34359738368 r419 = ~r419;
  always #68719476736 r420 = ~r420;
  always #137438953472 r421 = ~r421;
  always #274877906944 r422 = ~r422;
  always #549755813888 r423 = ~r423;
  always #1099511627776 r424 = ~r424;
  always #2199023255552 r425 = ~r425;
  always #4398046511104 r426 = ~r426;
  always #8796093022208 r427 = ~r427;
  always #17592186044416 r428 = ~r428;
  always #35184372088832 r429 = ~r429;
  always #70368744177664 r430 = ~r430;
  always #140737488355328 r431 = ~r431;
  always #281474976710656 r432 = ~r432;
  always #562949953421312 r433 = ~r433;
  always #1125899906842624 r434 = ~r434;
  always #2251799813685248 r435 = ~r435;
  always #4503599627370496 r436 = ~r436;
  always #9007199254740992 r437 = ~r437;
  always #18014398509481984 r438 = ~r438;
  always #36028797018963968 r439 = ~r439;
  always #72057594037927936 r440 = ~r440;
  always #144115188075855872 r441 = ~r441;
  always #288230376151711744 r442 = ~r442;
  always #576460752303423488 r443 = ~r443;
  always #1152921504606846976 r444 = ~r444;
  always #2305843009213693952 r445 = ~r445;
  always #4611686018427387904 r446 = ~r446;
  always #9223372036854775808 r447 = ~r447;
  always #1 r448 = ~r448;
  always #2 r449 = ~r449;
  always #4 r450 = ~r450;
  always #8 r451 = ~r451;
  always #16 r452 = ~r452;
  always #32 r453 = ~r453;
  always #64 r454 = ~r454;
  always #128 r455 = ~r455;
  always #256 r456 = ~r456;
  always #512 r457 = ~r457;
  always #1024 r458 = ~r458;
  always #2048 r459 = ~r459;
  always #4096 r460 = ~r460;
  always #8192 r461 = ~r461;
  always #16384 r462 = ~r462;
  always #32768 r463 = ~r463;
  always #65536 r464 = ~r464;
  always #131072 r465 = ~r465;
  always #262144 r466 = ~r466;
  always #524288 r467 = ~r467;
  always #1048576 r468 = ~r468;
  always #2097152 r469 = ~r469;
  always #4194304 r470 = ~r470;
  always #8388608 r471 = ~r471;
  always #16777216 r472 = ~r472;
  always #33554432 r473 = ~r473;
  always #67108864 r474 = ~r474;
  always #134217728 r475 = ~r475;
  always #268435456 r476 = ~r476;
  always #536870912 r477 = ~r477;
  always #1073741824 r478 = ~r478;
  always #2147483648 r479 = ~r479;
  always #4294967296 r480 = ~r480;
  always #8589934592 r481 = ~r481;
  always #17179869184 r482 = ~r482;
  always #34359738368 r483 = ~r483;
  always #68719476736 r484 = ~r484;
  always #137438953472 r485 = ~r485;
  always #274877906944 r486 = ~r486;
  always #549755813888 r487 = ~r487;
  always #1099511627776 r488 = ~r488;
  always #2199023255552 r489 = ~r489;
  always #4398046511104 r490 = ~r490;
  always #8796093022208 r491 = ~r491;
  always #17592186044416 r492 = ~r492;
  always #35184372088832 r493 = ~r493;
  always #70368744177664 r494 = ~r494;
  always #140737488355328 r495 = ~r495;
  always #281474976710656 r496 = ~r496;
  always #562949953421312 r497 = ~r497;
  always #1125899906842624 r498 = ~r498;
  always #2251799813685248 r499 = ~r499;
  always #4503599627370496 r500 = ~r500;
  always #9007199254740992 r501 = ~r501;
  always #18014398509481984 r502 = ~r502;
  always #36028797018963968 r503 = ~r503;
  always #72057594037927936 r504 = ~r504;
  always #144115188075855872 r505 = ~r505;
  always #288230376151711744 r506 = ~r506;
  always #576460752303423488 r507 = ~r507;
  always #1152921504606846976 r508 = ~r508;
  always #2305843009213693952 r509 = ~r509;
  always #4611686018427387904 r510 = ~r510;
  always #9223372036854775808 r511 = ~r511;
  always #1 r512 = ~r512;
  always #2 r513 = ~r513;
  always #4 r514 = ~r514;
  always #8 r515 = ~r515;
  always #16 r516 = ~r516;
  always #32 r517 = ~r517;
  always #64 r518 = ~r518;
  always #128 r519 = ~r519;
  always #256 r520 = ~r520;
  always #512 r521 = ~r521;
  always #1024 r522 = ~r522;
  always #2048 r523 = ~r523;
  always #4096 r524 = ~r524;
  always #8192 r525 = ~r525;
  always #16384 r526 = ~r526;
  always #32768 r527 = ~r527;
  always #65536 r528 = ~r528;
  always #131072 r529 = ~r529;
  always #262144 r530 = ~r530;
  always #524288 r531 = ~r531;
  always #1048576 r532 = ~r532;
  always #2097152 r533 = ~r533;
  always #4194304 r534 = ~r534;
  always #8388608 r535 = ~r535;
  always #16777216 r536 = ~r536;
  always #33554432 r537 = ~r537;
  always #67108864 r538 = ~r538;
  always #134217728 r539 = ~r539;
  always #268435456 r540 = ~r540;
  always #536870912 r541 = ~r541;
  always #1073741824 r542 = ~r542;
  always #2147483648 r543 = ~r543;
  always #4294967296 r544 = ~r544;
  always #8589934592 r545 = ~r545;
  always #17179869184 r546 = ~r546;
  always #34359738368 r547 = ~r547;
  always #68719476736 r548 = ~r548;
  always #137438953472 r549 = ~r549;
  always #274877906944 r550 = ~r550;
  always #549755813888 r551 = ~r551;
  always #1099511627776 r552 = ~r552;
  always #2199023255552 r553 = ~r553;
  always #4398046511104 r554 = ~r554;
  always #8796093022208 r555 = ~r555;
  always #17592186044416 r556 = ~r556;
  always #35184372088832 r557 = ~r557;
  always #70368744177664 r558 = ~r558;
  always #140737488355328 r559 = ~r559;
  always #281474976710656 r560 = ~r560;
  always #562949953421312 r561 = ~r561;
  always #1125899906842624 r562 = ~r562;
  always #2251799813685248 r563 = ~r563;
  always #4503599627370496 r564 = ~r564;
  always #9007199254740992 r565 = ~r565;
  always #18014398509481984 r566 = ~r566;
  always #36028797018963968 r567 = ~r567;
  always #72057594037927936 r568 = ~r568;
  always #144115188075855872 r569 = ~r569;
  always #288230376151711744 r570 = ~r570;
  always #576460752303423488 r571 = ~r571;
  always #1152921504606846976 r572 = ~r572;
  always #2305843009213693952 r573 = ~r573;
  always #4611686018427387904 r574 = ~r574;
  always #9223372036854775808 r575 = ~r575;
  always #1 r576 = ~r576;
  always #2 r577 = ~r577;
  always #4 r578 = ~r578;
  always #8 r579 = ~r579;
  always #16 r580 = ~r580;
  always #32 r581 = ~r581;
  always #64 r582 = ~r582;
  always #128 r583 = ~r583;
  always #256 r584 = ~r584;
  always #512 r585 = ~r585;
  always #1024 r586 = ~r586;
  always #2048 r587 = ~r587;
  always #4096 r588 = ~r588;
  always #8192 r589 = ~r589;
  always #16384 r590 = ~r590;
  always #32768 r591 = ~r591;
  always #65536 r592 = ~r592;
  always #131072 r593 = ~r593;
  always #262144 r594 = ~r594;
  always #524288 r595 = ~r595;
  always #1048576 r596 = ~r596;
  always #2097152 r597 = ~r597;
  always #4194304 r598 = ~r598;
  always #8388608 r599 = ~r599;
  always #16777216 r600 = ~r600;
  always #33554432 r601 = ~r601;
  always #67108864 r602 = ~r602;
  always #134217728 r603 = ~r603;
  always #268435456 r604 = ~r604;
  always #536870912 r605 = ~r605;
  always #1073741824 r606 = ~r606;
  always #2147483648 r607 = ~r607;
  always #4294967296 r608 = ~r608;
  always #8589934592 r609 = ~r609;
  always #17179869184 r610 = ~r610;
  always #34359738368 r611 = ~r611;
  always #68719476736 r612 = ~r612;
  always #137438953472 r613 = ~r613;
  always #274877906944 r614 = ~r614;
  always #549755813888 r615 = ~r615;
  always #1099511627776 r616 = ~r616;
  always #2199023255552 r617 = ~r617;
  always #4398046511104 r618 = ~r618;
  always #8796093022208 r619 = ~r619;
  always #17592186044416 r620 = ~r620;
  always #35184372088832 r621 = ~r621;
  always #70368744177664 r622 = ~r622;
  always #140737488355328 r623 = ~r623;
  always #281474976710656 r624 = ~r624;
  always #562949953421312 r625 = ~r625;
  always #1125899906842624 r626 = ~r626;
  always #2251799813685248 r627 = ~r627;
  always #4503599627370496 r628 = ~r628;
  always #9007199254740992 r629 = ~r629;
  always #18014398509481984 r630 = ~r630;
  always #36028797018963968 r631 = ~r631;
  always #72057594037927936 r632 = ~r632;
  always #144115188075855872 r633 = ~r633;
  always #288230376151711744 r634 = ~r634;
  always #576460752303423488 r635 = ~r635;
  always #1152921504606846976 r636 = ~r636;
  always #2305843009213693952 r637 = ~r637;
  always #4611686018427387904 r638 = ~r638;
  always #9223372036854775808 r639 = ~r639;
  always #1 r640 = ~r640;
  always #2 r641 = ~r641;
  always #4 r642 = ~r642;
  always #8 r643 = ~r643;
  always #16 r644 = ~r644;
  always #32 r645 = ~r645;
  always #64 r646 = ~r646;
  always #128 r647 = ~r647;
  always #256 r648 = ~r648;
  always #512 r649 = ~r649;
  always #1024 r650 = ~r650;
  always #2048 r651 = ~r651;
  always #4096 r652 = ~r652;
  always #8192 r653 = ~r653;
  always #16384 r654 = ~r654;
  always #32768 r655 = ~r655;
  always #65536 r656 = ~r656;
  always #131072 r657 = ~r657;
  always #262144 r658 = ~r658;
  always #524288 r659 = ~r659;
  always #1048576 r660 = ~r660;
  always #2097152 r661 = ~r661;
  always #4194304 r662 = ~r662;
  always #8388608 r663 = ~r663;
  always #16777216 r664 = ~r664;
  always #33554432 r665 = ~r665;
  always #67108864 r666 = ~r666;
  always #134217728 r667 = ~r667;
  always #268435456 r668 = ~r668;
  always #536870912 r669 = ~r669;
  always #1073741824 r670 = ~r670;
  always #2147483648 r671 = ~r671;
  always #4294967296 r672 = ~r672;
  always #8589934592 r673 = ~r673;
  always #17179869184 r674 = ~r674;
  always #34359738368 r675 = ~r675;
  always #68719476736 r676 = ~r676;
  always #137438953472 r677 = ~r677;
  always #274877906944 r678 = ~r678;
  always #549755813888 r679 = ~r679;
  always #1099511627776 r680 = ~r680;
  always #2199023255552 r681 = ~r681;
  always #4398046511104 r682 = ~r682;
  always #8796093022208 r683 = ~r683;
  always #17592186044416 r684 = ~r684;
  always #35184372088832 r685 = ~r685;
  always #70368744177664 r686 = ~r686;
  always #140737488355328 r687 = ~r687;
  always #281474976710656 r688 = ~r688;
  always #562949953421312 r689 = ~r689;
  always #1125899906842624 r690 = ~r690;
  always #2251799813685248 r691 = ~r691;
  always #4503599627370496 r692 = ~r692;
  always #9007199254740992 r693 = ~r693;
  always #18014398509481984 r694 = ~r694;
  always #36028797018963968 r695 = ~r695;
  always #72057594037927936 r696 = ~r696;
  always #144115188075855872 r697 = ~r697;
  always #288230376151711744 r698 = ~r698;
  always #576460752303423488 r699 = ~r699;
  always #1152921504606846976 r700 = ~r700;
  always #2305843009213693952 r701 = ~r701;
  always #4611686018427387904 r702 = ~r702;
  always #9223372036854775808 r703 = ~r703;
  always #1 r704 = ~r704;
  always #2 r705 = ~r705;
  always #4 r706 = ~r706;
  always #8 r707 = ~r707;
  always #16 r708 = ~r708;
  always #32 r709 = ~r709;
  always #64 r710 = ~r710;
  always #128 r711 = ~r711;
  always #256 r712 = ~r712;
  always #512 r713 = ~r713;
  always #1024 r714 = ~r714;
  always #2048 r715 = ~r715;
  always #4096 r716 = ~r716;
  always #8192 r717 = ~r717;
  always #16384 r718 = ~r718;
  always #32768 r719 = ~r719;
  always #65536 r720 = ~r720;
  always #131072 r721 = ~r721;
  always #262144 r722 = ~r722;
  always #524288 r723 = ~r723;
  always #1048576 r724 = ~r724;
  always #2097152 r725 = ~r725;
  always #4194304 r726 = ~r726;
  always #8388608 r727 = ~r727;
  always #16777216 r728 = ~r728;
  always #33554432 r729 = ~r729;
  always #67108864 r730 = ~r730;
  always #134217728 r731 = ~r731;
  always #268435456 r732 = ~r732;
  always #536870912 r733 = ~r733;
  always #1073741824 r734 = ~r734;
  always #2147483648 r735 = ~r735;
  always #4294967296 r736 = ~r736;
  always #8589934592 r737 = ~r737;
  always #17179869184 r738 = ~r738;
  always #34359738368 r739 = ~r739;
  always #68719476736 r740 = ~r740;
  always #137438953472 r741 = ~r741;
  always #274877906944 r742 = ~r742;
  always #549755813888 r743 = ~r743;
  always #1099511627776 r744 = ~r744;
  always #2199023255552 r745 = ~r745;
  always #4398046511104 r746 = ~r746;
  always #8796093022208 r747 = ~r747;
  always #17592186044416 r748 = ~r748;
  always #35184372088832 r749 = ~r749;
  always #70368744177664 r750 = ~r750;
  always #140737488355328 r751 = ~r751;
  always #281474976710656 r752 = ~r752;
  always #562949953421312 r753 = ~r753;
  always #1125899906842624 r754 = ~r754;
  always #2251799813685248 r755 = ~r755;
  always #4503599627370496 r756 = ~r756;
  always #9007199254740992 r757 = ~r757;
  always #18014398509481984 r758 = ~r758;
  always #36028797018963968 r759 = ~r759;
  always #72057594037927936 r760 = ~r760;
  always #144115188075855872 r761 = ~r761;
  always #288230376151711744 r762 = ~r762;
  always #576460752303423488 r763 = ~r763;
  always #1152921504606846976 r764 = ~r764;
  always #2305843009213693952 r765 = ~r765;
  always #4611686018427387904 r766 = ~r766;
  always #9223372036854775808 r767 = ~r767;
  always #1 r768 = ~r768;
  always #2 r769 = ~r769;
  always #4 r770 = ~r770;
  always #8 r771 = ~r771;
  always #16 r772 = ~r772;
  always #32 r773 = ~r773;
  always #64 r774 = ~r774;
  always #128 r775 = ~r775;
  always #256 r776 = ~r776;
  always #512 r777 = ~r777;
  always #1024 r778 = ~r778;
  always #2048 r779 = ~r779;
  always #4096 r780 = ~r780;
  always #8192 r781 = ~r781;
  always #16384 r782 = ~r782;
  always #32768 r783 = ~r783;
  always #65536 r784 = ~r784;
  always #131072 r785 = ~r785;
  always #262144 r786 = ~r786;
  always #524288 r787 = ~r787;
  always #1048576 r788 = ~r788;
  always #2097152 r789 = ~r789;
  always #4194304 r790 = ~r790;
  always #8388608 r791 = ~r791;
  always #16777216 r792 = ~r792;
  always #33554432 r793 = ~r793;
  always #67108864 r794 = ~r794;
  always #134217728 r795 = ~r795;
  always #268435456 r796 = ~r796;
  always #536870912 r797 = ~r797;
endmodule
*/
// ****** TestBench Module Defination End ******


// Gate Level Verilog Code Generated!
// GateLvl:30 GateNum:30 GateInputNum:2
// ****** Basic Gate Module Defination ******
module or2(out, in1, in2);
  output out;
  input in1, in2;
  wire in1, in2, out;
  assign out = in1 || in2;
endmodule

module and2(out, in1, in2);
  output out;
  input in1, in2;
  wire in1, in2, out;
  assign out = in1 && in2;
endmodule

module not1(out, in);
  output out;
  input in;
  wire in,out;
  assign out = ~in;
endmodule

module nand2(out, in1, in2);
  output out;
  input in1, in2;
  wire in1, in2, out;
  assign out = ~(in1 && in2);
endmodule
// ****** Basic Gate Module Defination End ******

// ****** Combined Logic Module Defination ******
module combLogic( w_000_000, w_000_001, w_000_002, w_000_003, w_000_004, w_000_005, w_000_006, w_000_007, w_000_008, w_000_009, w_000_010, w_000_011, w_000_012, w_000_013, w_000_014, w_000_015, w_000_016, w_000_017, w_000_018, w_000_019, w_000_021, w_000_022, w_000_024, w_000_025, w_000_029, w_030_000 );
  inout w_000_000, w_000_001, w_000_002, w_000_003, w_000_004, w_000_005, w_000_006, w_000_007, w_000_008, w_000_009, w_000_010, w_000_011, w_000_012, w_000_013, w_000_014, w_000_015, w_000_016, w_000_017, w_000_018, w_000_019, w_000_021, w_000_022, w_000_024, w_000_025, w_000_029;
  output w_030_000;
  wire w_000_000, w_000_001, w_000_002, w_000_003, w_000_004, w_000_005, w_000_006, w_000_007, w_000_008, w_000_009, w_000_010, w_000_011, w_000_012, w_000_013, w_000_014, w_000_015, w_000_016, w_000_017, w_000_018, w_000_019, w_000_021, w_000_022, w_000_024, w_000_025, w_000_029;
  wire w_001_000, w_001_001, w_001_002, w_001_003, w_001_004, w_001_005, w_001_006, w_001_007, w_001_008, w_001_009;
  wire w_002_000, w_002_001, w_002_002, w_002_003, w_002_004, w_002_005, w_002_006, w_002_007, w_002_008, w_002_009, w_002_011, w_002_012, w_002_013;
  wire w_003_003, w_003_004, w_003_005, w_003_007, w_003_008, w_003_010, w_003_011, w_003_012, w_003_013, w_003_014, w_003_017, w_003_019, w_003_020;
  wire w_004_000, w_004_001, w_004_002, w_004_004, w_004_008, w_004_011, w_004_012, w_004_013, w_004_015, w_004_016, w_004_018, w_004_019, w_004_020, w_004_021;
  wire w_005_002, w_005_004, w_005_007, w_005_008, w_005_010, w_005_011, w_005_013, w_005_014;
  wire w_006_002, w_006_004, w_006_013, w_006_019, w_006_021, w_006_022, w_006_024;
  wire w_007_005, w_007_008, w_007_009, w_007_010, w_007_012, w_007_015;
  wire w_008_000, w_008_001, w_008_002;
  wire w_009_000, w_009_001;
  wire w_010_000, w_010_002, w_010_003, w_010_006, w_010_008, w_010_015, w_010_022, w_010_025, w_010_026;
  wire w_011_001, w_011_002, w_011_003, w_011_004, w_011_005, w_011_006, w_011_007;
  wire w_012_003, w_012_006, w_012_022, w_012_029, w_012_030, w_012_031, w_012_032, w_012_033, w_012_034, w_012_035, w_012_036, w_012_037, w_012_039, w_012_041, w_012_042, w_012_043, w_012_044, w_012_045, w_012_046, w_012_047, w_012_048, w_012_049, w_012_050, w_012_051, w_012_053;
  wire w_013_000, w_013_002, w_013_004, w_013_005;
  wire w_014_000, w_014_001, w_014_003, w_014_005, w_014_006, w_014_007;
  wire w_015_000, w_015_007, w_015_011, w_015_017, w_015_021;
  wire w_016_023, w_016_028, w_016_029, w_016_030;
  wire w_018_031, w_018_032, w_018_033, w_018_034, w_018_035, w_018_036, w_018_037, w_018_038, w_018_039, w_018_043, w_018_044, w_018_045, w_018_046, w_018_047, w_018_048, w_018_049, w_018_051;
  wire w_019_003, w_019_012, w_019_019;
  wire w_020_007, w_020_021;
  wire w_021_000;
  wire w_022_030, w_022_031, w_022_032, w_022_033, w_022_034, w_022_035, w_022_036, w_022_040, w_022_041, w_022_042, w_022_043, w_022_044, w_022_045, w_022_046, w_022_047, w_022_048, w_022_049, w_022_050, w_022_051, w_022_053;
  wire w_023_000;
  wire w_024_010, w_024_011, w_024_012, w_024_013, w_024_014, w_024_015, w_024_016, w_024_017, w_024_018, w_024_019, w_024_020, w_024_024, w_024_025, w_024_026, w_024_027, w_024_028, w_024_029, w_024_030, w_024_031, w_024_032, w_024_033, w_024_035;
  wire w_030_000;
  not1 I001_000(w_001_000, w_000_000);
  nand2 I001_001(w_001_001, w_000_001, w_000_002);
  not1 I001_002(w_001_002, w_000_003);
  or2  I001_003(w_001_003, w_000_001, w_000_002);
  nand2 I001_004(w_001_004, w_000_004, w_000_005);
  nand2 I001_005(w_001_005, w_000_006, w_000_000);
  not1 I001_006(w_001_006, w_000_007);
  and2 I001_007(w_001_007, w_000_008, w_000_009);
  or2  I001_008(w_001_008, w_000_002, w_000_010);
  not1 I001_009(w_001_009, w_000_011);
  nand2 I002_000(w_002_000, w_001_002, w_000_012);
  or2  I002_001(w_002_001, w_001_003, w_000_001);
  not1 I002_002(w_002_002, w_001_003);
  or2  I002_003(w_002_003, w_001_004, w_001_008);
  and2 I002_004(w_002_004, w_001_000, w_001_006);
  nand2 I002_005(w_002_005, w_000_013, w_001_002);
  not1 I002_006(w_002_006, w_000_001);
  or2  I002_007(w_002_007, w_001_004, w_001_006);
  or2  I002_008(w_002_008, w_000_009, w_001_007);
  and2 I002_009(w_002_009, w_001_002, w_001_004);
  nand2 I002_011(w_002_011, w_000_006, w_000_008);
  and2 I002_012(w_002_012, w_001_001, w_000_015);
  and2 I002_013(w_002_013, w_000_016, w_000_017);
  and2 I003_003(w_003_003, w_001_006, w_001_000);
  not1 I003_004(w_003_004, w_001_005);
  or2  I003_005(w_003_005, w_001_009, w_000_007);
  nand2 I003_007(w_003_007, w_000_016, w_002_003);
  not1 I003_008(w_003_008, w_002_002);
  and2 I003_010(w_003_010, w_002_003, w_002_000);
  and2 I003_011(w_003_011, w_001_005, w_001_009);
  and2 I003_012(w_003_012, w_002_008, w_001_006);
  nand2 I003_013(w_003_013, w_001_005, w_002_000);
  and2 I003_014(w_003_014, w_002_001, w_002_013);
  or2  I003_017(w_003_017, w_000_016, w_001_001);
  nand2 I003_018(w_003_020, w_001_008, w_003_019);
  and2 I003_019(w_003_019, w_003_020, w_002_002);
  and2 I004_000(w_004_000, w_003_017, w_002_001);
  not1 I004_001(w_004_001, w_003_011);
  or2  I004_002(w_004_002, w_003_013, w_002_008);
  and2 I004_004(w_004_004, w_003_013, w_001_008);
  nand2 I004_008(w_004_008, w_002_009, w_002_001);
  not1 I004_011(w_004_011, w_000_007);
  nand2 I004_012(w_004_012, w_003_004, w_000_011);
  not1 I004_013(w_004_013, w_000_019);
  nand2 I004_015(w_004_015, w_002_001, w_001_001);
  not1 I004_016(w_004_016, w_002_005);
  or2  I004_018(w_004_018, w_000_016, w_002_008);
  and2 I004_019(w_004_019, w_001_002, w_000_000);
  and2 I004_020(w_004_020, w_000_021, w_003_010);
  and2 I004_021(w_004_021, w_003_003, w_002_013);
  not1 I005_002(w_005_002, w_001_003);
  or2  I005_004(w_005_004, w_004_019, w_001_000);
  or2  I005_007(w_005_007, w_001_001, w_000_014);
  and2 I005_008(w_005_008, w_002_002, w_000_022);
  not1 I005_010(w_005_010, w_003_008);
  not1 I005_011(w_005_011, w_004_020);
  nand2 I005_013(w_005_013, w_004_004, w_004_001);
  or2  I005_014(w_005_014, w_001_000, w_000_010);
  and2 I006_002(w_006_002, w_001_002, w_000_018);
  and2 I006_004(w_006_004, w_000_013, w_002_003);
  and2 I006_013(w_006_013, w_004_002, w_002_013);
  nand2 I006_019(w_006_019, w_003_010, w_004_011);
  nand2 I006_021(w_006_021, w_005_007, w_003_010);
  not1 I006_022(w_006_022, w_002_007);
  and2 I006_024(w_006_024, w_003_003, w_005_004);
  and2 I007_005(w_007_005, w_005_002, w_000_010);
  not1 I007_008(w_007_008, w_001_002);
  not1 I007_009(w_007_009, w_002_009);
  not1 I007_010(w_007_010, w_000_009);
  and2 I007_012(w_007_012, w_002_013, w_004_000);
  or2  I007_015(w_007_015, w_000_019, w_004_018);
  nand2 I008_000(w_008_000, w_001_008, w_001_007);
  or2  I008_001(w_008_001, w_003_007, w_006_002);
  not1 I008_002(w_008_002, w_007_009);
  nand2 I009_000(w_009_000, w_005_011, w_002_004);
  not1 I009_001(w_009_001, w_002_007);
  or2  I010_000(w_010_000, w_008_001, w_009_001);
  or2  I010_002(w_010_002, w_007_005, w_002_012);
  not1 I010_003(w_010_003, w_002_001);
  or2  I010_006(w_010_006, w_000_024, w_000_008);
  nand2 I010_008(w_010_008, w_009_000, w_004_008);
  or2  I010_015(w_010_015, w_004_021, w_005_014);
  nand2 I010_022(w_010_022, w_007_012, w_005_008);
  nand2 I010_025(w_010_025, w_003_005, w_003_008);
  or2  I010_026(w_010_026, w_001_000, w_008_001);
  and2 I011_001(w_011_001, w_002_007, w_004_015);
  or2  I011_002(w_011_002, w_006_024, w_009_001);
  not1 I011_003(w_011_003, w_003_005);
  or2  I011_004(w_011_004, w_004_015, w_004_019);
  and2 I011_005(w_011_005, w_010_026, w_009_001);
  and2 I011_006(w_011_006, w_000_025, w_002_012);
  nand2 I011_007(w_011_007, w_004_018, w_004_012);
  not1 I012_003(w_012_003, w_006_013);
  and2 I012_006(w_012_006, w_010_003, w_002_006);
  or2  I012_022(w_012_022, w_002_011, w_001_003);
  nand2 I012_028(w_012_030, w_012_029, w_009_000);
  nand2 I012_029(w_012_031, w_009_000, w_012_030);
  not1 I012_030(w_012_032, w_012_031);
  or2  I012_031(w_012_033, w_004_002, w_012_032);
  nand2 I012_032(w_012_034, w_012_033, w_003_012);
  not1 I012_033(w_012_035, w_012_034);
  and2 I012_034(w_012_036, w_003_003, w_012_035);
  nand2 I012_035(w_012_037, w_012_036, w_012_053);
  not1 I012_036(w_012_029, w_012_037);
  nand2 I012_037(w_012_042, w_005_008, w_012_041);
  and2 I012_038(w_012_043, w_011_001, w_012_042);
  not1 I012_039(w_012_044, w_012_043);
  not1 I012_040(w_012_045, w_012_044);
  or2  I012_041(w_012_046, w_012_045, w_011_005);
  and2 I012_042(w_012_047, w_004_016, w_012_046);
  nand2 I012_043(w_012_048, w_012_047, w_003_014);
  and2 I012_044(w_012_049, w_012_048, w_008_002);
  not1 I012_045(w_012_050, w_012_049);
  not1 I012_046(w_012_051, w_012_050);
  not1 I012_047(w_012_041, w_012_037);
  and2 I012_048(w_012_053, w_010_006, w_012_051);
  not1 I013_000(w_013_000, w_005_002);
  nand2 I013_002(w_013_002, w_009_000, w_010_025);
  not1 I013_004(w_013_004, w_005_007);
  and2 I013_005(w_013_005, w_007_010, w_007_015);
  and2 I013_009(w_012_039, w_002_002, w_012_029);
  and2 I014_000(w_014_000, w_013_005, w_010_000);
  or2  I014_001(w_014_001, w_012_039, w_009_000);
  nand2 I014_003(w_014_003, w_001_009, w_000_018);
  or2  I014_005(w_014_005, w_012_006, w_013_004);
  nand2 I014_006(w_014_006, w_005_010, w_012_022);
  or2  I014_007(w_014_007, w_001_005, w_010_008);
  or2  I015_000(w_015_000, w_010_022, w_009_001);
  not1 I015_007(w_015_007, w_008_000);
  nand2 I015_011(w_015_011, w_005_010, w_011_002);
  or2  I015_017(w_015_017, w_001_000, w_011_004);
  or2  I015_021(w_015_021, w_000_029, w_014_001);
  or2  I016_023(w_016_023, w_014_003, w_015_007);
  not1 I016_027(w_016_029, w_016_028);
  not1 I016_028(w_016_030, w_016_029);
  nand2 I016_029(w_016_028, w_015_011, w_016_030);
  and2 I018_030(w_018_032, w_018_031, w_011_007);
  and2 I018_031(w_018_033, w_015_021, w_018_032);
  not1 I018_032(w_018_034, w_018_033);
  and2 I018_033(w_018_035, w_018_034, w_001_009);
  nand2 I018_034(w_018_036, w_010_002, w_018_035);
  not1 I018_035(w_018_037, w_018_036);
  not1 I018_036(w_018_038, w_018_037);
  not1 I018_037(w_018_039, w_018_038);
  and2 I018_038(w_018_031, w_018_051, w_018_039);
  or2  I018_039(w_018_044, w_014_007, w_018_043);
  or2  I018_040(w_018_045, w_018_044, w_011_006);
  and2 I018_041(w_018_046, w_018_045, w_011_003);
  or2  I018_042(w_018_047, w_011_001, w_018_046);
  nand2 I018_043(w_018_048, w_013_004, w_018_047);
  not1 I018_044(w_018_049, w_018_048);
  not1 I018_045(w_018_043, w_018_031);
  and2 I018_046(w_018_051, w_008_002, w_018_049);
  and2 I019_003(w_019_003, w_009_000, w_014_005);
  and2 I019_012(w_019_012, w_009_001, w_013_000);
  or2  I019_019(w_019_019, w_014_000, w_007_008);
  nand2 I020_007(w_020_007, w_014_006, w_008_002);
  not1 I020_021(w_020_021, w_002_004);
  nand2 I021_000(w_021_000, w_006_021, w_008_001);
  nand2 I022_029(w_022_031, w_004_011, w_022_030);
  or2  I022_030(w_022_032, w_022_031, w_022_053);
  and2 I022_031(w_022_033, w_022_032, w_005_013);
  nand2 I022_032(w_022_034, w_019_012, w_022_033);
  or2  I022_033(w_022_035, w_013_002, w_022_034);
  and2 I022_034(w_022_036, w_022_035, w_014_001);
  not1 I022_035(w_022_030, w_022_036);
  nand2 I022_036(w_022_041, w_022_040, w_004_013);
  or2  I022_037(w_022_042, w_022_041, w_015_017);
  and2 I022_038(w_022_043, w_001_005, w_022_042);
  not1 I022_039(w_022_044, w_022_043);
  nand2 I022_040(w_022_045, w_005_013, w_022_044);
  and2 I022_041(w_022_046, w_022_045, w_018_037);
  nand2 I022_042(w_022_047, w_022_046, w_011_002);
  or2  I022_043(w_022_048, w_022_047, w_020_021);
  not1 I022_044(w_022_049, w_022_048);
  not1 I022_045(w_022_050, w_022_049);
  or2  I022_046(w_022_051, w_006_022, w_022_050);
  not1 I022_047(w_022_040, w_022_032);
  and2 I022_048(w_022_053, w_015_000, w_022_051);
  nand2 I023_000(w_023_000, w_009_000, w_000_022);
  or2  I024_009(w_024_011, w_024_010, w_006_019);
  and2 I024_010(w_024_012, w_010_015, w_024_011);
  or2  I024_011(w_024_013, w_024_035, w_024_012);
  and2 I024_012(w_024_014, w_024_013, w_007_015);
  nand2 I024_013(w_024_015, w_024_014, w_012_003);
  or2  I024_014(w_024_016, w_024_015, w_002_002);
  not1 I024_015(w_024_017, w_024_016);
  or2  I024_016(w_024_018, w_024_017, w_005_007);
  not1 I024_017(w_024_019, w_024_018);
  not1 I024_018(w_024_020, w_024_019);
  or2  I024_019(w_024_010, w_024_020, w_019_019);
  and2 I024_020(w_024_025, w_006_004, w_024_024);
  not1 I024_021(w_024_026, w_024_025);
  or2  I024_022(w_024_027, w_024_026, w_021_000);
  nand2 I024_023(w_024_028, w_024_027, w_011_006);
  and2 I024_024(w_024_029, w_024_028, w_023_000);
  not1 I024_025(w_024_030, w_024_029);
  or2  I024_026(w_024_031, w_014_006, w_024_030);
  and2 I024_027(w_024_032, w_020_007, w_024_031);
  or2  I024_028(w_024_033, w_024_032, w_008_001);
  not1 I024_029(w_024_024, w_024_013);
  and2 I024_030(w_024_035, w_011_007, w_024_033);
  and2 I030_000(w_030_000, w_019_003, w_016_023);

  initial begin
    $get_module_info();
  end
endmodule

// ****** Combined Logic Module Defination ******

// ****** TestBench Module Defination ******

/*
module tb();
  wire  w_000_000, w_000_001, w_000_002, w_000_003, w_000_004, w_000_005, w_000_006, w_000_007, w_000_008, w_000_009, w_000_010, w_000_011, w_000_012, w_000_013, w_000_014, w_000_015, w_000_016, w_000_017, w_000_018, w_000_019, w_000_021, w_000_022, w_000_024, w_000_025, w_000_029, w_030_000 ;
  combLogic I0(  w_000_000, w_000_001, w_000_002, w_000_003, w_000_004, w_000_005, w_000_006, w_000_007, w_000_008, w_000_009, w_000_010, w_000_011, w_000_012, w_000_013, w_000_014, w_000_015, w_000_016, w_000_017, w_000_018, w_000_019, w_000_021, w_000_022, w_000_024, w_000_025, w_000_029, w_030_000  );

  reg r0, r1, r2, r3, r4, r5, r6, r7, r8, r9, r10, r11, r12, r13, r14, r15, r16, r17, r18, r19, r20, r21, r22, r23, r24, r25, r26, r27, r28, r29, rEnd; 

  assign w_000_000 = r0;
  assign w_000_001 = r1;
  assign w_000_002 = r2;
  assign w_000_003 = r3;
  assign w_000_004 = r4;
  assign w_000_005 = r5;
  assign w_000_006 = r6;
  assign w_000_007 = r7;
  assign w_000_008 = r8;
  assign w_000_009 = r9;
  assign w_000_010 = r10;
  assign w_000_011 = r11;
  assign w_000_012 = r12;
  assign w_000_013 = r13;
  assign w_000_014 = r14;
  assign w_000_015 = r15;
  assign w_000_016 = r16;
  assign w_000_017 = r17;
  assign w_000_018 = r18;
  assign w_000_019 = r19;
  assign w_000_020 = r20;
  assign w_000_021 = r21;
  assign w_000_022 = r22;
  assign w_000_023 = r23;
  assign w_000_024 = r24;
  assign w_000_025 = r25;
  assign w_000_026 = r26;
  assign w_000_027 = r27;
  assign w_000_028 = r28;
  assign w_000_029 = r29;

  initial begin 
    r0 = 1'b0; 
    r1 = 1'b0; 
    r2 = 1'b0; 
    r3 = 1'b0; 
    r4 = 1'b0; 
    r5 = 1'b0; 
    r6 = 1'b0; 
    r7 = 1'b0; 
    r8 = 1'b0; 
    r9 = 1'b0; 
    r10 = 1'b0; 
    r11 = 1'b0; 
    r12 = 1'b0; 
    r13 = 1'b0; 
    r14 = 1'b0; 
    r15 = 1'b0; 
    r16 = 1'b0; 
    r17 = 1'b0; 
    r18 = 1'b0; 
    r19 = 1'b0; 
    r20 = 1'b0; 
    r21 = 1'b0; 
    r22 = 1'b0; 
    r23 = 1'b0; 
    r24 = 1'b0; 
    r25 = 1'b0; 
    r26 = 1'b0; 
    r27 = 1'b0; 
    r28 = 1'b0; 
    r29 = 1'b0; 
    $monitor("%t %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b  ", $time, w_000_000, w_000_001, w_000_002, w_000_003, w_000_004, w_000_005, w_000_006, w_000_007, w_000_008, w_000_009, w_000_010, w_000_011, w_000_012, w_000_013, w_000_014, w_000_015, w_000_016, w_000_017, w_000_018, w_000_019, w_000_020, w_000_021, w_000_022, w_000_023, w_000_024, w_000_025, w_000_026, w_000_027, w_000_028, w_000_029, w_030_000);
    #100;
    $finish;
  end
  always #1 r0 = ~r0;
  always #2 r1 = ~r1;
  always #4 r2 = ~r2;
  always #8 r3 = ~r3;
  always #16 r4 = ~r4;
  always #32 r5 = ~r5;
  always #64 r6 = ~r6;
  always #128 r7 = ~r7;
  always #256 r8 = ~r8;
  always #512 r9 = ~r9;
  always #1024 r10 = ~r10;
  always #2048 r11 = ~r11;
  always #4096 r12 = ~r12;
  always #8192 r13 = ~r13;
  always #16384 r14 = ~r14;
  always #32768 r15 = ~r15;
  always #65536 r16 = ~r16;
  always #131072 r17 = ~r17;
  always #262144 r18 = ~r18;
  always #524288 r19 = ~r19;
  always #1048576 r20 = ~r20;
  always #2097152 r21 = ~r21;
  always #4194304 r22 = ~r22;
  always #8388608 r23 = ~r23;
  always #16777216 r24 = ~r24;
  always #33554432 r25 = ~r25;
  always #67108864 r26 = ~r26;
  always #134217728 r27 = ~r27;
  always #268435456 r28 = ~r28;
  always #536870912 r29 = ~r29;
endmodule
*/
// ****** TestBench Module Defination End ******

/*
// ******* The results for this case *********
******* result_1.txt *********
1)
  Loop Signals: w_018_031, w_018_032, w_018_033, w_018_034, w_018_035, w_018_036, w_018_037, w_018_038, w_018_039, 
  Loop Gates: I018_030.port1, I018_031.port2, I018_032.port1, I018_033.port1, I018_034.port2, I018_035.port1, I018_036.port1, I018_037.port1, I018_038.port2, 

2)
  Loop Signals: w_018_031, w_018_043, w_018_044, w_018_045, w_018_046, w_018_047, w_018_048, w_018_049, w_018_051, 
  Loop Gates: I018_038.port1, I018_039.port2, I018_040.port1, I018_041.port1, I018_042.port2, I018_043.port2, I018_044.port1, I018_045.port1, I018_046.port2, 

3)
  Loop Signals: w_016_028, w_016_029, w_016_030, 
  Loop Gates: I016_027.port1, I016_028.port1, I016_029.port2, 

4)
  Loop Signals: w_022_030, w_022_031, w_022_032, w_022_033, w_022_034, w_022_035, w_022_036, 
  Loop Gates: I022_029.port2, I022_030.port1, I022_031.port1, I022_032.port2, I022_033.port2, I022_034.port1, I022_035.port1, 

5)
  Loop Signals: w_022_032, w_022_040, w_022_041, w_022_042, w_022_043, w_022_044, w_022_045, w_022_046, w_022_047, w_022_048, w_022_049, w_022_050, w_022_051, w_022_053, 
  Loop Gates: I022_030.port2, I022_036.port1, I022_037.port1, I022_038.port2, I022_039.port1, I022_040.port2, I022_041.port1, I022_042.port1, I022_043.port1, I022_044.port1, I022_045.port1, I022_046.port2, I022_047.port1, I022_048.port2, 

6)
  Loop Signals: w_012_029, w_012_030, w_012_031, w_012_032, w_012_033, w_012_034, w_012_035, w_012_036, w_012_037, 
  Loop Gates: I012_028.port1, I012_029.port2, I012_030.port1, I012_031.port2, I012_032.port1, I012_033.port1, I012_034.port2, I012_035.port1, I012_036.port1, 

7)
  Loop Signals: w_012_037, w_012_041, w_012_042, w_012_043, w_012_044, w_012_045, w_012_046, w_012_047, w_012_048, w_012_049, w_012_050, w_012_051, w_012_053, 
  Loop Gates: I012_035.port2, I012_037.port2, I012_038.port2, I012_039.port1, I012_040.port1, I012_041.port1, I012_042.port2, I012_043.port1, I012_044.port1, I012_045.port1, I012_046.port1, I012_047.port1, I012_048.port2, 

8)
  Loop Signals: w_024_010, w_024_011, w_024_012, w_024_013, w_024_014, w_024_015, w_024_016, w_024_017, w_024_018, w_024_019, w_024_020, 
  Loop Gates: I024_009.port1, I024_010.port2, I024_011.port2, I024_012.port1, I024_013.port1, I024_014.port1, I024_015.port1, I024_016.port1, I024_017.port1, I024_018.port1, I024_019.port1, 

9)
  Loop Signals: w_024_013, w_024_024, w_024_025, w_024_026, w_024_027, w_024_028, w_024_029, w_024_030, w_024_031, w_024_032, w_024_033, w_024_035, 
  Loop Gates: I024_011.port1, I024_020.port2, I024_021.port1, I024_022.port1, I024_023.port1, I024_024.port1, I024_025.port1, I024_026.port2, I024_027.port2, I024_028.port1, I024_029.port1, I024_030.port2, 

10)
  Loop Signals: w_003_019, w_003_020, 
  Loop Gates: I003_018.port2, I003_019.port1, 

******* result_2.txt *********
1)
  Loop Signals: w_012_037, w_012_041, w_012_042, w_012_043, w_012_044, w_012_045, w_012_046, w_012_047, w_012_048, w_012_049, w_012_050, w_012_051, w_012_053, 
  Loop Gates: I012_035.port2, I012_037.port2, I012_038.port2, I012_039.port1, I012_040.port1, I012_041.port1, I012_042.port2, I012_043.port1, I012_044.port1, I012_045.port1, I012_046.port1, I012_047.port1, I012_048.port2, 

2)
  Loop Signals: w_024_010, w_024_011, w_024_012, w_024_013, w_024_014, w_024_015, w_024_016, w_024_017, w_024_018, w_024_019, w_024_020, 
  Loop Gates: I024_009.port1, I024_010.port2, I024_011.port2, I024_012.port1, I024_013.port1, I024_014.port1, I024_015.port1, I024_016.port1, I024_017.port1, I024_018.port1, I024_019.port1, 

3)
  Loop Signals: w_024_013, w_024_024, w_024_025, w_024_026, w_024_027, w_024_028, w_024_029, w_024_030, w_024_031, w_024_032, w_024_033, w_024_035, 
  Loop Gates: I024_011.port1, I024_020.port2, I024_021.port1, I024_022.port1, I024_023.port1, I024_024.port1, I024_025.port1, I024_026.port2, I024_027.port2, I024_028.port1, I024_029.port1, I024_030.port2, 

******* result_3.txt *********
1)
  Loop Signals: w_018_031, w_018_032, w_018_033, w_018_034, w_018_035, w_018_036, w_018_037, w_018_038, w_018_039, 
  Loop Gates: I018_030.port1, I018_031.port2, I018_032.port1, I018_033.port1, I018_034.port2, I018_035.port1, I018_036.port1, I018_037.port1, I018_038.port2, 
  Loop Conditions: I018_030.port2=1, I018_031.port1=1, I018_033.port2=1, I018_034.port1=1, I018_038.port2=1, 
  (Signal Values: w_001_009=1, w_010_002=1, w_011_007=1, w_015_021=1, w_018_039=1, )

2)
  Loop Signals: w_018_031, w_018_043, w_018_044, w_018_045, w_018_046, w_018_047, w_018_048, w_018_049, w_018_051, 
  Loop Gates: I018_038.port1, I018_039.port2, I018_040.port1, I018_041.port1, I018_042.port2, I018_043.port2, I018_044.port1, I018_045.port1, I018_046.port2, 
  Loop Conditions: I018_038.port2=1, I018_039.port1=0, I018_040.port2=0, I018_041.port2=1, I018_042.port1=0, I018_043.port1=1, I018_046.port2=1, 
  (Signal Values: w_011_003=1, w_011_001=0, w_011_006=0, w_013_004=1, w_014_007=0, w_018_039=1, w_018_049=1, )

3)
  Loop Signals: w_016_028, w_016_029, w_016_030, 
  Loop Gates: I016_027.port1, I016_028.port1, I016_029.port2, 
  Loop Conditions: I016_029.port1=1, 
  (Signal Values: w_015_011=1, )

4)
  Loop Signals: w_022_030, w_022_031, w_022_032, w_022_033, w_022_034, w_022_035, w_022_036, 
  Loop Gates: I022_029.port2, I022_030.port1, I022_031.port1, I022_032.port2, I022_033.port2, I022_034.port1, I022_035.port1, 
  Loop Conditions: I022_029.port1=1, I022_030.port2=0, I022_031.port2=1, I022_032.port1=1, I022_033.port1=0, I022_034.port2=1, 
  (Signal Values: w_004_011=1, w_005_013=1, w_013_002=0, w_014_001=1, w_019_012=1, w_022_053=0, )

5)
  Loop Signals: w_022_032, w_022_040, w_022_041, w_022_042, w_022_043, w_022_044, w_022_045, w_022_046, w_022_047, w_022_048, w_022_049, w_022_050, w_022_051, w_022_053, 
  Loop Gates: I022_030.port2, I022_036.port1, I022_037.port1, I022_038.port2, I022_039.port1, I022_040.port2, I022_041.port1, I022_042.port1, I022_043.port1, I022_044.port1, I022_045.port1, I022_046.port2, I022_047.port1, I022_048.port2, 
  Loop Conditions: I022_030.port2=0, I022_036.port2=1, I022_037.port2=0, I022_038.port1=1, I022_040.port1=1, I022_041.port2=1, I022_042.port2=1, I022_043.port2=0, I022_046.port1=0, I022_048.port2=1, 
  (Signal Values: w_001_005=1, w_004_013=1, w_005_013=1, w_006_022=0, w_011_002=1, w_015_017=0, w_018_037=1, w_020_021=0, w_022_051=1, w_022_053=0, )

6)
  Loop Signals: w_012_029, w_012_030, w_012_031, w_012_032, w_012_033, w_012_034, w_012_035, w_012_036, w_012_037, 
  Loop Gates: I012_028.port1, I012_029.port2, I012_030.port1, I012_031.port2, I012_032.port1, I012_033.port1, I012_034.port2, I012_035.port1, I012_036.port1, 
  Loop Conditions: I012_028.port2=1, I012_029.port1=1, I012_031.port1=0, I012_032.port2=1, I012_034.port1=1, I012_035.port2=1, 
  (Signal Values: w_003_003=1, w_003_012=1, w_004_002=0, w_009_000=1, w_012_053=1, )

7)
  Loop Signals: w_003_019, w_003_020, 
  Loop Gates: I003_018.port2, I003_019.port1, 
  Loop Conditions: I003_018.port1=1, I003_019.port2=1, 
  (Signal Values: w_001_008=1, w_002_002=1, )

******* result_4.txt *********
1)
  Loop Breaker: I018_038.port0-w_018_031-Register-w_018_031'-I018_030.port1 

2)
  Loop Breaker: I018_038.port0-w_018_031-Register-w_018_031'-I018_045.port1 

3)
  Loop Breaker: I016_027.port0-w_016_029-Register-w_016_029'-I016_028.port1 

4)
  Loop Breaker: I022_030.port0-w_022_032-Register-w_022_032'-I022_031.port1 

5)
  Loop Breaker: I022_030.port0-w_022_032-Register-w_022_032'-I022_047.port1 

6)
  Loop Breaker: I012_035.port0-w_012_037-Register-w_012_037'-I012_036.port1 

7)
  Loop Breaker: I003_018.port0-w_003_020-Register-w_003_020'-I003_019.port1 

// ******* The results for this case End *********
*/

// Gate Level Verilog Code Generated!
// GateLvl:2000 GateNum:2000 GateInputNum:2
// ****** Basic Gate Module Defination ******
module or2(out, in1, in2);
  output out;
  input in1, in2;
  wire in1, in2, out;
  assign out = in1 || in2;
endmodule

module and2(out, in1, in2);
  output out;
  input in1, in2;
  wire in1, in2, out;
  assign out = in1 && in2;
endmodule

module not1(out, in);
  output out;
  input in;
  wire in,out;
  assign out = ~in;
endmodule

module nand2(out, in1, in2);
  output out;
  input in1, in2;
  wire in1, in2, out;
  assign out = ~(in1 && in2);
endmodule
// ****** Basic Gate Module Defination End ******

// ****** Combined Logic Module Defination ******
module combLogic( w_000_000, w_000_001, w_000_002, w_000_003, w_000_004, w_000_005, w_000_006, w_000_007, w_000_008, w_000_009, w_000_010, w_000_011, w_000_012, w_000_013, w_000_014, w_000_015, w_000_016, w_000_017, w_000_018, w_000_019, w_000_020, w_000_021, w_000_022, w_000_023, w_000_024, w_000_025, w_000_026, w_000_027, w_000_028, w_000_029, w_000_030, w_000_031, w_000_032, w_000_033, w_000_034, w_000_035, w_000_036, w_000_037, w_000_038, w_000_039, w_000_040, w_000_041, w_000_042, w_000_043, w_000_044, w_000_045, w_000_046, w_000_047, w_000_048, w_000_049, w_000_050, w_000_051, w_000_052, w_000_053, w_000_054, w_000_055, w_000_056, w_000_057, w_000_058, w_000_059, w_000_060, w_000_061, w_000_062, w_000_063, w_000_065, w_000_066, w_000_067, w_000_068, w_000_069, w_000_070, w_000_071, w_000_072, w_000_073, w_000_074, w_000_075, w_000_076, w_000_077, w_000_078, w_000_079, w_000_080, w_000_081, w_000_082, w_000_083, w_000_084, w_000_085, w_000_086, w_000_087, w_000_088, w_000_089, w_000_090, w_000_091, w_000_092, w_000_093, w_000_094, w_000_095, w_000_096, w_000_097, w_000_098, w_000_099, w_000_100, w_000_101, w_000_102, w_000_103, w_000_104, w_000_105, w_000_106, w_000_107, w_000_108, w_000_109, w_000_110, w_000_111, w_000_112, w_000_113, w_000_114, w_000_115, w_000_116, w_000_117, w_000_118, w_000_119, w_000_120, w_000_121, w_000_122, w_000_123, w_000_124, w_000_125, w_000_126, w_000_127, w_000_128, w_000_129, w_000_130, w_000_131, w_000_132, w_000_133, w_000_134, w_000_135, w_000_136, w_000_137, w_000_138, w_000_139, w_000_140, w_000_141, w_000_142, w_000_143, w_000_144, w_000_145, w_000_146, w_000_147, w_000_148, w_000_149, w_000_150, w_000_151, w_000_152, w_000_153, w_000_154, w_000_155, w_000_156, w_000_157, w_000_158, w_000_159, w_000_160, w_000_161, w_000_162, w_000_163, w_000_164, w_000_165, w_000_166, w_000_167, w_000_168, w_000_169, w_000_170, w_000_171, w_000_172, w_000_173, w_000_174, w_000_175, w_000_176, w_000_177, w_000_178, w_000_179, w_000_180, w_000_181, w_000_182, w_000_183, w_000_184, w_000_185, w_000_186, w_000_187, w_000_188, w_000_189, w_000_190, w_000_191, w_000_192, w_000_193, w_000_194, w_000_195, w_000_196, w_000_197, w_000_198, w_000_199, w_000_200, w_000_201, w_000_202, w_000_203, w_000_204, w_000_205, w_000_206, w_000_207, w_000_208, w_000_209, w_000_210, w_000_211, w_000_212, w_000_213, w_000_214, w_000_215, w_000_216, w_000_217, w_000_218, w_000_219, w_000_220, w_000_221, w_000_222, w_000_223, w_000_224, w_000_225, w_000_226, w_000_227, w_000_228, w_000_229, w_000_230, w_000_231, w_000_232, w_000_233, w_000_234, w_000_235, w_000_236, w_000_237, w_000_238, w_000_239, w_000_240, w_000_241, w_000_242, w_000_243, w_000_244, w_000_245, w_000_246, w_000_247, w_000_248, w_000_249, w_000_250, w_000_251, w_000_252, w_000_253, w_000_254, w_000_255, w_000_256, w_000_257, w_000_258, w_000_259, w_000_260, w_000_261, w_000_262, w_000_263, w_000_264, w_000_265, w_000_266, w_000_267, w_000_268, w_000_269, w_000_270, w_000_271, w_000_272, w_000_273, w_000_274, w_000_275, w_000_276, w_000_277, w_000_278, w_000_279, w_000_280, w_000_281, w_000_282, w_000_283, w_000_284, w_000_285, w_000_286, w_000_287, w_000_289, w_000_290, w_000_291, w_000_292, w_000_293, w_000_294, w_000_295, w_000_296, w_000_297, w_000_298, w_000_299, w_000_300, w_000_301, w_000_302, w_000_303, w_000_304, w_000_305, w_000_306, w_000_307, w_000_308, w_000_309, w_000_310, w_000_311, w_000_312, w_000_313, w_000_314, w_000_315, w_000_316, w_000_317, w_000_318, w_000_319, w_000_320, w_000_321, w_000_322, w_000_323, w_000_324, w_000_325, w_000_326, w_000_327, w_000_328, w_000_329, w_000_330, w_000_331, w_000_332, w_000_333, w_000_334, w_000_335, w_000_336, w_000_337, w_000_338, w_000_339, w_000_340, w_000_341, w_000_342, w_000_343, w_000_344, w_000_345, w_000_346, w_000_347, w_000_348, w_000_349, w_000_350, w_000_351, w_000_352, w_000_353, w_000_354, w_000_355, w_000_356, w_000_357, w_000_358, w_000_359, w_000_360, w_000_361, w_000_362, w_000_363, w_000_364, w_000_365, w_000_366, w_000_367, w_000_368, w_000_369, w_000_370, w_000_371, w_000_372, w_000_373, w_000_374, w_000_375, w_000_376, w_000_377, w_000_378, w_000_379, w_000_380, w_000_381, w_000_382, w_000_383, w_000_384, w_000_385, w_000_386, w_000_387, w_000_388, w_000_389, w_000_390, w_000_391, w_000_392, w_000_393, w_000_394, w_000_395, w_000_396, w_000_397, w_000_398, w_000_399, w_000_400, w_000_401, w_000_402, w_000_403, w_000_404, w_000_405, w_000_406, w_000_407, w_000_408, w_000_409, w_000_410, w_000_411, w_000_412, w_000_413, w_000_414, w_000_415, w_000_416, w_000_417, w_000_418, w_000_419, w_000_420, w_000_421, w_000_422, w_000_423, w_000_424, w_000_425, w_000_426, w_000_427, w_000_428, w_000_429, w_000_430, w_000_431, w_000_432, w_000_433, w_000_434, w_000_435, w_000_436, w_000_437, w_000_438, w_000_439, w_000_440, w_000_441, w_000_442, w_000_443, w_000_444, w_000_445, w_000_446, w_000_447, w_000_448, w_000_449, w_000_450, w_000_451, w_000_452, w_000_453, w_000_454, w_000_455, w_000_456, w_000_457, w_000_458, w_000_459, w_000_460, w_000_461, w_000_462, w_000_463, w_000_464, w_000_465, w_000_466, w_000_467, w_000_468, w_000_469, w_000_470, w_000_471, w_000_472, w_000_473, w_000_474, w_000_475, w_000_476, w_000_477, w_000_478, w_000_479, w_000_480, w_000_481, w_000_482, w_000_483, w_000_484, w_000_485, w_000_486, w_000_487, w_000_488, w_000_489, w_000_490, w_000_491, w_000_492, w_000_493, w_000_494, w_000_495, w_000_496, w_000_498, w_000_499, w_000_500, w_000_501, w_000_502, w_000_503, w_000_504, w_000_505, w_000_506, w_000_507, w_000_508, w_000_509, w_000_510, w_000_511, w_000_512, w_000_513, w_000_514, w_000_515, w_000_516, w_000_517, w_000_518, w_000_519, w_000_520, w_000_521, w_000_522, w_000_523, w_000_524, w_000_525, w_000_526, w_000_527, w_000_528, w_000_529, w_000_530, w_000_531, w_000_532, w_000_533, w_000_534, w_000_535, w_000_536, w_000_537, w_000_538, w_000_539, w_000_540, w_000_541, w_000_542, w_000_543, w_000_544, w_000_545, w_000_546, w_000_547, w_000_548, w_000_549, w_000_550, w_000_551, w_000_552, w_000_553, w_000_554, w_000_555, w_000_556, w_000_557, w_000_558, w_000_559, w_000_560, w_000_561, w_000_562, w_000_563, w_000_564, w_000_565, w_000_566, w_000_567, w_000_568, w_000_569, w_000_570, w_000_571, w_000_572, w_000_573, w_000_575, w_000_576, w_000_577, w_000_578, w_000_579, w_000_580, w_000_581, w_000_582, w_000_583, w_000_584, w_000_585, w_000_586, w_000_587, w_000_588, w_000_589, w_000_590, w_000_591, w_000_592, w_000_593, w_000_594, w_000_595, w_000_596, w_000_597, w_000_598, w_000_599, w_000_600, w_000_601, w_000_602, w_000_603, w_000_604, w_000_605, w_000_606, w_000_607, w_000_608, w_000_609, w_000_610, w_000_611, w_000_612, w_000_613, w_000_614, w_000_615, w_000_616, w_000_617, w_000_618, w_000_619, w_000_620, w_000_621, w_000_622, w_000_623, w_000_624, w_000_625, w_000_626, w_000_627, w_000_628, w_000_629, w_000_630, w_000_631, w_000_632, w_000_633, w_000_634, w_000_635, w_000_636, w_000_638, w_000_639, w_000_640, w_000_641, w_000_643, w_000_644, w_000_645, w_000_646, w_000_647, w_000_648, w_000_649, w_000_650, w_000_651, w_000_652, w_000_653, w_000_654, w_000_655, w_000_656, w_000_657, w_000_658, w_000_659, w_000_660, w_000_661, w_000_662, w_000_663, w_000_664, w_000_665, w_000_667, w_000_668, w_000_669, w_000_670, w_000_671, w_000_672, w_000_673, w_000_674, w_000_675, w_000_676, w_000_677, w_000_678, w_000_679, w_000_680, w_000_681, w_000_682, w_000_683, w_000_684, w_000_685, w_000_686, w_000_687, w_000_688, w_000_689, w_000_690, w_000_691, w_000_692, w_000_693, w_000_694, w_000_695, w_000_696, w_000_697, w_000_698, w_000_699, w_000_700, w_000_701, w_000_702, w_000_703, w_000_704, w_000_705, w_000_706, w_000_707, w_000_708, w_000_709, w_000_710, w_000_711, w_000_712, w_000_713, w_000_714, w_000_715, w_000_716, w_000_717, w_000_718, w_000_719, w_000_720, w_000_721, w_000_722, w_000_723, w_000_724, w_000_725, w_000_726, w_000_727, w_000_728, w_000_729, w_000_730, w_000_731, w_000_732, w_000_733, w_000_734, w_000_735, w_000_736, w_000_737, w_000_738, w_000_739, w_000_740, w_000_741, w_000_742, w_000_743, w_000_744, w_000_745, w_000_746, w_000_747, w_000_748, w_000_749, w_000_750, w_000_751, w_000_752, w_000_753, w_000_754, w_000_755, w_000_756, w_000_757, w_000_758, w_000_759, w_000_760, w_000_761, w_000_762, w_000_763, w_000_764, w_000_765, w_000_766, w_000_767, w_000_768, w_000_769, w_000_770, w_000_771, w_000_772, w_000_773, w_000_774, w_000_775, w_000_776, w_000_777, w_000_778, w_000_779, w_000_780, w_000_781, w_000_782, w_000_783, w_000_784, w_000_785, w_000_786, w_000_787, w_000_788, w_000_789, w_000_790, w_000_791, w_000_792, w_000_793, w_000_794, w_000_795, w_000_796, w_000_797, w_000_798, w_000_799, w_000_800, w_000_801, w_000_802, w_000_803, w_000_804, w_000_805, w_000_806, w_000_807, w_000_808, w_000_809, w_000_810, w_000_811, w_000_812, w_000_813, w_000_814, w_000_815, w_000_816, w_000_817, w_000_818, w_000_819, w_000_820, w_000_821, w_000_822, w_000_823, w_000_824, w_000_825, w_000_826, w_000_827, w_000_828, w_000_829, w_000_830, w_000_831, w_000_832, w_000_833, w_000_835, w_000_836, w_000_837, w_000_838, w_000_839, w_000_840, w_000_841, w_000_842, w_000_843, w_000_844, w_000_845, w_000_846, w_000_847, w_000_848, w_000_849, w_000_850, w_000_851, w_000_852, w_000_853, w_000_854, w_000_855, w_000_856, w_000_857, w_000_858, w_000_859, w_000_860, w_000_861, w_000_862, w_000_863, w_000_864, w_000_865, w_000_866, w_000_867, w_000_868, w_000_869, w_000_870, w_000_871, w_000_872, w_000_873, w_000_874, w_000_875, w_000_876, w_000_877, w_000_878, w_000_879, w_000_880, w_000_881, w_000_882, w_000_883, w_000_884, w_000_885, w_000_886, w_000_887, w_000_888, w_000_889, w_000_890, w_000_891, w_000_892, w_000_893, w_000_894, w_000_895, w_000_896, w_000_897, w_000_898, w_000_899, w_000_900, w_000_901, w_000_902, w_000_903, w_000_904, w_000_905, w_000_906, w_000_907, w_000_908, w_000_909, w_000_910, w_000_911, w_000_912, w_000_913, w_000_914, w_000_915, w_000_916, w_000_917, w_000_918, w_000_919, w_000_920, w_000_921, w_000_922, w_000_923, w_000_924, w_000_925, w_000_926, w_000_927, w_000_928, w_000_929, w_000_930, w_000_931, w_000_932, w_000_933, w_000_935, w_000_936, w_000_937, w_000_938, w_000_939, w_000_940, w_000_941, w_000_942, w_000_943, w_000_944, w_000_945, w_000_946, w_000_947, w_000_948, w_000_949, w_000_950, w_000_951, w_000_952, w_000_953, w_000_954, w_000_955, w_000_956, w_000_957, w_000_958, w_000_959, w_000_960, w_000_961, w_000_962, w_000_963, w_000_964, w_000_965, w_000_966, w_000_967, w_000_968, w_000_969, w_000_970, w_000_971, w_000_972, w_000_973, w_000_974, w_000_975, w_000_976, w_000_977, w_000_978, w_000_979, w_000_980, w_000_981, w_000_982, w_000_983, w_000_984, w_000_985, w_000_986, w_000_987, w_000_988, w_000_989, w_000_990, w_000_991, w_000_992, w_000_993, w_000_994, w_000_995, w_000_996, w_000_997, w_000_998, w_000_999, w_000_1000, w_000_1001, w_000_1002, w_000_1003, w_000_1004, w_000_1005, w_000_1006, w_000_1007, w_000_1008, w_000_1009, w_000_1010, w_000_1011, w_000_1012, w_000_1013, w_000_1014, w_000_1015, w_000_1016, w_000_1017, w_000_1018, w_000_1019, w_000_1020, w_000_1021, w_000_1022, w_000_1023, w_000_1024, w_000_1025, w_000_1026, w_000_1027, w_000_1028, w_000_1029, w_000_1030, w_000_1031, w_000_1032, w_000_1033, w_000_1034, w_000_1035, w_000_1036, w_000_1037, w_000_1038, w_000_1039, w_000_1040, w_000_1041, w_000_1042, w_000_1043, w_000_1044, w_000_1045, w_000_1046, w_000_1047, w_000_1048, w_000_1049, w_000_1050, w_000_1051, w_000_1052, w_000_1053, w_000_1054, w_000_1055, w_000_1056, w_000_1057, w_000_1058, w_000_1060, w_000_1061, w_000_1062, w_000_1063, w_000_1064, w_000_1065, w_000_1066, w_000_1067, w_000_1068, w_000_1069, w_000_1070, w_000_1071, w_000_1072, w_000_1073, w_000_1074, w_000_1075, w_000_1076, w_000_1077, w_000_1078, w_000_1079, w_000_1080, w_000_1081, w_000_1082, w_000_1083, w_000_1084, w_000_1085, w_000_1086, w_000_1087, w_000_1088, w_000_1089, w_000_1090, w_000_1091, w_000_1093, w_000_1094, w_000_1095, w_000_1096, w_000_1097, w_000_1098, w_000_1099, w_000_1101, w_000_1102, w_000_1103, w_000_1104, w_000_1105, w_000_1106, w_000_1107, w_000_1108, w_000_1109, w_000_1110, w_000_1111, w_000_1112, w_000_1113, w_000_1114, w_000_1115, w_000_1116, w_000_1117, w_000_1118, w_000_1119, w_000_1120, w_000_1121, w_000_1122, w_000_1123, w_000_1124, w_000_1125, w_000_1126, w_000_1127, w_000_1128, w_000_1129, w_000_1130, w_000_1131, w_000_1132, w_000_1133, w_000_1134, w_000_1136, w_000_1137, w_000_1138, w_000_1139, w_000_1140, w_000_1141, w_000_1142, w_000_1143, w_000_1144, w_000_1145, w_000_1146, w_000_1147, w_000_1148, w_000_1149, w_000_1150, w_000_1151, w_000_1152, w_000_1153, w_000_1154, w_000_1155, w_000_1156, w_000_1157, w_000_1158, w_000_1159, w_000_1160, w_000_1161, w_000_1162, w_000_1163, w_000_1165, w_000_1166, w_000_1168, w_000_1169, w_000_1171, w_000_1172, w_000_1173, w_000_1174, w_000_1175, w_000_1176, w_000_1177, w_000_1178, w_000_1179, w_000_1180, w_000_1181, w_000_1182, w_000_1183, w_000_1184, w_000_1185, w_000_1186, w_000_1187, w_000_1188, w_000_1189, w_000_1190, w_000_1191, w_000_1192, w_000_1193, w_000_1194, w_000_1195, w_000_1196, w_000_1197, w_000_1198, w_000_1199, w_000_1200, w_000_1201, w_000_1202, w_000_1203, w_000_1204, w_000_1205, w_000_1206, w_000_1207, w_000_1208, w_000_1209, w_000_1210, w_000_1211, w_000_1212, w_000_1213, w_000_1214, w_000_1215, w_000_1216, w_000_1217, w_000_1218, w_000_1219, w_000_1220, w_000_1221, w_000_1222, w_000_1223, w_000_1224, w_000_1225, w_000_1226, w_000_1227, w_000_1228, w_000_1229, w_000_1230, w_000_1231, w_000_1232, w_000_1233, w_000_1234, w_000_1235, w_000_1236, w_000_1237, w_000_1238, w_000_1239, w_000_1240, w_000_1241, w_000_1242, w_000_1243, w_000_1244, w_000_1245, w_000_1246, w_000_1247, w_000_1248, w_000_1249, w_000_1250, w_000_1251, w_000_1252, w_000_1253, w_000_1254, w_000_1255, w_000_1256, w_000_1257, w_000_1258, w_000_1259, w_000_1260, w_000_1261, w_000_1262, w_000_1264, w_000_1265, w_000_1266, w_000_1267, w_000_1268, w_000_1270, w_000_1271, w_000_1272, w_000_1274, w_000_1275, w_000_1276, w_000_1277, w_000_1278, w_000_1279, w_000_1282, w_000_1283, w_000_1284, w_000_1285, w_000_1286, w_000_1287, w_000_1288, w_000_1289, w_000_1290, w_000_1291, w_000_1293, w_000_1294, w_000_1295, w_000_1296, w_000_1297, w_000_1298, w_000_1299, w_000_1300, w_000_1301, w_000_1302, w_000_1303, w_000_1304, w_000_1305, w_000_1306, w_000_1307, w_000_1308, w_000_1309, w_000_1310, w_000_1311, w_000_1312, w_000_1313, w_000_1314, w_000_1315, w_000_1316, w_000_1317, w_000_1318, w_000_1320, w_000_1321, w_000_1322, w_000_1323, w_000_1324, w_000_1325, w_000_1326, w_000_1327, w_000_1328, w_000_1329, w_000_1330, w_000_1331, w_000_1332, w_000_1333, w_000_1334, w_000_1335, w_000_1338, w_000_1339, w_000_1340, w_000_1341, w_000_1342, w_000_1343, w_000_1344, w_000_1345, w_000_1346, w_000_1347, w_000_1348, w_000_1349, w_000_1350, w_000_1351, w_000_1352, w_000_1353, w_000_1354, w_000_1355, w_000_1356, w_000_1357, w_000_1358, w_000_1359, w_000_1360, w_000_1361, w_000_1362, w_000_1363, w_000_1365, w_000_1366, w_000_1367, w_000_1368, w_000_1369, w_000_1370, w_000_1371, w_000_1372, w_000_1373, w_000_1374, w_000_1375, w_000_1376, w_000_1377, w_000_1378, w_000_1379, w_000_1380, w_000_1381, w_000_1382, w_000_1383, w_000_1385, w_000_1386, w_000_1387, w_000_1388, w_000_1389, w_000_1390, w_000_1391, w_000_1392, w_000_1393, w_000_1394, w_000_1395, w_000_1396, w_000_1397, w_000_1398, w_000_1399, w_000_1400, w_000_1401, w_000_1402, w_000_1403, w_000_1405, w_000_1406, w_000_1407, w_000_1408, w_000_1409, w_000_1410, w_000_1411, w_000_1412, w_000_1413, w_000_1414, w_000_1415, w_000_1417, w_000_1418, w_000_1419, w_000_1421, w_000_1422, w_000_1423, w_000_1424, w_000_1425, w_000_1426, w_000_1427, w_000_1428, w_000_1429, w_000_1430, w_000_1431, w_000_1432, w_000_1433, w_000_1434, w_000_1435, w_000_1436, w_000_1437, w_000_1438, w_000_1439, w_000_1440, w_000_1441, w_000_1442, w_000_1443, w_000_1444, w_000_1445, w_000_1447, w_000_1448, w_000_1449, w_000_1450, w_000_1451, w_000_1452, w_000_1453, w_000_1454, w_000_1455, w_000_1457, w_000_1458, w_000_1459, w_000_1460, w_000_1461, w_000_1462, w_000_1463, w_000_1464, w_000_1465, w_000_1466, w_000_1467, w_000_1469, w_000_1470, w_000_1471, w_000_1472, w_000_1473, w_000_1474, w_000_1475, w_000_1476, w_000_1477, w_000_1478, w_000_1480, w_000_1481, w_000_1482, w_000_1483, w_000_1484, w_000_1485, w_000_1486, w_000_1487, w_000_1488, w_000_1489, w_000_1490, w_000_1491, w_000_1492, w_000_1493, w_000_1494, w_000_1495, w_000_1496, w_000_1497, w_000_1498, w_000_1499, w_000_1500, w_000_1501, w_000_1502, w_000_1503, w_000_1504, w_000_1505, w_000_1506, w_000_1507, w_000_1508, w_000_1509, w_000_1510, w_000_1511, w_000_1512, w_000_1513, w_000_1514, w_000_1515, w_000_1516, w_000_1518, w_000_1519, w_000_1520, w_000_1521, w_000_1522, w_000_1523, w_000_1524, w_000_1525, w_000_1526, w_000_1527, w_000_1528, w_000_1529, w_000_1530, w_000_1531, w_000_1532, w_000_1533, w_000_1534, w_000_1535, w_000_1536, w_000_1537, w_000_1538, w_000_1539, w_000_1540, w_000_1541, w_000_1542, w_000_1543, w_000_1544, w_000_1545, w_000_1546, w_000_1547, w_000_1548, w_000_1549, w_000_1550, w_000_1551, w_000_1552, w_000_1553, w_000_1554, w_000_1555, w_000_1556, w_000_1557, w_000_1558, w_000_1559, w_000_1560, w_000_1561, w_000_1562, w_000_1563, w_000_1564, w_000_1565, w_000_1566, w_000_1567, w_000_1568, w_000_1569, w_000_1570, w_000_1571, w_000_1572, w_000_1573, w_000_1574, w_000_1575, w_000_1576, w_000_1577, w_000_1578, w_000_1579, w_000_1580, w_000_1581, w_000_1583, w_000_1584, w_000_1585, w_000_1586, w_000_1587, w_000_1588, w_000_1589, w_000_1590, w_000_1591, w_000_1592, w_000_1593, w_000_1594, w_000_1595, w_000_1596, w_000_1597, w_000_1598, w_000_1599, w_000_1600, w_000_1601, w_000_1602, w_000_1603, w_000_1604, w_000_1605, w_000_1606, w_000_1607, w_000_1608, w_000_1609, w_000_1610, w_000_1611, w_000_1612, w_000_1613, w_000_1614, w_000_1615, w_000_1616, w_000_1617, w_000_1618, w_000_1619, w_000_1620, w_000_1621, w_000_1622, w_000_1623, w_000_1624, w_000_1625, w_000_1626, w_000_1627, w_000_1628, w_000_1629, w_000_1630, w_000_1631, w_000_1632, w_000_1633, w_000_1634, w_000_1635, w_000_1636, w_000_1637, w_000_1638, w_000_1639, w_000_1640, w_000_1641, w_000_1642, w_000_1643, w_000_1644, w_000_1645, w_000_1646, w_000_1647, w_000_1648, w_000_1649, w_000_1650, w_000_1651, w_000_1652, w_000_1653, w_000_1654, w_000_1655, w_000_1656, w_000_1657, w_000_1658, w_000_1659, w_000_1660, w_000_1661, w_000_1662, w_000_1663, w_000_1664, w_000_1665, w_000_1666, w_000_1667, w_000_1669, w_000_1671, w_000_1672, w_000_1673, w_000_1674, w_000_1675, w_000_1676, w_000_1677, w_000_1678, w_000_1679, w_000_1680, w_000_1682, w_000_1683, w_000_1684, w_000_1685, w_000_1686, w_000_1687, w_000_1688, w_000_1690, w_000_1691, w_000_1692, w_000_1693, w_000_1694, w_000_1695, w_000_1696, w_000_1698, w_000_1699, w_000_1700, w_000_1701, w_000_1702, w_000_1703, w_000_1704, w_000_1705, w_000_1706, w_000_1707, w_000_1709, w_000_1710, w_000_1711, w_000_1712, w_000_1713, w_000_1716, w_000_1717, w_000_1719, w_000_1720, w_000_1722, w_000_1723, w_000_1725, w_000_1726, w_000_1727, w_000_1728, w_000_1729, w_000_1730, w_000_1732, w_000_1733, w_000_1734, w_000_1736, w_000_1737, w_000_1739, w_000_1740, w_000_1741, w_000_1742, w_000_1744, w_000_1745, w_000_1746, w_000_1747, w_000_1748, w_000_1749, w_000_1752, w_000_1753, w_000_1754, w_000_1755, w_000_1756, w_000_1757, w_000_1758, w_000_1759, w_000_1760, w_000_1761, w_000_1762, w_000_1763, w_000_1764, w_000_1765, w_000_1766, w_000_1768, w_000_1769, w_000_1770, w_000_1771, w_000_1772, w_000_1774, w_000_1775, w_000_1776, w_000_1778, w_000_1779, w_000_1780, w_000_1781, w_000_1782, w_000_1783, w_000_1784, w_000_1785, w_000_1787, w_000_1788, w_000_1789, w_000_1790, w_000_1791, w_000_1792, w_000_1794, w_000_1795, w_000_1796, w_000_1797, w_000_1800, w_000_1801, w_000_1802, w_000_1803, w_000_1804, w_000_1805, w_000_1806, w_000_1807, w_000_1808, w_000_1809, w_000_1810, w_000_1811, w_000_1812, w_000_1813, w_000_1814, w_000_1815, w_000_1816, w_000_1817, w_000_1818, w_000_1819, w_000_1820, w_000_1821, w_000_1822, w_000_1823, w_000_1824, w_000_1826, w_000_1827, w_000_1828, w_000_1829, w_000_1830, w_000_1831, w_000_1832, w_000_1833, w_000_1834, w_000_1835, w_000_1836, w_000_1837, w_000_1838, w_000_1839, w_000_1840, w_000_1841, w_000_1842, w_000_1843, w_000_1844, w_000_1845, w_000_1846, w_000_1847, w_000_1848, w_000_1849, w_000_1850, w_000_1851, w_000_1852, w_000_1857, w_000_1859, w_000_1861, w_000_1862, w_000_1863, w_000_1864, w_000_1865, w_000_1866, w_000_1868, w_000_1869, w_000_1870, w_000_1871, w_000_1873, w_000_1875, w_000_1876, w_000_1877, w_000_1878, w_000_1879, w_000_1880, w_000_1881, w_000_1882, w_000_1883, w_000_1885, w_000_1886, w_000_1887, w_000_1888, w_000_1889, w_000_1890, w_000_1893, w_000_1894, w_000_1895, w_000_1896, w_000_1899, w_000_1900, w_000_1902, w_000_1904, w_000_1905, w_000_1906, w_000_1907, w_000_1908, w_000_1909, w_000_1910, w_000_1912, w_000_1913, w_000_1914, w_000_1916, w_000_1917, w_000_1921, w_000_1922, w_000_1923, w_000_1924, w_000_1925, w_000_1926, w_000_1929, w_000_1931, w_000_1932, w_000_1935, w_000_1939, w_000_1942, w_000_1943, w_000_1946, w_000_1947, w_000_1949, w_000_1951, w_000_1962, w_000_1969, w_000_1971, w_000_1975, w_000_1977, w_2000_000, w_2000_001, w_2000_002, w_2000_003, w_2000_004, w_2000_005, w_2000_006, w_2000_007, w_2000_008, w_2000_009, w_2000_010, w_2000_011, w_2000_012, w_2000_013, w_2000_014, w_2000_015, w_2000_016, w_2000_017, w_2000_018, w_2000_019, w_2000_020, w_2000_021, w_2000_022, w_2000_023, w_2000_024, w_2000_025, w_2000_026, w_2000_027, w_2000_028, w_2000_029, w_2000_030, w_2000_031, w_2000_032, w_2000_033, w_2000_034, w_2000_035, w_2000_036, w_2000_037, w_2000_038, w_2000_039, w_2000_040, w_2000_041, w_2000_042, w_2000_043, w_2000_044, w_2000_045, w_2000_046, w_2000_047, w_2000_048, w_2000_049, w_2000_050, w_2000_051, w_2000_052, w_2000_053, w_2000_054, w_2000_055, w_2000_056, w_2000_057, w_2000_058, w_2000_059, w_2000_060, w_2000_061, w_2000_062, w_2000_063, w_2000_064, w_2000_065, w_2000_066, w_2000_067, w_2000_068, w_2000_069, w_2000_070, w_2000_071, w_2000_072, w_2000_073, w_2000_074, w_2000_075, w_2000_076, w_2000_077, w_2000_078, w_2000_079, w_2000_080, w_2000_081, w_2000_082, w_2000_083, w_2000_084, w_2000_085, w_2000_086, w_2000_087, w_2000_088, w_2000_089, w_2000_090, w_2000_091, w_2000_092, w_2000_093, w_2000_094, w_2000_095, w_2000_096, w_2000_097, w_2000_098, w_2000_099, w_2000_100, w_2000_101, w_2000_102, w_2000_103, w_2000_104, w_2000_105, w_2000_106, w_2000_107, w_2000_108, w_2000_109, w_2000_110 );
  inout w_000_000, w_000_001, w_000_002, w_000_003, w_000_004, w_000_005, w_000_006, w_000_007, w_000_008, w_000_009, w_000_010, w_000_011, w_000_012, w_000_013, w_000_014, w_000_015, w_000_016, w_000_017, w_000_018, w_000_019, w_000_020, w_000_021, w_000_022, w_000_023, w_000_024, w_000_025, w_000_026, w_000_027, w_000_028, w_000_029, w_000_030, w_000_031, w_000_032, w_000_033, w_000_034, w_000_035, w_000_036, w_000_037, w_000_038, w_000_039, w_000_040, w_000_041, w_000_042, w_000_043, w_000_044, w_000_045, w_000_046, w_000_047, w_000_048, w_000_049, w_000_050, w_000_051, w_000_052, w_000_053, w_000_054, w_000_055, w_000_056, w_000_057, w_000_058, w_000_059, w_000_060, w_000_061, w_000_062, w_000_063, w_000_065, w_000_066, w_000_067, w_000_068, w_000_069, w_000_070, w_000_071, w_000_072, w_000_073, w_000_074, w_000_075, w_000_076, w_000_077, w_000_078, w_000_079, w_000_080, w_000_081, w_000_082, w_000_083, w_000_084, w_000_085, w_000_086, w_000_087, w_000_088, w_000_089, w_000_090, w_000_091, w_000_092, w_000_093, w_000_094, w_000_095, w_000_096, w_000_097, w_000_098, w_000_099, w_000_100, w_000_101, w_000_102, w_000_103, w_000_104, w_000_105, w_000_106, w_000_107, w_000_108, w_000_109, w_000_110, w_000_111, w_000_112, w_000_113, w_000_114, w_000_115, w_000_116, w_000_117, w_000_118, w_000_119, w_000_120, w_000_121, w_000_122, w_000_123, w_000_124, w_000_125, w_000_126, w_000_127, w_000_128, w_000_129, w_000_130, w_000_131, w_000_132, w_000_133, w_000_134, w_000_135, w_000_136, w_000_137, w_000_138, w_000_139, w_000_140, w_000_141, w_000_142, w_000_143, w_000_144, w_000_145, w_000_146, w_000_147, w_000_148, w_000_149, w_000_150, w_000_151, w_000_152, w_000_153, w_000_154, w_000_155, w_000_156, w_000_157, w_000_158, w_000_159, w_000_160, w_000_161, w_000_162, w_000_163, w_000_164, w_000_165, w_000_166, w_000_167, w_000_168, w_000_169, w_000_170, w_000_171, w_000_172, w_000_173, w_000_174, w_000_175, w_000_176, w_000_177, w_000_178, w_000_179, w_000_180, w_000_181, w_000_182, w_000_183, w_000_184, w_000_185, w_000_186, w_000_187, w_000_188, w_000_189, w_000_190, w_000_191, w_000_192, w_000_193, w_000_194, w_000_195, w_000_196, w_000_197, w_000_198, w_000_199, w_000_200, w_000_201, w_000_202, w_000_203, w_000_204, w_000_205, w_000_206, w_000_207, w_000_208, w_000_209, w_000_210, w_000_211, w_000_212, w_000_213, w_000_214, w_000_215, w_000_216, w_000_217, w_000_218, w_000_219, w_000_220, w_000_221, w_000_222, w_000_223, w_000_224, w_000_225, w_000_226, w_000_227, w_000_228, w_000_229, w_000_230, w_000_231, w_000_232, w_000_233, w_000_234, w_000_235, w_000_236, w_000_237, w_000_238, w_000_239, w_000_240, w_000_241, w_000_242, w_000_243, w_000_244, w_000_245, w_000_246, w_000_247, w_000_248, w_000_249, w_000_250, w_000_251, w_000_252, w_000_253, w_000_254, w_000_255, w_000_256, w_000_257, w_000_258, w_000_259, w_000_260, w_000_261, w_000_262, w_000_263, w_000_264, w_000_265, w_000_266, w_000_267, w_000_268, w_000_269, w_000_270, w_000_271, w_000_272, w_000_273, w_000_274, w_000_275, w_000_276, w_000_277, w_000_278, w_000_279, w_000_280, w_000_281, w_000_282, w_000_283, w_000_284, w_000_285, w_000_286, w_000_287, w_000_289, w_000_290, w_000_291, w_000_292, w_000_293, w_000_294, w_000_295, w_000_296, w_000_297, w_000_298, w_000_299, w_000_300, w_000_301, w_000_302, w_000_303, w_000_304, w_000_305, w_000_306, w_000_307, w_000_308, w_000_309, w_000_310, w_000_311, w_000_312, w_000_313, w_000_314, w_000_315, w_000_316, w_000_317, w_000_318, w_000_319, w_000_320, w_000_321, w_000_322, w_000_323, w_000_324, w_000_325, w_000_326, w_000_327, w_000_328, w_000_329, w_000_330, w_000_331, w_000_332, w_000_333, w_000_334, w_000_335, w_000_336, w_000_337, w_000_338, w_000_339, w_000_340, w_000_341, w_000_342, w_000_343, w_000_344, w_000_345, w_000_346, w_000_347, w_000_348, w_000_349, w_000_350, w_000_351, w_000_352, w_000_353, w_000_354, w_000_355, w_000_356, w_000_357, w_000_358, w_000_359, w_000_360, w_000_361, w_000_362, w_000_363, w_000_364, w_000_365, w_000_366, w_000_367, w_000_368, w_000_369, w_000_370, w_000_371, w_000_372, w_000_373, w_000_374, w_000_375, w_000_376, w_000_377, w_000_378, w_000_379, w_000_380, w_000_381, w_000_382, w_000_383, w_000_384, w_000_385, w_000_386, w_000_387, w_000_388, w_000_389, w_000_390, w_000_391, w_000_392, w_000_393, w_000_394, w_000_395, w_000_396, w_000_397, w_000_398, w_000_399, w_000_400, w_000_401, w_000_402, w_000_403, w_000_404, w_000_405, w_000_406, w_000_407, w_000_408, w_000_409, w_000_410, w_000_411, w_000_412, w_000_413, w_000_414, w_000_415, w_000_416, w_000_417, w_000_418, w_000_419, w_000_420, w_000_421, w_000_422, w_000_423, w_000_424, w_000_425, w_000_426, w_000_427, w_000_428, w_000_429, w_000_430, w_000_431, w_000_432, w_000_433, w_000_434, w_000_435, w_000_436, w_000_437, w_000_438, w_000_439, w_000_440, w_000_441, w_000_442, w_000_443, w_000_444, w_000_445, w_000_446, w_000_447, w_000_448, w_000_449, w_000_450, w_000_451, w_000_452, w_000_453, w_000_454, w_000_455, w_000_456, w_000_457, w_000_458, w_000_459, w_000_460, w_000_461, w_000_462, w_000_463, w_000_464, w_000_465, w_000_466, w_000_467, w_000_468, w_000_469, w_000_470, w_000_471, w_000_472, w_000_473, w_000_474, w_000_475, w_000_476, w_000_477, w_000_478, w_000_479, w_000_480, w_000_481, w_000_482, w_000_483, w_000_484, w_000_485, w_000_486, w_000_487, w_000_488, w_000_489, w_000_490, w_000_491, w_000_492, w_000_493, w_000_494, w_000_495, w_000_496, w_000_498, w_000_499, w_000_500, w_000_501, w_000_502, w_000_503, w_000_504, w_000_505, w_000_506, w_000_507, w_000_508, w_000_509, w_000_510, w_000_511, w_000_512, w_000_513, w_000_514, w_000_515, w_000_516, w_000_517, w_000_518, w_000_519, w_000_520, w_000_521, w_000_522, w_000_523, w_000_524, w_000_525, w_000_526, w_000_527, w_000_528, w_000_529, w_000_530, w_000_531, w_000_532, w_000_533, w_000_534, w_000_535, w_000_536, w_000_537, w_000_538, w_000_539, w_000_540, w_000_541, w_000_542, w_000_543, w_000_544, w_000_545, w_000_546, w_000_547, w_000_548, w_000_549, w_000_550, w_000_551, w_000_552, w_000_553, w_000_554, w_000_555, w_000_556, w_000_557, w_000_558, w_000_559, w_000_560, w_000_561, w_000_562, w_000_563, w_000_564, w_000_565, w_000_566, w_000_567, w_000_568, w_000_569, w_000_570, w_000_571, w_000_572, w_000_573, w_000_575, w_000_576, w_000_577, w_000_578, w_000_579, w_000_580, w_000_581, w_000_582, w_000_583, w_000_584, w_000_585, w_000_586, w_000_587, w_000_588, w_000_589, w_000_590, w_000_591, w_000_592, w_000_593, w_000_594, w_000_595, w_000_596, w_000_597, w_000_598, w_000_599, w_000_600, w_000_601, w_000_602, w_000_603, w_000_604, w_000_605, w_000_606, w_000_607, w_000_608, w_000_609, w_000_610, w_000_611, w_000_612, w_000_613, w_000_614, w_000_615, w_000_616, w_000_617, w_000_618, w_000_619, w_000_620, w_000_621, w_000_622, w_000_623, w_000_624, w_000_625, w_000_626, w_000_627, w_000_628, w_000_629, w_000_630, w_000_631, w_000_632, w_000_633, w_000_634, w_000_635, w_000_636, w_000_638, w_000_639, w_000_640, w_000_641, w_000_643, w_000_644, w_000_645, w_000_646, w_000_647, w_000_648, w_000_649, w_000_650, w_000_651, w_000_652, w_000_653, w_000_654, w_000_655, w_000_656, w_000_657, w_000_658, w_000_659, w_000_660, w_000_661, w_000_662, w_000_663, w_000_664, w_000_665, w_000_667, w_000_668, w_000_669, w_000_670, w_000_671, w_000_672, w_000_673, w_000_674, w_000_675, w_000_676, w_000_677, w_000_678, w_000_679, w_000_680, w_000_681, w_000_682, w_000_683, w_000_684, w_000_685, w_000_686, w_000_687, w_000_688, w_000_689, w_000_690, w_000_691, w_000_692, w_000_693, w_000_694, w_000_695, w_000_696, w_000_697, w_000_698, w_000_699, w_000_700, w_000_701, w_000_702, w_000_703, w_000_704, w_000_705, w_000_706, w_000_707, w_000_708, w_000_709, w_000_710, w_000_711, w_000_712, w_000_713, w_000_714, w_000_715, w_000_716, w_000_717, w_000_718, w_000_719, w_000_720, w_000_721, w_000_722, w_000_723, w_000_724, w_000_725, w_000_726, w_000_727, w_000_728, w_000_729, w_000_730, w_000_731, w_000_732, w_000_733, w_000_734, w_000_735, w_000_736, w_000_737, w_000_738, w_000_739, w_000_740, w_000_741, w_000_742, w_000_743, w_000_744, w_000_745, w_000_746, w_000_747, w_000_748, w_000_749, w_000_750, w_000_751, w_000_752, w_000_753, w_000_754, w_000_755, w_000_756, w_000_757, w_000_758, w_000_759, w_000_760, w_000_761, w_000_762, w_000_763, w_000_764, w_000_765, w_000_766, w_000_767, w_000_768, w_000_769, w_000_770, w_000_771, w_000_772, w_000_773, w_000_774, w_000_775, w_000_776, w_000_777, w_000_778, w_000_779, w_000_780, w_000_781, w_000_782, w_000_783, w_000_784, w_000_785, w_000_786, w_000_787, w_000_788, w_000_789, w_000_790, w_000_791, w_000_792, w_000_793, w_000_794, w_000_795, w_000_796, w_000_797, w_000_798, w_000_799, w_000_800, w_000_801, w_000_802, w_000_803, w_000_804, w_000_805, w_000_806, w_000_807, w_000_808, w_000_809, w_000_810, w_000_811, w_000_812, w_000_813, w_000_814, w_000_815, w_000_816, w_000_817, w_000_818, w_000_819, w_000_820, w_000_821, w_000_822, w_000_823, w_000_824, w_000_825, w_000_826, w_000_827, w_000_828, w_000_829, w_000_830, w_000_831, w_000_832, w_000_833, w_000_835, w_000_836, w_000_837, w_000_838, w_000_839, w_000_840, w_000_841, w_000_842, w_000_843, w_000_844, w_000_845, w_000_846, w_000_847, w_000_848, w_000_849, w_000_850, w_000_851, w_000_852, w_000_853, w_000_854, w_000_855, w_000_856, w_000_857, w_000_858, w_000_859, w_000_860, w_000_861, w_000_862, w_000_863, w_000_864, w_000_865, w_000_866, w_000_867, w_000_868, w_000_869, w_000_870, w_000_871, w_000_872, w_000_873, w_000_874, w_000_875, w_000_876, w_000_877, w_000_878, w_000_879, w_000_880, w_000_881, w_000_882, w_000_883, w_000_884, w_000_885, w_000_886, w_000_887, w_000_888, w_000_889, w_000_890, w_000_891, w_000_892, w_000_893, w_000_894, w_000_895, w_000_896, w_000_897, w_000_898, w_000_899, w_000_900, w_000_901, w_000_902, w_000_903, w_000_904, w_000_905, w_000_906, w_000_907, w_000_908, w_000_909, w_000_910, w_000_911, w_000_912, w_000_913, w_000_914, w_000_915, w_000_916, w_000_917, w_000_918, w_000_919, w_000_920, w_000_921, w_000_922, w_000_923, w_000_924, w_000_925, w_000_926, w_000_927, w_000_928, w_000_929, w_000_930, w_000_931, w_000_932, w_000_933, w_000_935, w_000_936, w_000_937, w_000_938, w_000_939, w_000_940, w_000_941, w_000_942, w_000_943, w_000_944, w_000_945, w_000_946, w_000_947, w_000_948, w_000_949, w_000_950, w_000_951, w_000_952, w_000_953, w_000_954, w_000_955, w_000_956, w_000_957, w_000_958, w_000_959, w_000_960, w_000_961, w_000_962, w_000_963, w_000_964, w_000_965, w_000_966, w_000_967, w_000_968, w_000_969, w_000_970, w_000_971, w_000_972, w_000_973, w_000_974, w_000_975, w_000_976, w_000_977, w_000_978, w_000_979, w_000_980, w_000_981, w_000_982, w_000_983, w_000_984, w_000_985, w_000_986, w_000_987, w_000_988, w_000_989, w_000_990, w_000_991, w_000_992, w_000_993, w_000_994, w_000_995, w_000_996, w_000_997, w_000_998, w_000_999, w_000_1000, w_000_1001, w_000_1002, w_000_1003, w_000_1004, w_000_1005, w_000_1006, w_000_1007, w_000_1008, w_000_1009, w_000_1010, w_000_1011, w_000_1012, w_000_1013, w_000_1014, w_000_1015, w_000_1016, w_000_1017, w_000_1018, w_000_1019, w_000_1020, w_000_1021, w_000_1022, w_000_1023, w_000_1024, w_000_1025, w_000_1026, w_000_1027, w_000_1028, w_000_1029, w_000_1030, w_000_1031, w_000_1032, w_000_1033, w_000_1034, w_000_1035, w_000_1036, w_000_1037, w_000_1038, w_000_1039, w_000_1040, w_000_1041, w_000_1042, w_000_1043, w_000_1044, w_000_1045, w_000_1046, w_000_1047, w_000_1048, w_000_1049, w_000_1050, w_000_1051, w_000_1052, w_000_1053, w_000_1054, w_000_1055, w_000_1056, w_000_1057, w_000_1058, w_000_1060, w_000_1061, w_000_1062, w_000_1063, w_000_1064, w_000_1065, w_000_1066, w_000_1067, w_000_1068, w_000_1069, w_000_1070, w_000_1071, w_000_1072, w_000_1073, w_000_1074, w_000_1075, w_000_1076, w_000_1077, w_000_1078, w_000_1079, w_000_1080, w_000_1081, w_000_1082, w_000_1083, w_000_1084, w_000_1085, w_000_1086, w_000_1087, w_000_1088, w_000_1089, w_000_1090, w_000_1091, w_000_1093, w_000_1094, w_000_1095, w_000_1096, w_000_1097, w_000_1098, w_000_1099, w_000_1101, w_000_1102, w_000_1103, w_000_1104, w_000_1105, w_000_1106, w_000_1107, w_000_1108, w_000_1109, w_000_1110, w_000_1111, w_000_1112, w_000_1113, w_000_1114, w_000_1115, w_000_1116, w_000_1117, w_000_1118, w_000_1119, w_000_1120, w_000_1121, w_000_1122, w_000_1123, w_000_1124, w_000_1125, w_000_1126, w_000_1127, w_000_1128, w_000_1129, w_000_1130, w_000_1131, w_000_1132, w_000_1133, w_000_1134, w_000_1136, w_000_1137, w_000_1138, w_000_1139, w_000_1140, w_000_1141, w_000_1142, w_000_1143, w_000_1144, w_000_1145, w_000_1146, w_000_1147, w_000_1148, w_000_1149, w_000_1150, w_000_1151, w_000_1152, w_000_1153, w_000_1154, w_000_1155, w_000_1156, w_000_1157, w_000_1158, w_000_1159, w_000_1160, w_000_1161, w_000_1162, w_000_1163, w_000_1165, w_000_1166, w_000_1168, w_000_1169, w_000_1171, w_000_1172, w_000_1173, w_000_1174, w_000_1175, w_000_1176, w_000_1177, w_000_1178, w_000_1179, w_000_1180, w_000_1181, w_000_1182, w_000_1183, w_000_1184, w_000_1185, w_000_1186, w_000_1187, w_000_1188, w_000_1189, w_000_1190, w_000_1191, w_000_1192, w_000_1193, w_000_1194, w_000_1195, w_000_1196, w_000_1197, w_000_1198, w_000_1199, w_000_1200, w_000_1201, w_000_1202, w_000_1203, w_000_1204, w_000_1205, w_000_1206, w_000_1207, w_000_1208, w_000_1209, w_000_1210, w_000_1211, w_000_1212, w_000_1213, w_000_1214, w_000_1215, w_000_1216, w_000_1217, w_000_1218, w_000_1219, w_000_1220, w_000_1221, w_000_1222, w_000_1223, w_000_1224, w_000_1225, w_000_1226, w_000_1227, w_000_1228, w_000_1229, w_000_1230, w_000_1231, w_000_1232, w_000_1233, w_000_1234, w_000_1235, w_000_1236, w_000_1237, w_000_1238, w_000_1239, w_000_1240, w_000_1241, w_000_1242, w_000_1243, w_000_1244, w_000_1245, w_000_1246, w_000_1247, w_000_1248, w_000_1249, w_000_1250, w_000_1251, w_000_1252, w_000_1253, w_000_1254, w_000_1255, w_000_1256, w_000_1257, w_000_1258, w_000_1259, w_000_1260, w_000_1261, w_000_1262, w_000_1264, w_000_1265, w_000_1266, w_000_1267, w_000_1268, w_000_1270, w_000_1271, w_000_1272, w_000_1274, w_000_1275, w_000_1276, w_000_1277, w_000_1278, w_000_1279, w_000_1282, w_000_1283, w_000_1284, w_000_1285, w_000_1286, w_000_1287, w_000_1288, w_000_1289, w_000_1290, w_000_1291, w_000_1293, w_000_1294, w_000_1295, w_000_1296, w_000_1297, w_000_1298, w_000_1299, w_000_1300, w_000_1301, w_000_1302, w_000_1303, w_000_1304, w_000_1305, w_000_1306, w_000_1307, w_000_1308, w_000_1309, w_000_1310, w_000_1311, w_000_1312, w_000_1313, w_000_1314, w_000_1315, w_000_1316, w_000_1317, w_000_1318, w_000_1320, w_000_1321, w_000_1322, w_000_1323, w_000_1324, w_000_1325, w_000_1326, w_000_1327, w_000_1328, w_000_1329, w_000_1330, w_000_1331, w_000_1332, w_000_1333, w_000_1334, w_000_1335, w_000_1338, w_000_1339, w_000_1340, w_000_1341, w_000_1342, w_000_1343, w_000_1344, w_000_1345, w_000_1346, w_000_1347, w_000_1348, w_000_1349, w_000_1350, w_000_1351, w_000_1352, w_000_1353, w_000_1354, w_000_1355, w_000_1356, w_000_1357, w_000_1358, w_000_1359, w_000_1360, w_000_1361, w_000_1362, w_000_1363, w_000_1365, w_000_1366, w_000_1367, w_000_1368, w_000_1369, w_000_1370, w_000_1371, w_000_1372, w_000_1373, w_000_1374, w_000_1375, w_000_1376, w_000_1377, w_000_1378, w_000_1379, w_000_1380, w_000_1381, w_000_1382, w_000_1383, w_000_1385, w_000_1386, w_000_1387, w_000_1388, w_000_1389, w_000_1390, w_000_1391, w_000_1392, w_000_1393, w_000_1394, w_000_1395, w_000_1396, w_000_1397, w_000_1398, w_000_1399, w_000_1400, w_000_1401, w_000_1402, w_000_1403, w_000_1405, w_000_1406, w_000_1407, w_000_1408, w_000_1409, w_000_1410, w_000_1411, w_000_1412, w_000_1413, w_000_1414, w_000_1415, w_000_1417, w_000_1418, w_000_1419, w_000_1421, w_000_1422, w_000_1423, w_000_1424, w_000_1425, w_000_1426, w_000_1427, w_000_1428, w_000_1429, w_000_1430, w_000_1431, w_000_1432, w_000_1433, w_000_1434, w_000_1435, w_000_1436, w_000_1437, w_000_1438, w_000_1439, w_000_1440, w_000_1441, w_000_1442, w_000_1443, w_000_1444, w_000_1445, w_000_1447, w_000_1448, w_000_1449, w_000_1450, w_000_1451, w_000_1452, w_000_1453, w_000_1454, w_000_1455, w_000_1457, w_000_1458, w_000_1459, w_000_1460, w_000_1461, w_000_1462, w_000_1463, w_000_1464, w_000_1465, w_000_1466, w_000_1467, w_000_1469, w_000_1470, w_000_1471, w_000_1472, w_000_1473, w_000_1474, w_000_1475, w_000_1476, w_000_1477, w_000_1478, w_000_1480, w_000_1481, w_000_1482, w_000_1483, w_000_1484, w_000_1485, w_000_1486, w_000_1487, w_000_1488, w_000_1489, w_000_1490, w_000_1491, w_000_1492, w_000_1493, w_000_1494, w_000_1495, w_000_1496, w_000_1497, w_000_1498, w_000_1499, w_000_1500, w_000_1501, w_000_1502, w_000_1503, w_000_1504, w_000_1505, w_000_1506, w_000_1507, w_000_1508, w_000_1509, w_000_1510, w_000_1511, w_000_1512, w_000_1513, w_000_1514, w_000_1515, w_000_1516, w_000_1518, w_000_1519, w_000_1520, w_000_1521, w_000_1522, w_000_1523, w_000_1524, w_000_1525, w_000_1526, w_000_1527, w_000_1528, w_000_1529, w_000_1530, w_000_1531, w_000_1532, w_000_1533, w_000_1534, w_000_1535, w_000_1536, w_000_1537, w_000_1538, w_000_1539, w_000_1540, w_000_1541, w_000_1542, w_000_1543, w_000_1544, w_000_1545, w_000_1546, w_000_1547, w_000_1548, w_000_1549, w_000_1550, w_000_1551, w_000_1552, w_000_1553, w_000_1554, w_000_1555, w_000_1556, w_000_1557, w_000_1558, w_000_1559, w_000_1560, w_000_1561, w_000_1562, w_000_1563, w_000_1564, w_000_1565, w_000_1566, w_000_1567, w_000_1568, w_000_1569, w_000_1570, w_000_1571, w_000_1572, w_000_1573, w_000_1574, w_000_1575, w_000_1576, w_000_1577, w_000_1578, w_000_1579, w_000_1580, w_000_1581, w_000_1583, w_000_1584, w_000_1585, w_000_1586, w_000_1587, w_000_1588, w_000_1589, w_000_1590, w_000_1591, w_000_1592, w_000_1593, w_000_1594, w_000_1595, w_000_1596, w_000_1597, w_000_1598, w_000_1599, w_000_1600, w_000_1601, w_000_1602, w_000_1603, w_000_1604, w_000_1605, w_000_1606, w_000_1607, w_000_1608, w_000_1609, w_000_1610, w_000_1611, w_000_1612, w_000_1613, w_000_1614, w_000_1615, w_000_1616, w_000_1617, w_000_1618, w_000_1619, w_000_1620, w_000_1621, w_000_1622, w_000_1623, w_000_1624, w_000_1625, w_000_1626, w_000_1627, w_000_1628, w_000_1629, w_000_1630, w_000_1631, w_000_1632, w_000_1633, w_000_1634, w_000_1635, w_000_1636, w_000_1637, w_000_1638, w_000_1639, w_000_1640, w_000_1641, w_000_1642, w_000_1643, w_000_1644, w_000_1645, w_000_1646, w_000_1647, w_000_1648, w_000_1649, w_000_1650, w_000_1651, w_000_1652, w_000_1653, w_000_1654, w_000_1655, w_000_1656, w_000_1657, w_000_1658, w_000_1659, w_000_1660, w_000_1661, w_000_1662, w_000_1663, w_000_1664, w_000_1665, w_000_1666, w_000_1667, w_000_1669, w_000_1671, w_000_1672, w_000_1673, w_000_1674, w_000_1675, w_000_1676, w_000_1677, w_000_1678, w_000_1679, w_000_1680, w_000_1682, w_000_1683, w_000_1684, w_000_1685, w_000_1686, w_000_1687, w_000_1688, w_000_1690, w_000_1691, w_000_1692, w_000_1693, w_000_1694, w_000_1695, w_000_1696, w_000_1698, w_000_1699, w_000_1700, w_000_1701, w_000_1702, w_000_1703, w_000_1704, w_000_1705, w_000_1706, w_000_1707, w_000_1709, w_000_1710, w_000_1711, w_000_1712, w_000_1713, w_000_1716, w_000_1717, w_000_1719, w_000_1720, w_000_1722, w_000_1723, w_000_1725, w_000_1726, w_000_1727, w_000_1728, w_000_1729, w_000_1730, w_000_1732, w_000_1733, w_000_1734, w_000_1736, w_000_1737, w_000_1739, w_000_1740, w_000_1741, w_000_1742, w_000_1744, w_000_1745, w_000_1746, w_000_1747, w_000_1748, w_000_1749, w_000_1752, w_000_1753, w_000_1754, w_000_1755, w_000_1756, w_000_1757, w_000_1758, w_000_1759, w_000_1760, w_000_1761, w_000_1762, w_000_1763, w_000_1764, w_000_1765, w_000_1766, w_000_1768, w_000_1769, w_000_1770, w_000_1771, w_000_1772, w_000_1774, w_000_1775, w_000_1776, w_000_1778, w_000_1779, w_000_1780, w_000_1781, w_000_1782, w_000_1783, w_000_1784, w_000_1785, w_000_1787, w_000_1788, w_000_1789, w_000_1790, w_000_1791, w_000_1792, w_000_1794, w_000_1795, w_000_1796, w_000_1797, w_000_1800, w_000_1801, w_000_1802, w_000_1803, w_000_1804, w_000_1805, w_000_1806, w_000_1807, w_000_1808, w_000_1809, w_000_1810, w_000_1811, w_000_1812, w_000_1813, w_000_1814, w_000_1815, w_000_1816, w_000_1817, w_000_1818, w_000_1819, w_000_1820, w_000_1821, w_000_1822, w_000_1823, w_000_1824, w_000_1826, w_000_1827, w_000_1828, w_000_1829, w_000_1830, w_000_1831, w_000_1832, w_000_1833, w_000_1834, w_000_1835, w_000_1836, w_000_1837, w_000_1838, w_000_1839, w_000_1840, w_000_1841, w_000_1842, w_000_1843, w_000_1844, w_000_1845, w_000_1846, w_000_1847, w_000_1848, w_000_1849, w_000_1850, w_000_1851, w_000_1852, w_000_1857, w_000_1859, w_000_1861, w_000_1862, w_000_1863, w_000_1864, w_000_1865, w_000_1866, w_000_1868, w_000_1869, w_000_1870, w_000_1871, w_000_1873, w_000_1875, w_000_1876, w_000_1877, w_000_1878, w_000_1879, w_000_1880, w_000_1881, w_000_1882, w_000_1883, w_000_1885, w_000_1886, w_000_1887, w_000_1888, w_000_1889, w_000_1890, w_000_1893, w_000_1894, w_000_1895, w_000_1896, w_000_1899, w_000_1900, w_000_1902, w_000_1904, w_000_1905, w_000_1906, w_000_1907, w_000_1908, w_000_1909, w_000_1910, w_000_1912, w_000_1913, w_000_1914, w_000_1916, w_000_1917, w_000_1921, w_000_1922, w_000_1923, w_000_1924, w_000_1925, w_000_1926, w_000_1929, w_000_1931, w_000_1932, w_000_1935, w_000_1939, w_000_1942, w_000_1943, w_000_1946, w_000_1947, w_000_1949, w_000_1951, w_000_1962, w_000_1969, w_000_1971, w_000_1975, w_000_1977;
  output w_2000_000, w_2000_001, w_2000_002, w_2000_003, w_2000_004, w_2000_005, w_2000_006, w_2000_007, w_2000_008, w_2000_009, w_2000_010, w_2000_011, w_2000_012, w_2000_013, w_2000_014, w_2000_015, w_2000_016, w_2000_017, w_2000_018, w_2000_019, w_2000_020, w_2000_021, w_2000_022, w_2000_023, w_2000_024, w_2000_025, w_2000_026, w_2000_027, w_2000_028, w_2000_029, w_2000_030, w_2000_031, w_2000_032, w_2000_033, w_2000_034, w_2000_035, w_2000_036, w_2000_037, w_2000_038, w_2000_039, w_2000_040, w_2000_041, w_2000_042, w_2000_043, w_2000_044, w_2000_045, w_2000_046, w_2000_047, w_2000_048, w_2000_049, w_2000_050, w_2000_051, w_2000_052, w_2000_053, w_2000_054, w_2000_055, w_2000_056, w_2000_057, w_2000_058, w_2000_059, w_2000_060, w_2000_061, w_2000_062, w_2000_063, w_2000_064, w_2000_065, w_2000_066, w_2000_067, w_2000_068, w_2000_069, w_2000_070, w_2000_071, w_2000_072, w_2000_073, w_2000_074, w_2000_075, w_2000_076, w_2000_077, w_2000_078, w_2000_079, w_2000_080, w_2000_081, w_2000_082, w_2000_083, w_2000_084, w_2000_085, w_2000_086, w_2000_087, w_2000_088, w_2000_089, w_2000_090, w_2000_091, w_2000_092, w_2000_093, w_2000_094, w_2000_095, w_2000_096, w_2000_097, w_2000_098, w_2000_099, w_2000_100, w_2000_101, w_2000_102, w_2000_103, w_2000_104, w_2000_105, w_2000_106, w_2000_107, w_2000_108, w_2000_109, w_2000_110;
  wire w_000_000, w_000_001, w_000_002, w_000_003, w_000_004, w_000_005, w_000_006, w_000_007, w_000_008, w_000_009, w_000_010, w_000_011, w_000_012, w_000_013, w_000_014, w_000_015, w_000_016, w_000_017, w_000_018, w_000_019, w_000_020, w_000_021, w_000_022, w_000_023, w_000_024, w_000_025, w_000_026, w_000_027, w_000_028, w_000_029, w_000_030, w_000_031, w_000_032, w_000_033, w_000_034, w_000_035, w_000_036, w_000_037, w_000_038, w_000_039, w_000_040, w_000_041, w_000_042, w_000_043, w_000_044, w_000_045, w_000_046, w_000_047, w_000_048, w_000_049, w_000_050, w_000_051, w_000_052, w_000_053, w_000_054, w_000_055, w_000_056, w_000_057, w_000_058, w_000_059, w_000_060, w_000_061, w_000_062, w_000_063, w_000_065, w_000_066, w_000_067, w_000_068, w_000_069, w_000_070, w_000_071, w_000_072, w_000_073, w_000_074, w_000_075, w_000_076, w_000_077, w_000_078, w_000_079, w_000_080, w_000_081, w_000_082, w_000_083, w_000_084, w_000_085, w_000_086, w_000_087, w_000_088, w_000_089, w_000_090, w_000_091, w_000_092, w_000_093, w_000_094, w_000_095, w_000_096, w_000_097, w_000_098, w_000_099, w_000_100, w_000_101, w_000_102, w_000_103, w_000_104, w_000_105, w_000_106, w_000_107, w_000_108, w_000_109, w_000_110, w_000_111, w_000_112, w_000_113, w_000_114, w_000_115, w_000_116, w_000_117, w_000_118, w_000_119, w_000_120, w_000_121, w_000_122, w_000_123, w_000_124, w_000_125, w_000_126, w_000_127, w_000_128, w_000_129, w_000_130, w_000_131, w_000_132, w_000_133, w_000_134, w_000_135, w_000_136, w_000_137, w_000_138, w_000_139, w_000_140, w_000_141, w_000_142, w_000_143, w_000_144, w_000_145, w_000_146, w_000_147, w_000_148, w_000_149, w_000_150, w_000_151, w_000_152, w_000_153, w_000_154, w_000_155, w_000_156, w_000_157, w_000_158, w_000_159, w_000_160, w_000_161, w_000_162, w_000_163, w_000_164, w_000_165, w_000_166, w_000_167, w_000_168, w_000_169, w_000_170, w_000_171, w_000_172, w_000_173, w_000_174, w_000_175, w_000_176, w_000_177, w_000_178, w_000_179, w_000_180, w_000_181, w_000_182, w_000_183, w_000_184, w_000_185, w_000_186, w_000_187, w_000_188, w_000_189, w_000_190, w_000_191, w_000_192, w_000_193, w_000_194, w_000_195, w_000_196, w_000_197, w_000_198, w_000_199, w_000_200, w_000_201, w_000_202, w_000_203, w_000_204, w_000_205, w_000_206, w_000_207, w_000_208, w_000_209, w_000_210, w_000_211, w_000_212, w_000_213, w_000_214, w_000_215, w_000_216, w_000_217, w_000_218, w_000_219, w_000_220, w_000_221, w_000_222, w_000_223, w_000_224, w_000_225, w_000_226, w_000_227, w_000_228, w_000_229, w_000_230, w_000_231, w_000_232, w_000_233, w_000_234, w_000_235, w_000_236, w_000_237, w_000_238, w_000_239, w_000_240, w_000_241, w_000_242, w_000_243, w_000_244, w_000_245, w_000_246, w_000_247, w_000_248, w_000_249, w_000_250, w_000_251, w_000_252, w_000_253, w_000_254, w_000_255, w_000_256, w_000_257, w_000_258, w_000_259, w_000_260, w_000_261, w_000_262, w_000_263, w_000_264, w_000_265, w_000_266, w_000_267, w_000_268, w_000_269, w_000_270, w_000_271, w_000_272, w_000_273, w_000_274, w_000_275, w_000_276, w_000_277, w_000_278, w_000_279, w_000_280, w_000_281, w_000_282, w_000_283, w_000_284, w_000_285, w_000_286, w_000_287, w_000_289, w_000_290, w_000_291, w_000_292, w_000_293, w_000_294, w_000_295, w_000_296, w_000_297, w_000_298, w_000_299, w_000_300, w_000_301, w_000_302, w_000_303, w_000_304, w_000_305, w_000_306, w_000_307, w_000_308, w_000_309, w_000_310, w_000_311, w_000_312, w_000_313, w_000_314, w_000_315, w_000_316, w_000_317, w_000_318, w_000_319, w_000_320, w_000_321, w_000_322, w_000_323, w_000_324, w_000_325, w_000_326, w_000_327, w_000_328, w_000_329, w_000_330, w_000_331, w_000_332, w_000_333, w_000_334, w_000_335, w_000_336, w_000_337, w_000_338, w_000_339, w_000_340, w_000_341, w_000_342, w_000_343, w_000_344, w_000_345, w_000_346, w_000_347, w_000_348, w_000_349, w_000_350, w_000_351, w_000_352, w_000_353, w_000_354, w_000_355, w_000_356, w_000_357, w_000_358, w_000_359, w_000_360, w_000_361, w_000_362, w_000_363, w_000_364, w_000_365, w_000_366, w_000_367, w_000_368, w_000_369, w_000_370, w_000_371, w_000_372, w_000_373, w_000_374, w_000_375, w_000_376, w_000_377, w_000_378, w_000_379, w_000_380, w_000_381, w_000_382, w_000_383, w_000_384, w_000_385, w_000_386, w_000_387, w_000_388, w_000_389, w_000_390, w_000_391, w_000_392, w_000_393, w_000_394, w_000_395, w_000_396, w_000_397, w_000_398, w_000_399, w_000_400, w_000_401, w_000_402, w_000_403, w_000_404, w_000_405, w_000_406, w_000_407, w_000_408, w_000_409, w_000_410, w_000_411, w_000_412, w_000_413, w_000_414, w_000_415, w_000_416, w_000_417, w_000_418, w_000_419, w_000_420, w_000_421, w_000_422, w_000_423, w_000_424, w_000_425, w_000_426, w_000_427, w_000_428, w_000_429, w_000_430, w_000_431, w_000_432, w_000_433, w_000_434, w_000_435, w_000_436, w_000_437, w_000_438, w_000_439, w_000_440, w_000_441, w_000_442, w_000_443, w_000_444, w_000_445, w_000_446, w_000_447, w_000_448, w_000_449, w_000_450, w_000_451, w_000_452, w_000_453, w_000_454, w_000_455, w_000_456, w_000_457, w_000_458, w_000_459, w_000_460, w_000_461, w_000_462, w_000_463, w_000_464, w_000_465, w_000_466, w_000_467, w_000_468, w_000_469, w_000_470, w_000_471, w_000_472, w_000_473, w_000_474, w_000_475, w_000_476, w_000_477, w_000_478, w_000_479, w_000_480, w_000_481, w_000_482, w_000_483, w_000_484, w_000_485, w_000_486, w_000_487, w_000_488, w_000_489, w_000_490, w_000_491, w_000_492, w_000_493, w_000_494, w_000_495, w_000_496, w_000_498, w_000_499, w_000_500, w_000_501, w_000_502, w_000_503, w_000_504, w_000_505, w_000_506, w_000_507, w_000_508, w_000_509, w_000_510, w_000_511, w_000_512, w_000_513, w_000_514, w_000_515, w_000_516, w_000_517, w_000_518, w_000_519, w_000_520, w_000_521, w_000_522, w_000_523, w_000_524, w_000_525, w_000_526, w_000_527, w_000_528, w_000_529, w_000_530, w_000_531, w_000_532, w_000_533, w_000_534, w_000_535, w_000_536, w_000_537, w_000_538, w_000_539, w_000_540, w_000_541, w_000_542, w_000_543, w_000_544, w_000_545, w_000_546, w_000_547, w_000_548, w_000_549, w_000_550, w_000_551, w_000_552, w_000_553, w_000_554, w_000_555, w_000_556, w_000_557, w_000_558, w_000_559, w_000_560, w_000_561, w_000_562, w_000_563, w_000_564, w_000_565, w_000_566, w_000_567, w_000_568, w_000_569, w_000_570, w_000_571, w_000_572, w_000_573, w_000_575, w_000_576, w_000_577, w_000_578, w_000_579, w_000_580, w_000_581, w_000_582, w_000_583, w_000_584, w_000_585, w_000_586, w_000_587, w_000_588, w_000_589, w_000_590, w_000_591, w_000_592, w_000_593, w_000_594, w_000_595, w_000_596, w_000_597, w_000_598, w_000_599, w_000_600, w_000_601, w_000_602, w_000_603, w_000_604, w_000_605, w_000_606, w_000_607, w_000_608, w_000_609, w_000_610, w_000_611, w_000_612, w_000_613, w_000_614, w_000_615, w_000_616, w_000_617, w_000_618, w_000_619, w_000_620, w_000_621, w_000_622, w_000_623, w_000_624, w_000_625, w_000_626, w_000_627, w_000_628, w_000_629, w_000_630, w_000_631, w_000_632, w_000_633, w_000_634, w_000_635, w_000_636, w_000_638, w_000_639, w_000_640, w_000_641, w_000_643, w_000_644, w_000_645, w_000_646, w_000_647, w_000_648, w_000_649, w_000_650, w_000_651, w_000_652, w_000_653, w_000_654, w_000_655, w_000_656, w_000_657, w_000_658, w_000_659, w_000_660, w_000_661, w_000_662, w_000_663, w_000_664, w_000_665, w_000_667, w_000_668, w_000_669, w_000_670, w_000_671, w_000_672, w_000_673, w_000_674, w_000_675, w_000_676, w_000_677, w_000_678, w_000_679, w_000_680, w_000_681, w_000_682, w_000_683, w_000_684, w_000_685, w_000_686, w_000_687, w_000_688, w_000_689, w_000_690, w_000_691, w_000_692, w_000_693, w_000_694, w_000_695, w_000_696, w_000_697, w_000_698, w_000_699, w_000_700, w_000_701, w_000_702, w_000_703, w_000_704, w_000_705, w_000_706, w_000_707, w_000_708, w_000_709, w_000_710, w_000_711, w_000_712, w_000_713, w_000_714, w_000_715, w_000_716, w_000_717, w_000_718, w_000_719, w_000_720, w_000_721, w_000_722, w_000_723, w_000_724, w_000_725, w_000_726, w_000_727, w_000_728, w_000_729, w_000_730, w_000_731, w_000_732, w_000_733, w_000_734, w_000_735, w_000_736, w_000_737, w_000_738, w_000_739, w_000_740, w_000_741, w_000_742, w_000_743, w_000_744, w_000_745, w_000_746, w_000_747, w_000_748, w_000_749, w_000_750, w_000_751, w_000_752, w_000_753, w_000_754, w_000_755, w_000_756, w_000_757, w_000_758, w_000_759, w_000_760, w_000_761, w_000_762, w_000_763, w_000_764, w_000_765, w_000_766, w_000_767, w_000_768, w_000_769, w_000_770, w_000_771, w_000_772, w_000_773, w_000_774, w_000_775, w_000_776, w_000_777, w_000_778, w_000_779, w_000_780, w_000_781, w_000_782, w_000_783, w_000_784, w_000_785, w_000_786, w_000_787, w_000_788, w_000_789, w_000_790, w_000_791, w_000_792, w_000_793, w_000_794, w_000_795, w_000_796, w_000_797, w_000_798, w_000_799, w_000_800, w_000_801, w_000_802, w_000_803, w_000_804, w_000_805, w_000_806, w_000_807, w_000_808, w_000_809, w_000_810, w_000_811, w_000_812, w_000_813, w_000_814, w_000_815, w_000_816, w_000_817, w_000_818, w_000_819, w_000_820, w_000_821, w_000_822, w_000_823, w_000_824, w_000_825, w_000_826, w_000_827, w_000_828, w_000_829, w_000_830, w_000_831, w_000_832, w_000_833, w_000_835, w_000_836, w_000_837, w_000_838, w_000_839, w_000_840, w_000_841, w_000_842, w_000_843, w_000_844, w_000_845, w_000_846, w_000_847, w_000_848, w_000_849, w_000_850, w_000_851, w_000_852, w_000_853, w_000_854, w_000_855, w_000_856, w_000_857, w_000_858, w_000_859, w_000_860, w_000_861, w_000_862, w_000_863, w_000_864, w_000_865, w_000_866, w_000_867, w_000_868, w_000_869, w_000_870, w_000_871, w_000_872, w_000_873, w_000_874, w_000_875, w_000_876, w_000_877, w_000_878, w_000_879, w_000_880, w_000_881, w_000_882, w_000_883, w_000_884, w_000_885, w_000_886, w_000_887, w_000_888, w_000_889, w_000_890, w_000_891, w_000_892, w_000_893, w_000_894, w_000_895, w_000_896, w_000_897, w_000_898, w_000_899, w_000_900, w_000_901, w_000_902, w_000_903, w_000_904, w_000_905, w_000_906, w_000_907, w_000_908, w_000_909, w_000_910, w_000_911, w_000_912, w_000_913, w_000_914, w_000_915, w_000_916, w_000_917, w_000_918, w_000_919, w_000_920, w_000_921, w_000_922, w_000_923, w_000_924, w_000_925, w_000_926, w_000_927, w_000_928, w_000_929, w_000_930, w_000_931, w_000_932, w_000_933, w_000_935, w_000_936, w_000_937, w_000_938, w_000_939, w_000_940, w_000_941, w_000_942, w_000_943, w_000_944, w_000_945, w_000_946, w_000_947, w_000_948, w_000_949, w_000_950, w_000_951, w_000_952, w_000_953, w_000_954, w_000_955, w_000_956, w_000_957, w_000_958, w_000_959, w_000_960, w_000_961, w_000_962, w_000_963, w_000_964, w_000_965, w_000_966, w_000_967, w_000_968, w_000_969, w_000_970, w_000_971, w_000_972, w_000_973, w_000_974, w_000_975, w_000_976, w_000_977, w_000_978, w_000_979, w_000_980, w_000_981, w_000_982, w_000_983, w_000_984, w_000_985, w_000_986, w_000_987, w_000_988, w_000_989, w_000_990, w_000_991, w_000_992, w_000_993, w_000_994, w_000_995, w_000_996, w_000_997, w_000_998, w_000_999, w_000_1000, w_000_1001, w_000_1002, w_000_1003, w_000_1004, w_000_1005, w_000_1006, w_000_1007, w_000_1008, w_000_1009, w_000_1010, w_000_1011, w_000_1012, w_000_1013, w_000_1014, w_000_1015, w_000_1016, w_000_1017, w_000_1018, w_000_1019, w_000_1020, w_000_1021, w_000_1022, w_000_1023, w_000_1024, w_000_1025, w_000_1026, w_000_1027, w_000_1028, w_000_1029, w_000_1030, w_000_1031, w_000_1032, w_000_1033, w_000_1034, w_000_1035, w_000_1036, w_000_1037, w_000_1038, w_000_1039, w_000_1040, w_000_1041, w_000_1042, w_000_1043, w_000_1044, w_000_1045, w_000_1046, w_000_1047, w_000_1048, w_000_1049, w_000_1050, w_000_1051, w_000_1052, w_000_1053, w_000_1054, w_000_1055, w_000_1056, w_000_1057, w_000_1058, w_000_1060, w_000_1061, w_000_1062, w_000_1063, w_000_1064, w_000_1065, w_000_1066, w_000_1067, w_000_1068, w_000_1069, w_000_1070, w_000_1071, w_000_1072, w_000_1073, w_000_1074, w_000_1075, w_000_1076, w_000_1077, w_000_1078, w_000_1079, w_000_1080, w_000_1081, w_000_1082, w_000_1083, w_000_1084, w_000_1085, w_000_1086, w_000_1087, w_000_1088, w_000_1089, w_000_1090, w_000_1091, w_000_1093, w_000_1094, w_000_1095, w_000_1096, w_000_1097, w_000_1098, w_000_1099, w_000_1101, w_000_1102, w_000_1103, w_000_1104, w_000_1105, w_000_1106, w_000_1107, w_000_1108, w_000_1109, w_000_1110, w_000_1111, w_000_1112, w_000_1113, w_000_1114, w_000_1115, w_000_1116, w_000_1117, w_000_1118, w_000_1119, w_000_1120, w_000_1121, w_000_1122, w_000_1123, w_000_1124, w_000_1125, w_000_1126, w_000_1127, w_000_1128, w_000_1129, w_000_1130, w_000_1131, w_000_1132, w_000_1133, w_000_1134, w_000_1136, w_000_1137, w_000_1138, w_000_1139, w_000_1140, w_000_1141, w_000_1142, w_000_1143, w_000_1144, w_000_1145, w_000_1146, w_000_1147, w_000_1148, w_000_1149, w_000_1150, w_000_1151, w_000_1152, w_000_1153, w_000_1154, w_000_1155, w_000_1156, w_000_1157, w_000_1158, w_000_1159, w_000_1160, w_000_1161, w_000_1162, w_000_1163, w_000_1165, w_000_1166, w_000_1168, w_000_1169, w_000_1171, w_000_1172, w_000_1173, w_000_1174, w_000_1175, w_000_1176, w_000_1177, w_000_1178, w_000_1179, w_000_1180, w_000_1181, w_000_1182, w_000_1183, w_000_1184, w_000_1185, w_000_1186, w_000_1187, w_000_1188, w_000_1189, w_000_1190, w_000_1191, w_000_1192, w_000_1193, w_000_1194, w_000_1195, w_000_1196, w_000_1197, w_000_1198, w_000_1199, w_000_1200, w_000_1201, w_000_1202, w_000_1203, w_000_1204, w_000_1205, w_000_1206, w_000_1207, w_000_1208, w_000_1209, w_000_1210, w_000_1211, w_000_1212, w_000_1213, w_000_1214, w_000_1215, w_000_1216, w_000_1217, w_000_1218, w_000_1219, w_000_1220, w_000_1221, w_000_1222, w_000_1223, w_000_1224, w_000_1225, w_000_1226, w_000_1227, w_000_1228, w_000_1229, w_000_1230, w_000_1231, w_000_1232, w_000_1233, w_000_1234, w_000_1235, w_000_1236, w_000_1237, w_000_1238, w_000_1239, w_000_1240, w_000_1241, w_000_1242, w_000_1243, w_000_1244, w_000_1245, w_000_1246, w_000_1247, w_000_1248, w_000_1249, w_000_1250, w_000_1251, w_000_1252, w_000_1253, w_000_1254, w_000_1255, w_000_1256, w_000_1257, w_000_1258, w_000_1259, w_000_1260, w_000_1261, w_000_1262, w_000_1264, w_000_1265, w_000_1266, w_000_1267, w_000_1268, w_000_1270, w_000_1271, w_000_1272, w_000_1274, w_000_1275, w_000_1276, w_000_1277, w_000_1278, w_000_1279, w_000_1282, w_000_1283, w_000_1284, w_000_1285, w_000_1286, w_000_1287, w_000_1288, w_000_1289, w_000_1290, w_000_1291, w_000_1293, w_000_1294, w_000_1295, w_000_1296, w_000_1297, w_000_1298, w_000_1299, w_000_1300, w_000_1301, w_000_1302, w_000_1303, w_000_1304, w_000_1305, w_000_1306, w_000_1307, w_000_1308, w_000_1309, w_000_1310, w_000_1311, w_000_1312, w_000_1313, w_000_1314, w_000_1315, w_000_1316, w_000_1317, w_000_1318, w_000_1320, w_000_1321, w_000_1322, w_000_1323, w_000_1324, w_000_1325, w_000_1326, w_000_1327, w_000_1328, w_000_1329, w_000_1330, w_000_1331, w_000_1332, w_000_1333, w_000_1334, w_000_1335, w_000_1338, w_000_1339, w_000_1340, w_000_1341, w_000_1342, w_000_1343, w_000_1344, w_000_1345, w_000_1346, w_000_1347, w_000_1348, w_000_1349, w_000_1350, w_000_1351, w_000_1352, w_000_1353, w_000_1354, w_000_1355, w_000_1356, w_000_1357, w_000_1358, w_000_1359, w_000_1360, w_000_1361, w_000_1362, w_000_1363, w_000_1365, w_000_1366, w_000_1367, w_000_1368, w_000_1369, w_000_1370, w_000_1371, w_000_1372, w_000_1373, w_000_1374, w_000_1375, w_000_1376, w_000_1377, w_000_1378, w_000_1379, w_000_1380, w_000_1381, w_000_1382, w_000_1383, w_000_1385, w_000_1386, w_000_1387, w_000_1388, w_000_1389, w_000_1390, w_000_1391, w_000_1392, w_000_1393, w_000_1394, w_000_1395, w_000_1396, w_000_1397, w_000_1398, w_000_1399, w_000_1400, w_000_1401, w_000_1402, w_000_1403, w_000_1405, w_000_1406, w_000_1407, w_000_1408, w_000_1409, w_000_1410, w_000_1411, w_000_1412, w_000_1413, w_000_1414, w_000_1415, w_000_1417, w_000_1418, w_000_1419, w_000_1421, w_000_1422, w_000_1423, w_000_1424, w_000_1425, w_000_1426, w_000_1427, w_000_1428, w_000_1429, w_000_1430, w_000_1431, w_000_1432, w_000_1433, w_000_1434, w_000_1435, w_000_1436, w_000_1437, w_000_1438, w_000_1439, w_000_1440, w_000_1441, w_000_1442, w_000_1443, w_000_1444, w_000_1445, w_000_1447, w_000_1448, w_000_1449, w_000_1450, w_000_1451, w_000_1452, w_000_1453, w_000_1454, w_000_1455, w_000_1457, w_000_1458, w_000_1459, w_000_1460, w_000_1461, w_000_1462, w_000_1463, w_000_1464, w_000_1465, w_000_1466, w_000_1467, w_000_1469, w_000_1470, w_000_1471, w_000_1472, w_000_1473, w_000_1474, w_000_1475, w_000_1476, w_000_1477, w_000_1478, w_000_1480, w_000_1481, w_000_1482, w_000_1483, w_000_1484, w_000_1485, w_000_1486, w_000_1487, w_000_1488, w_000_1489, w_000_1490, w_000_1491, w_000_1492, w_000_1493, w_000_1494, w_000_1495, w_000_1496, w_000_1497, w_000_1498, w_000_1499, w_000_1500, w_000_1501, w_000_1502, w_000_1503, w_000_1504, w_000_1505, w_000_1506, w_000_1507, w_000_1508, w_000_1509, w_000_1510, w_000_1511, w_000_1512, w_000_1513, w_000_1514, w_000_1515, w_000_1516, w_000_1518, w_000_1519, w_000_1520, w_000_1521, w_000_1522, w_000_1523, w_000_1524, w_000_1525, w_000_1526, w_000_1527, w_000_1528, w_000_1529, w_000_1530, w_000_1531, w_000_1532, w_000_1533, w_000_1534, w_000_1535, w_000_1536, w_000_1537, w_000_1538, w_000_1539, w_000_1540, w_000_1541, w_000_1542, w_000_1543, w_000_1544, w_000_1545, w_000_1546, w_000_1547, w_000_1548, w_000_1549, w_000_1550, w_000_1551, w_000_1552, w_000_1553, w_000_1554, w_000_1555, w_000_1556, w_000_1557, w_000_1558, w_000_1559, w_000_1560, w_000_1561, w_000_1562, w_000_1563, w_000_1564, w_000_1565, w_000_1566, w_000_1567, w_000_1568, w_000_1569, w_000_1570, w_000_1571, w_000_1572, w_000_1573, w_000_1574, w_000_1575, w_000_1576, w_000_1577, w_000_1578, w_000_1579, w_000_1580, w_000_1581, w_000_1583, w_000_1584, w_000_1585, w_000_1586, w_000_1587, w_000_1588, w_000_1589, w_000_1590, w_000_1591, w_000_1592, w_000_1593, w_000_1594, w_000_1595, w_000_1596, w_000_1597, w_000_1598, w_000_1599, w_000_1600, w_000_1601, w_000_1602, w_000_1603, w_000_1604, w_000_1605, w_000_1606, w_000_1607, w_000_1608, w_000_1609, w_000_1610, w_000_1611, w_000_1612, w_000_1613, w_000_1614, w_000_1615, w_000_1616, w_000_1617, w_000_1618, w_000_1619, w_000_1620, w_000_1621, w_000_1622, w_000_1623, w_000_1624, w_000_1625, w_000_1626, w_000_1627, w_000_1628, w_000_1629, w_000_1630, w_000_1631, w_000_1632, w_000_1633, w_000_1634, w_000_1635, w_000_1636, w_000_1637, w_000_1638, w_000_1639, w_000_1640, w_000_1641, w_000_1642, w_000_1643, w_000_1644, w_000_1645, w_000_1646, w_000_1647, w_000_1648, w_000_1649, w_000_1650, w_000_1651, w_000_1652, w_000_1653, w_000_1654, w_000_1655, w_000_1656, w_000_1657, w_000_1658, w_000_1659, w_000_1660, w_000_1661, w_000_1662, w_000_1663, w_000_1664, w_000_1665, w_000_1666, w_000_1667, w_000_1669, w_000_1671, w_000_1672, w_000_1673, w_000_1674, w_000_1675, w_000_1676, w_000_1677, w_000_1678, w_000_1679, w_000_1680, w_000_1682, w_000_1683, w_000_1684, w_000_1685, w_000_1686, w_000_1687, w_000_1688, w_000_1690, w_000_1691, w_000_1692, w_000_1693, w_000_1694, w_000_1695, w_000_1696, w_000_1698, w_000_1699, w_000_1700, w_000_1701, w_000_1702, w_000_1703, w_000_1704, w_000_1705, w_000_1706, w_000_1707, w_000_1709, w_000_1710, w_000_1711, w_000_1712, w_000_1713, w_000_1716, w_000_1717, w_000_1719, w_000_1720, w_000_1722, w_000_1723, w_000_1725, w_000_1726, w_000_1727, w_000_1728, w_000_1729, w_000_1730, w_000_1732, w_000_1733, w_000_1734, w_000_1736, w_000_1737, w_000_1739, w_000_1740, w_000_1741, w_000_1742, w_000_1744, w_000_1745, w_000_1746, w_000_1747, w_000_1748, w_000_1749, w_000_1752, w_000_1753, w_000_1754, w_000_1755, w_000_1756, w_000_1757, w_000_1758, w_000_1759, w_000_1760, w_000_1761, w_000_1762, w_000_1763, w_000_1764, w_000_1765, w_000_1766, w_000_1768, w_000_1769, w_000_1770, w_000_1771, w_000_1772, w_000_1774, w_000_1775, w_000_1776, w_000_1778, w_000_1779, w_000_1780, w_000_1781, w_000_1782, w_000_1783, w_000_1784, w_000_1785, w_000_1787, w_000_1788, w_000_1789, w_000_1790, w_000_1791, w_000_1792, w_000_1794, w_000_1795, w_000_1796, w_000_1797, w_000_1800, w_000_1801, w_000_1802, w_000_1803, w_000_1804, w_000_1805, w_000_1806, w_000_1807, w_000_1808, w_000_1809, w_000_1810, w_000_1811, w_000_1812, w_000_1813, w_000_1814, w_000_1815, w_000_1816, w_000_1817, w_000_1818, w_000_1819, w_000_1820, w_000_1821, w_000_1822, w_000_1823, w_000_1824, w_000_1826, w_000_1827, w_000_1828, w_000_1829, w_000_1830, w_000_1831, w_000_1832, w_000_1833, w_000_1834, w_000_1835, w_000_1836, w_000_1837, w_000_1838, w_000_1839, w_000_1840, w_000_1841, w_000_1842, w_000_1843, w_000_1844, w_000_1845, w_000_1846, w_000_1847, w_000_1848, w_000_1849, w_000_1850, w_000_1851, w_000_1852, w_000_1857, w_000_1859, w_000_1861, w_000_1862, w_000_1863, w_000_1864, w_000_1865, w_000_1866, w_000_1868, w_000_1869, w_000_1870, w_000_1871, w_000_1873, w_000_1875, w_000_1876, w_000_1877, w_000_1878, w_000_1879, w_000_1880, w_000_1881, w_000_1882, w_000_1883, w_000_1885, w_000_1886, w_000_1887, w_000_1888, w_000_1889, w_000_1890, w_000_1893, w_000_1894, w_000_1895, w_000_1896, w_000_1899, w_000_1900, w_000_1902, w_000_1904, w_000_1905, w_000_1906, w_000_1907, w_000_1908, w_000_1909, w_000_1910, w_000_1912, w_000_1913, w_000_1914, w_000_1916, w_000_1917, w_000_1921, w_000_1922, w_000_1923, w_000_1924, w_000_1925, w_000_1926, w_000_1929, w_000_1931, w_000_1932, w_000_1935, w_000_1939, w_000_1942, w_000_1943, w_000_1946, w_000_1947, w_000_1949, w_000_1951, w_000_1962, w_000_1969, w_000_1971, w_000_1975, w_000_1977;
  wire w_001_000, w_001_001, w_001_002, w_001_003, w_001_004, w_001_005, w_001_006, w_001_007, w_001_008, w_001_009, w_001_010, w_001_011, w_001_012, w_001_013, w_001_014, w_001_015, w_001_016, w_001_017, w_001_018, w_001_019, w_001_020, w_001_021, w_001_022, w_001_023, w_001_024, w_001_025, w_001_026, w_001_027, w_001_028, w_001_029, w_001_030, w_001_031, w_001_032, w_001_033, w_001_034, w_001_035, w_001_036, w_001_038, w_001_039, w_001_040, w_001_041, w_001_042, w_001_043, w_001_044, w_001_045, w_001_046, w_001_047, w_001_048, w_001_049, w_001_050, w_001_051, w_001_052, w_001_053, w_001_054, w_001_055, w_001_056, w_001_057, w_001_059, w_001_060, w_001_061, w_001_062, w_001_063, w_001_064, w_001_065, w_001_066, w_001_067, w_001_068, w_001_069, w_001_070, w_001_071, w_001_072, w_001_073, w_001_074, w_001_075, w_001_076, w_001_077, w_001_078, w_001_079, w_001_080, w_001_081, w_001_082, w_001_083, w_001_084, w_001_086, w_001_087, w_001_088, w_001_090, w_001_091, w_001_092, w_001_093, w_001_094, w_001_095, w_001_096, w_001_097, w_001_098, w_001_099, w_001_100, w_001_101, w_001_102, w_001_103, w_001_104, w_001_106, w_001_107, w_001_108, w_001_109, w_001_110, w_001_111, w_001_112, w_001_113, w_001_114, w_001_115, w_001_116, w_001_117, w_001_119, w_001_120, w_001_121, w_001_122, w_001_123, w_001_124, w_001_125, w_001_126, w_001_127, w_001_128, w_001_129, w_001_130, w_001_131, w_001_132, w_001_133, w_001_134, w_001_135, w_001_137, w_001_138, w_001_139, w_001_140, w_001_141, w_001_142, w_001_143, w_001_145, w_001_147, w_001_148, w_001_149, w_001_150, w_001_151, w_001_152, w_001_153, w_001_154, w_001_155, w_001_156, w_001_157, w_001_159, w_001_160, w_001_161, w_001_162, w_001_163, w_001_164, w_001_165, w_001_166, w_001_168, w_001_169, w_001_170, w_001_172, w_001_173, w_001_174, w_001_175, w_001_176, w_001_177, w_001_178, w_001_179, w_001_180, w_001_181, w_001_182, w_001_183, w_001_184, w_001_185, w_001_186, w_001_187, w_001_188, w_001_189, w_001_190, w_001_191, w_001_192, w_001_193, w_001_194, w_001_195, w_001_196, w_001_197, w_001_198, w_001_199, w_001_200, w_001_201, w_001_202, w_001_203, w_001_204, w_001_205, w_001_206, w_001_207, w_001_208, w_001_209, w_001_210, w_001_212, w_001_213, w_001_214, w_001_216, w_001_217, w_001_218, w_001_219, w_001_221, w_001_223, w_001_224, w_001_225, w_001_226, w_001_227, w_001_228, w_001_229, w_001_230, w_001_231, w_001_232, w_001_233, w_001_234, w_001_235, w_001_236, w_001_237, w_001_238, w_001_239, w_001_240, w_001_241, w_001_242, w_001_243, w_001_244, w_001_245, w_001_246, w_001_247, w_001_248, w_001_249, w_001_250, w_001_251, w_001_252, w_001_253, w_001_254, w_001_255, w_001_256, w_001_257, w_001_258, w_001_259, w_001_260, w_001_261, w_001_262, w_001_263, w_001_264, w_001_265, w_001_266, w_001_267, w_001_268, w_001_269, w_001_270, w_001_271, w_001_272, w_001_273, w_001_274, w_001_275, w_001_276, w_001_278, w_001_279, w_001_280, w_001_281, w_001_282, w_001_283, w_001_284, w_001_285, w_001_286, w_001_287, w_001_288, w_001_289, w_001_290, w_001_291, w_001_292, w_001_293, w_001_294, w_001_295, w_001_296, w_001_297, w_001_298, w_001_299, w_001_300, w_001_302, w_001_303, w_001_305, w_001_306, w_001_307, w_001_308, w_001_309, w_001_310, w_001_311, w_001_312, w_001_313, w_001_316, w_001_317, w_001_319, w_001_321, w_001_322, w_001_323, w_001_325, w_001_326, w_001_329, w_001_330, w_001_331, w_001_335, w_001_336, w_001_337, w_001_338, w_001_340, w_001_341, w_001_342, w_001_343, w_001_344, w_001_345, w_001_346, w_001_348, w_001_349, w_001_350, w_001_352, w_001_354, w_001_357, w_001_358, w_001_359, w_001_362, w_001_363, w_001_364, w_001_365, w_001_366, w_001_367, w_001_370, w_001_371, w_001_372, w_001_373, w_001_374, w_001_377, w_001_378, w_001_379, w_001_384, w_001_386, w_001_387, w_001_388, w_001_389, w_001_390, w_001_391, w_001_392, w_001_393, w_001_394, w_001_395, w_001_397, w_001_398, w_001_399, w_001_400, w_001_401, w_001_404, w_001_405, w_001_406, w_001_407, w_001_408, w_001_409, w_001_411, w_001_412, w_001_413, w_001_414, w_001_416, w_001_417, w_001_418, w_001_419, w_001_420, w_001_421, w_001_422, w_001_423, w_001_424, w_001_425, w_001_426, w_001_427, w_001_428, w_001_429, w_001_430, w_001_431, w_001_432, w_001_435, w_001_436, w_001_438, w_001_440, w_001_442, w_001_443, w_001_444, w_001_445, w_001_446, w_001_447, w_001_448, w_001_449, w_001_451, w_001_452, w_001_453, w_001_454, w_001_455, w_001_457, w_001_458, w_001_459, w_001_460, w_001_461, w_001_466, w_001_467, w_001_470, w_001_471, w_001_472, w_001_473, w_001_474, w_001_475, w_001_476, w_001_478, w_001_479, w_001_480, w_001_481, w_001_482, w_001_484, w_001_485, w_001_486, w_001_487, w_001_488, w_001_489, w_001_491, w_001_492, w_001_493, w_001_494, w_001_495, w_001_496, w_001_498, w_001_499, w_001_501, w_001_502, w_001_503, w_001_504, w_001_505, w_001_506, w_001_507, w_001_509, w_001_510, w_001_511, w_001_512, w_001_513, w_001_514, w_001_517, w_001_518, w_001_519, w_001_520, w_001_521, w_001_522, w_001_524, w_001_525, w_001_526, w_001_527, w_001_528, w_001_529, w_001_530, w_001_531, w_001_532, w_001_533, w_001_535, w_001_537, w_001_538, w_001_539, w_001_542, w_001_543, w_001_544, w_001_545, w_001_546, w_001_548, w_001_549, w_001_550, w_001_553, w_001_554, w_001_555, w_001_556, w_001_558, w_001_559, w_001_560, w_001_561, w_001_562, w_001_564, w_001_565, w_001_566, w_001_567, w_001_568, w_001_569, w_001_570, w_001_571, w_001_572, w_001_573, w_001_574, w_001_575, w_001_576, w_001_577, w_001_580, w_001_583, w_001_584, w_001_585, w_001_586, w_001_587, w_001_589, w_001_590, w_001_592, w_001_593, w_001_594, w_001_595, w_001_596, w_001_597, w_001_601, w_001_602, w_001_603, w_001_604, w_001_605, w_001_606, w_001_609, w_001_610, w_001_612, w_001_613, w_001_614, w_001_615, w_001_617, w_001_618, w_001_619, w_001_620, w_001_621, w_001_622, w_001_623, w_001_624, w_001_625, w_001_626, w_001_627, w_001_628, w_001_629, w_001_630, w_001_631, w_001_632, w_001_635, w_001_636, w_001_637, w_001_638, w_001_639, w_001_640, w_001_641, w_001_643, w_001_644, w_001_646, w_001_649, w_001_650, w_001_651, w_001_652, w_001_653, w_001_655, w_001_656, w_001_657, w_001_658, w_001_659, w_001_660, w_001_661, w_001_662, w_001_663, w_001_665, w_001_666, w_001_667, w_001_668, w_001_669, w_001_671, w_001_672, w_001_673, w_001_674, w_001_677, w_001_678, w_001_681, w_001_683, w_001_685, w_001_686, w_001_687, w_001_688, w_001_689, w_001_691, w_001_692, w_001_696, w_001_697, w_001_698, w_001_699, w_001_700, w_001_701, w_001_702, w_001_704, w_001_707, w_001_708, w_001_709, w_001_710, w_001_711, w_001_712, w_001_714, w_001_715, w_001_716, w_001_717, w_001_718, w_001_720, w_001_721, w_001_722, w_001_723, w_001_725, w_001_726, w_001_728, w_001_729, w_001_731, w_001_732, w_001_733, w_001_734, w_001_735, w_001_736, w_001_737, w_001_738, w_001_741, w_001_742, w_001_744, w_001_745, w_001_746, w_001_747, w_001_750, w_001_751, w_001_752, w_001_754, w_001_755, w_001_756, w_001_757, w_001_758, w_001_759, w_001_761, w_001_762, w_001_763, w_001_764, w_001_765, w_001_767, w_001_768, w_001_769, w_001_770, w_001_771, w_001_772, w_001_776, w_001_778, w_001_779, w_001_780, w_001_781, w_001_783, w_001_784, w_001_785, w_001_786, w_001_787, w_001_790, w_001_791, w_001_792, w_001_793, w_001_794, w_001_796, w_001_797, w_001_798, w_001_799, w_001_800, w_001_801, w_001_804, w_001_805, w_001_806, w_001_807, w_001_808, w_001_809, w_001_810, w_001_811, w_001_812, w_001_813, w_001_814, w_001_815, w_001_816, w_001_817, w_001_818, w_001_820, w_001_821, w_001_822, w_001_824, w_001_825, w_001_827, w_001_828, w_001_829, w_001_831, w_001_832, w_001_833, w_001_835, w_001_836, w_001_837, w_001_840, w_001_842, w_001_843, w_001_844, w_001_845, w_001_847, w_001_848, w_001_849, w_001_850, w_001_851, w_001_852, w_001_853, w_001_854, w_001_855, w_001_856, w_001_857, w_001_859, w_001_860, w_001_861, w_001_862, w_001_864, w_001_865, w_001_866, w_001_867, w_001_868, w_001_869, w_001_870, w_001_872, w_001_873, w_001_875, w_001_876, w_001_877, w_001_878, w_001_879, w_001_880, w_001_881, w_001_882, w_001_883, w_001_884, w_001_885, w_001_887, w_001_888, w_001_889, w_001_890, w_001_892, w_001_893, w_001_894, w_001_895, w_001_897, w_001_898, w_001_899, w_001_900, w_001_901, w_001_902, w_001_903, w_001_904, w_001_905, w_001_906, w_001_907, w_001_908, w_001_909, w_001_910, w_001_911, w_001_914, w_001_915, w_001_916, w_001_919, w_001_921, w_001_922, w_001_926, w_001_929, w_001_931, w_001_932, w_001_936, w_001_937, w_001_939, w_001_940, w_001_941, w_001_943, w_001_944, w_001_946, w_001_947, w_001_948, w_001_949, w_001_950, w_001_951, w_001_953, w_001_954, w_001_955, w_001_956, w_001_958, w_001_960, w_001_961, w_001_963, w_001_964, w_001_965, w_001_966, w_001_967, w_001_969, w_001_970, w_001_973, w_001_974, w_001_976, w_001_977, w_001_978, w_001_980, w_001_981, w_001_982, w_001_983, w_001_984, w_001_985, w_001_986, w_001_987, w_001_988, w_001_989, w_001_990, w_001_991, w_001_993, w_001_994, w_001_997, w_001_998, w_001_999, w_001_1000, w_001_1001, w_001_1002, w_001_1003, w_001_1005, w_001_1007, w_001_1008, w_001_1011, w_001_1012, w_001_1013, w_001_1014, w_001_1015, w_001_1019, w_001_1020, w_001_1022, w_001_1023, w_001_1025, w_001_1026, w_001_1027, w_001_1028, w_001_1030, w_001_1031, w_001_1033, w_001_1034, w_001_1035, w_001_1036, w_001_1037, w_001_1039, w_001_1040, w_001_1042, w_001_1044, w_001_1045, w_001_1046, w_001_1047, w_001_1049, w_001_1050, w_001_1051, w_001_1053, w_001_1054, w_001_1056, w_001_1057, w_001_1058, w_001_1059, w_001_1060, w_001_1061, w_001_1062, w_001_1063, w_001_1064, w_001_1065, w_001_1066, w_001_1067, w_001_1068, w_001_1070, w_001_1071, w_001_1072, w_001_1074, w_001_1076, w_001_1077, w_001_1078, w_001_1079, w_001_1081, w_001_1082, w_001_1083, w_001_1084, w_001_1085, w_001_1088, w_001_1089, w_001_1090, w_001_1092, w_001_1093, w_001_1094, w_001_1096, w_001_1097, w_001_1098, w_001_1099, w_001_1100, w_001_1101, w_001_1102, w_001_1104, w_001_1105, w_001_1106, w_001_1107, w_001_1108, w_001_1109, w_001_1111, w_001_1112, w_001_1113, w_001_1115, w_001_1117, w_001_1118, w_001_1119, w_001_1120, w_001_1121, w_001_1122, w_001_1123, w_001_1124, w_001_1125, w_001_1126, w_001_1127, w_001_1128, w_001_1129, w_001_1130, w_001_1131, w_001_1132, w_001_1133, w_001_1134, w_001_1135, w_001_1138, w_001_1140, w_001_1141, w_001_1142, w_001_1143, w_001_1144, w_001_1145, w_001_1146, w_001_1147, w_001_1148, w_001_1149, w_001_1151, w_001_1152, w_001_1153, w_001_1155, w_001_1156, w_001_1158, w_001_1159, w_001_1160, w_001_1161, w_001_1163, w_001_1164, w_001_1167, w_001_1170, w_001_1171, w_001_1172, w_001_1176, w_001_1177, w_001_1179, w_001_1181, w_001_1183, w_001_1184, w_001_1185, w_001_1186, w_001_1187, w_001_1188, w_001_1189, w_001_1191, w_001_1192, w_001_1193, w_001_1195, w_001_1196, w_001_1197, w_001_1198, w_001_1199, w_001_1200, w_001_1201, w_001_1202, w_001_1203, w_001_1204, w_001_1205, w_001_1206, w_001_1207, w_001_1209, w_001_1211, w_001_1212, w_001_1213, w_001_1215, w_001_1216, w_001_1217, w_001_1220, w_001_1221, w_001_1222, w_001_1225, w_001_1226, w_001_1227, w_001_1228, w_001_1229, w_001_1230, w_001_1231, w_001_1232, w_001_1233, w_001_1235, w_001_1236, w_001_1237, w_001_1238, w_001_1239, w_001_1240, w_001_1241, w_001_1242, w_001_1243, w_001_1246, w_001_1247, w_001_1248, w_001_1249, w_001_1250, w_001_1251, w_001_1253, w_001_1255, w_001_1256, w_001_1259, w_001_1260, w_001_1261, w_001_1262, w_001_1263, w_001_1264, w_001_1265, w_001_1266, w_001_1267, w_001_1268, w_001_1269, w_001_1270, w_001_1271, w_001_1272, w_001_1273, w_001_1274, w_001_1275, w_001_1276, w_001_1278, w_001_1279, w_001_1280, w_001_1281, w_001_1282, w_001_1284, w_001_1288, w_001_1289, w_001_1290, w_001_1293, w_001_1296, w_001_1298, w_001_1299, w_001_1300, w_001_1301, w_001_1302, w_001_1303, w_001_1304, w_001_1305, w_001_1306, w_001_1307, w_001_1308, w_001_1309, w_001_1310, w_001_1312, w_001_1314, w_001_1316, w_001_1317, w_001_1319, w_001_1320, w_001_1321, w_001_1322, w_001_1323, w_001_1324, w_001_1325, w_001_1327, w_001_1331, w_001_1332, w_001_1333, w_001_1335, w_001_1337, w_001_1339, w_001_1341, w_001_1342, w_001_1343, w_001_1345, w_001_1346, w_001_1349, w_001_1350, w_001_1351, w_001_1353, w_001_1354, w_001_1355, w_001_1356, w_001_1358, w_001_1359, w_001_1361, w_001_1362, w_001_1365, w_001_1366, w_001_1367, w_001_1369, w_001_1371, w_001_1373, w_001_1374, w_001_1376, w_001_1379, w_001_1380, w_001_1381, w_001_1382, w_001_1383, w_001_1384, w_001_1386, w_001_1387, w_001_1388, w_001_1390, w_001_1392, w_001_1393, w_001_1394, w_001_1396, w_001_1397, w_001_1398, w_001_1399, w_001_1400, w_001_1402, w_001_1403, w_001_1405, w_001_1406, w_001_1408, w_001_1409, w_001_1412, w_001_1413, w_001_1416, w_001_1417, w_001_1418, w_001_1422, w_001_1423, w_001_1424, w_001_1425, w_001_1426, w_001_1427, w_001_1428, w_001_1429, w_001_1430, w_001_1431, w_001_1432, w_001_1435, w_001_1436, w_001_1437, w_001_1438, w_001_1439, w_001_1440, w_001_1441, w_001_1444, w_001_1446, w_001_1447, w_001_1449, w_001_1452, w_001_1453, w_001_1454, w_001_1456, w_001_1457, w_001_1458, w_001_1459, w_001_1460, w_001_1461, w_001_1462, w_001_1463, w_001_1464, w_001_1465, w_001_1467, w_001_1469, w_001_1470, w_001_1474, w_001_1475, w_001_1476, w_001_1477, w_001_1479, w_001_1480, w_001_1482, w_001_1483, w_001_1484, w_001_1485, w_001_1486, w_001_1487, w_001_1488, w_001_1489, w_001_1491, w_001_1495, w_001_1496, w_001_1497, w_001_1498, w_001_1499, w_001_1500, w_001_1502, w_001_1503, w_001_1505, w_001_1506, w_001_1507, w_001_1508, w_001_1509, w_001_1511, w_001_1513, w_001_1514, w_001_1515, w_001_1516, w_001_1517, w_001_1520, w_001_1521, w_001_1522, w_001_1523, w_001_1524, w_001_1526, w_001_1527, w_001_1529, w_001_1531, w_001_1532, w_001_1533, w_001_1534, w_001_1536, w_001_1538, w_001_1540, w_001_1541, w_001_1544, w_001_1547, w_001_1548, w_001_1550, w_001_1551, w_001_1555, w_001_1556, w_001_1557, w_001_1559, w_001_1560, w_001_1561, w_001_1563, w_001_1564, w_001_1565, w_001_1566, w_001_1567, w_001_1568, w_001_1570, w_001_1571, w_001_1573, w_001_1575, w_001_1576, w_001_1578, w_001_1579, w_001_1580, w_001_1581, w_001_1582, w_001_1583, w_001_1585, w_001_1586, w_001_1587, w_001_1588, w_001_1589, w_001_1592, w_001_1593, w_001_1595, w_001_1597, w_001_1599, w_001_1600, w_001_1602, w_001_1603, w_001_1604, w_001_1605, w_001_1606, w_001_1607, w_001_1608, w_001_1609, w_001_1612, w_001_1613, w_001_1616, w_001_1617, w_001_1622, w_001_1625, w_001_1627, w_001_1628, w_001_1629, w_001_1630, w_001_1631, w_001_1632, w_001_1633, w_001_1634, w_001_1636, w_001_1637, w_001_1638, w_001_1639, w_001_1640, w_001_1641, w_001_1642, w_001_1643, w_001_1644, w_001_1645, w_001_1646, w_001_1647, w_001_1649, w_001_1651, w_001_1653, w_001_1654, w_001_1655, w_001_1656, w_001_1657, w_001_1659, w_001_1660, w_001_1661, w_001_1662, w_001_1664, w_001_1665, w_001_1666, w_001_1667, w_001_1669, w_001_1670, w_001_1671, w_001_1672, w_001_1673, w_001_1674, w_001_1675, w_001_1676, w_001_1677, w_001_1680, w_001_1681, w_001_1682, w_001_1683, w_001_1684, w_001_1685, w_001_1687, w_001_1688, w_001_1689;
  wire w_002_000, w_002_001, w_002_002, w_002_003, w_002_004, w_002_005, w_002_006, w_002_007, w_002_008, w_002_009, w_002_010, w_002_011, w_002_012, w_002_013, w_002_014, w_002_015, w_002_016, w_002_017, w_002_018, w_002_019, w_002_020, w_002_021, w_002_022, w_002_023, w_002_025, w_002_026, w_002_027, w_002_028, w_002_029, w_002_030, w_002_031, w_002_032, w_002_033, w_002_034, w_002_035, w_002_036, w_002_037, w_002_038, w_002_039, w_002_040, w_002_041, w_002_042, w_002_043, w_002_044, w_002_045, w_002_046, w_002_047, w_002_048, w_002_049, w_002_050, w_002_051, w_002_052, w_002_053, w_002_054, w_002_055, w_002_056, w_002_057, w_002_058, w_002_059, w_002_060, w_002_061, w_002_062, w_002_063, w_002_064, w_002_065, w_002_066, w_002_067, w_002_068, w_002_069, w_002_070, w_002_071, w_002_072, w_002_073, w_002_074, w_002_075, w_002_076, w_002_077, w_002_078, w_002_079, w_002_080, w_002_081, w_002_082, w_002_083, w_002_084, w_002_085, w_002_086, w_002_087, w_002_088, w_002_089, w_002_090, w_002_091, w_002_092, w_002_093, w_002_094, w_002_095, w_002_096, w_002_097, w_002_098, w_002_099, w_002_100, w_002_101, w_002_102, w_002_103, w_002_104, w_002_105, w_002_106, w_002_107, w_002_108, w_002_109, w_002_110, w_002_111, w_002_112, w_002_113, w_002_114, w_002_115, w_002_116, w_002_117, w_002_118, w_002_119, w_002_120, w_002_121, w_002_122, w_002_123, w_002_124, w_002_125, w_002_126, w_002_127, w_002_128, w_002_129, w_002_130, w_002_131, w_002_132, w_002_133, w_002_134, w_002_135, w_002_136, w_002_137, w_002_138, w_002_139, w_002_140, w_002_141, w_002_142, w_002_143, w_002_144, w_002_145, w_002_146, w_002_147, w_002_148, w_002_149, w_002_150, w_002_151, w_002_152, w_002_153, w_002_154, w_002_155, w_002_156, w_002_157, w_002_158, w_002_159, w_002_160, w_002_161, w_002_162, w_002_163, w_002_164, w_002_165, w_002_166, w_002_167, w_002_168, w_002_169, w_002_170, w_002_171, w_002_172, w_002_173, w_002_174, w_002_175, w_002_176, w_002_177, w_002_178, w_002_179, w_002_180, w_002_181, w_002_182, w_002_183, w_002_184, w_002_185, w_002_186, w_002_187, w_002_188, w_002_189, w_002_190, w_002_191, w_002_192, w_002_193, w_002_194, w_002_195, w_002_196, w_002_197, w_002_198, w_002_199, w_002_200, w_002_201, w_002_202, w_002_203, w_002_204, w_002_205, w_002_206, w_002_207, w_002_208, w_002_209, w_002_210, w_002_211, w_002_212, w_002_213, w_002_214, w_002_215, w_002_216, w_002_217, w_002_218, w_002_219, w_002_220, w_002_221, w_002_222, w_002_223, w_002_224, w_002_225, w_002_226, w_002_227, w_002_228, w_002_229, w_002_230, w_002_231, w_002_232, w_002_233, w_002_234, w_002_235, w_002_236, w_002_237, w_002_238, w_002_239, w_002_240, w_002_241, w_002_242, w_002_243, w_002_244, w_002_245, w_002_246, w_002_247, w_002_248, w_002_249, w_002_250, w_002_251, w_002_252, w_002_253, w_002_255, w_002_256, w_002_257, w_002_258, w_002_259, w_002_260, w_002_261, w_002_262, w_002_263, w_002_264, w_002_265, w_002_266, w_002_267, w_002_268, w_002_269, w_002_270, w_002_271, w_002_272, w_002_273, w_002_274, w_002_275, w_002_276, w_002_277, w_002_278, w_002_280, w_002_281, w_002_282, w_002_283, w_002_284, w_002_285, w_002_286, w_002_287, w_002_288, w_002_289, w_002_290, w_002_291, w_002_292, w_002_293, w_002_294, w_002_295, w_002_297, w_002_298, w_002_299, w_002_300, w_002_301, w_002_302, w_002_303, w_002_304, w_002_305, w_002_306, w_002_307, w_002_308, w_002_309, w_002_310, w_002_311, w_002_312, w_002_313, w_002_314, w_002_315, w_002_316, w_002_317, w_002_318, w_002_319, w_002_320, w_002_321, w_002_322, w_002_323, w_002_324, w_002_325, w_002_326, w_002_327, w_002_328, w_002_329, w_002_330, w_002_331, w_002_332, w_002_333, w_002_334, w_002_335, w_002_336, w_002_338, w_002_339, w_002_340, w_002_341, w_002_342, w_002_343, w_002_344, w_002_345, w_002_346, w_002_347, w_002_348, w_002_349, w_002_350, w_002_351, w_002_352, w_002_353, w_002_354, w_002_355, w_002_356, w_002_357, w_002_358, w_002_359, w_002_360, w_002_361, w_002_363, w_002_365, w_002_366, w_002_367, w_002_368, w_002_369, w_002_370, w_002_371, w_002_372, w_002_373, w_002_374, w_002_375, w_002_376, w_002_377, w_002_378, w_002_379, w_002_380, w_002_381, w_002_382, w_002_383, w_002_384, w_002_385, w_002_386, w_002_387, w_002_388, w_002_389, w_002_390, w_002_391, w_002_392, w_002_393, w_002_394, w_002_395, w_002_396, w_002_397, w_002_398, w_002_399, w_002_400, w_002_401, w_002_402, w_002_403, w_002_404, w_002_405, w_002_406, w_002_407, w_002_408, w_002_409, w_002_410, w_002_411, w_002_412, w_002_413, w_002_414, w_002_416, w_002_417, w_002_418, w_002_419, w_002_420, w_002_421, w_002_422, w_002_423, w_002_424, w_002_425, w_002_426, w_002_427, w_002_428, w_002_429, w_002_430, w_002_431, w_002_432, w_002_433, w_002_434, w_002_435, w_002_436, w_002_437, w_002_438, w_002_439, w_002_440, w_002_441, w_002_442, w_002_443, w_002_444, w_002_445, w_002_446, w_002_447, w_002_448, w_002_449, w_002_450, w_002_451, w_002_452, w_002_453, w_002_454, w_002_456, w_002_457, w_002_458, w_002_459, w_002_460, w_002_461, w_002_462, w_002_463, w_002_464, w_002_465, w_002_466, w_002_467, w_002_468, w_002_469, w_002_470, w_002_471, w_002_472, w_002_473, w_002_474, w_002_475, w_002_476, w_002_477, w_002_478, w_002_479, w_002_480, w_002_481, w_002_482, w_002_483, w_002_484, w_002_485, w_002_486, w_002_487, w_002_488, w_002_489, w_002_490, w_002_491, w_002_492, w_002_493, w_002_494, w_002_495, w_002_496, w_002_497, w_002_498, w_002_499, w_002_500, w_002_501, w_002_502, w_002_503, w_002_504, w_002_505, w_002_506, w_002_507, w_002_508, w_002_509, w_002_510, w_002_511, w_002_512, w_002_513, w_002_514, w_002_515, w_002_516, w_002_517, w_002_519, w_002_521, w_002_522, w_002_523, w_002_524, w_002_525, w_002_526, w_002_527, w_002_528, w_002_529, w_002_530, w_002_531, w_002_532, w_002_533, w_002_534, w_002_535, w_002_536, w_002_537, w_002_538, w_002_539, w_002_540, w_002_541, w_002_542, w_002_543, w_002_544, w_002_545, w_002_546, w_002_547, w_002_548, w_002_549, w_002_550, w_002_551, w_002_552, w_002_553, w_002_554, w_002_555, w_002_556, w_002_557, w_002_558, w_002_559, w_002_560, w_002_561, w_002_562, w_002_563, w_002_564, w_002_565, w_002_566, w_002_567, w_002_568, w_002_569, w_002_570, w_002_571, w_002_572, w_002_573, w_002_574, w_002_575, w_002_576, w_002_577, w_002_578, w_002_579, w_002_580, w_002_581, w_002_582, w_002_583, w_002_584, w_002_585, w_002_586, w_002_587, w_002_588, w_002_589, w_002_590, w_002_591, w_002_592, w_002_593;
  wire w_003_000, w_003_001, w_003_002, w_003_003, w_003_004, w_003_005, w_003_006, w_003_007, w_003_008, w_003_009, w_003_010, w_003_011, w_003_012, w_003_013, w_003_014, w_003_015, w_003_016, w_003_017, w_003_018, w_003_019, w_003_020, w_003_021, w_003_022, w_003_023, w_003_024, w_003_025, w_003_026, w_003_027, w_003_028, w_003_029, w_003_030, w_003_031, w_003_032, w_003_033, w_003_034, w_003_035, w_003_036, w_003_037, w_003_038, w_003_039, w_003_040, w_003_041, w_003_042, w_003_043, w_003_044, w_003_045, w_003_046, w_003_047, w_003_048, w_003_049, w_003_050, w_003_051, w_003_052, w_003_053, w_003_054, w_003_055, w_003_056, w_003_057, w_003_058, w_003_059, w_003_060, w_003_061, w_003_062, w_003_063, w_003_064, w_003_065, w_003_066, w_003_067, w_003_068, w_003_069, w_003_070, w_003_071, w_003_072, w_003_073, w_003_074, w_003_075, w_003_076, w_003_077, w_003_078, w_003_079, w_003_080, w_003_081, w_003_082, w_003_083, w_003_084, w_003_085, w_003_086, w_003_087, w_003_088, w_003_089, w_003_090, w_003_091, w_003_092, w_003_093, w_003_094, w_003_095, w_003_096, w_003_097, w_003_098, w_003_099, w_003_100, w_003_101, w_003_102, w_003_103, w_003_104, w_003_105, w_003_106, w_003_107, w_003_108, w_003_109, w_003_110, w_003_111, w_003_112, w_003_113, w_003_114, w_003_115, w_003_116, w_003_117, w_003_118, w_003_119, w_003_120, w_003_121, w_003_122, w_003_123, w_003_124, w_003_125, w_003_126, w_003_127, w_003_128, w_003_129, w_003_130, w_003_131, w_003_132, w_003_133, w_003_134, w_003_135, w_003_136, w_003_137, w_003_138, w_003_139, w_003_140, w_003_141, w_003_142, w_003_143, w_003_144, w_003_145, w_003_147, w_003_148, w_003_149, w_003_150, w_003_151, w_003_152, w_003_153, w_003_154, w_003_155, w_003_156, w_003_157, w_003_158, w_003_159, w_003_160, w_003_161, w_003_162, w_003_163, w_003_164, w_003_165, w_003_166, w_003_167, w_003_168, w_003_169, w_003_170, w_003_171, w_003_172, w_003_173, w_003_174, w_003_175, w_003_176, w_003_177, w_003_178, w_003_179, w_003_180, w_003_181, w_003_182, w_003_183, w_003_184, w_003_185, w_003_186, w_003_187, w_003_188, w_003_189, w_003_190, w_003_191, w_003_192, w_003_193, w_003_194, w_003_195, w_003_196, w_003_197, w_003_198, w_003_199, w_003_200, w_003_201, w_003_202, w_003_203, w_003_204, w_003_205, w_003_206, w_003_207, w_003_208, w_003_209, w_003_210, w_003_211, w_003_212, w_003_213, w_003_214, w_003_215, w_003_216, w_003_217, w_003_218, w_003_219, w_003_220, w_003_221, w_003_222, w_003_223, w_003_224, w_003_225, w_003_226, w_003_227, w_003_228, w_003_229, w_003_230, w_003_231, w_003_232, w_003_233, w_003_234, w_003_235, w_003_236, w_003_237, w_003_238, w_003_239, w_003_240, w_003_241, w_003_242, w_003_243, w_003_244, w_003_245, w_003_246, w_003_247, w_003_248, w_003_249, w_003_250, w_003_251, w_003_252, w_003_253, w_003_254, w_003_255, w_003_256, w_003_257, w_003_258, w_003_259, w_003_260, w_003_261, w_003_262, w_003_263, w_003_264, w_003_265, w_003_266, w_003_267, w_003_268, w_003_269, w_003_270, w_003_271, w_003_272, w_003_273, w_003_274, w_003_275, w_003_276, w_003_277, w_003_278, w_003_279, w_003_280, w_003_281, w_003_282, w_003_283, w_003_284, w_003_285, w_003_286, w_003_287, w_003_288, w_003_289, w_003_290, w_003_291, w_003_292, w_003_293, w_003_294, w_003_295, w_003_296, w_003_297, w_003_298, w_003_299, w_003_300, w_003_301, w_003_302, w_003_303, w_003_304, w_003_305, w_003_306, w_003_307, w_003_308, w_003_309, w_003_310, w_003_311, w_003_312, w_003_313, w_003_314, w_003_315, w_003_316, w_003_317, w_003_318, w_003_319;
  wire w_004_000, w_004_001, w_004_002, w_004_003, w_004_004, w_004_005, w_004_007, w_004_008, w_004_009, w_004_011, w_004_012, w_004_013, w_004_014, w_004_015, w_004_016, w_004_017, w_004_019, w_004_021, w_004_022, w_004_024, w_004_025, w_004_027, w_004_028, w_004_029, w_004_030, w_004_031, w_004_032, w_004_035, w_004_036, w_004_039, w_004_041, w_004_042, w_004_043, w_004_044, w_004_045, w_004_046, w_004_047, w_004_048, w_004_049, w_004_050, w_004_051, w_004_054, w_004_056, w_004_057, w_004_058, w_004_059, w_004_060, w_004_061, w_004_062, w_004_063, w_004_064, w_004_066, w_004_068, w_004_070, w_004_071, w_004_074, w_004_075, w_004_076, w_004_077, w_004_078, w_004_079, w_004_080, w_004_081, w_004_082, w_004_084, w_004_085, w_004_086, w_004_087, w_004_088, w_004_091, w_004_093, w_004_095, w_004_096, w_004_100, w_004_101, w_004_102, w_004_104, w_004_107, w_004_108, w_004_109, w_004_111, w_004_112, w_004_114, w_004_115, w_004_116, w_004_117, w_004_118, w_004_120, w_004_121, w_004_122, w_004_123, w_004_126, w_004_130, w_004_132, w_004_134, w_004_135, w_004_136, w_004_137, w_004_139, w_004_141, w_004_142, w_004_143, w_004_144, w_004_146, w_004_147, w_004_148, w_004_151, w_004_152, w_004_153, w_004_156, w_004_157, w_004_159, w_004_160, w_004_162, w_004_166, w_004_167, w_004_170, w_004_171, w_004_172, w_004_173, w_004_175, w_004_176, w_004_177, w_004_179, w_004_181, w_004_182, w_004_183, w_004_185, w_004_186, w_004_187, w_004_188, w_004_190, w_004_191, w_004_192, w_004_194, w_004_195, w_004_196, w_004_197, w_004_199, w_004_200, w_004_201, w_004_202, w_004_206, w_004_207, w_004_209, w_004_210, w_004_211, w_004_213, w_004_214, w_004_215, w_004_216, w_004_217, w_004_218, w_004_220, w_004_222, w_004_223, w_004_225, w_004_226, w_004_227, w_004_229, w_004_232, w_004_233, w_004_234, w_004_235, w_004_236, w_004_241, w_004_243, w_004_245, w_004_246, w_004_248, w_004_249, w_004_250, w_004_251, w_004_252, w_004_254, w_004_257, w_004_258, w_004_259, w_004_260, w_004_261, w_004_262, w_004_264, w_004_265, w_004_266, w_004_269, w_004_275, w_004_276, w_004_277, w_004_278, w_004_279, w_004_280, w_004_283, w_004_286, w_004_288, w_004_292, w_004_293, w_004_296, w_004_298, w_004_300, w_004_301, w_004_303, w_004_305, w_004_307, w_004_310, w_004_312, w_004_313, w_004_314, w_004_315, w_004_316, w_004_318, w_004_319, w_004_321, w_004_322, w_004_323, w_004_324, w_004_325, w_004_326, w_004_328, w_004_331, w_004_334, w_004_337, w_004_340, w_004_342, w_004_343, w_004_345, w_004_346, w_004_352, w_004_353, w_004_355, w_004_356, w_004_359, w_004_361, w_004_362, w_004_364, w_004_366, w_004_368, w_004_369, w_004_371, w_004_372, w_004_373, w_004_374, w_004_375, w_004_377, w_004_379, w_004_380, w_004_382, w_004_383, w_004_384, w_004_385, w_004_388, w_004_391, w_004_394, w_004_395, w_004_396, w_004_398, w_004_399, w_004_400, w_004_402, w_004_404, w_004_406, w_004_407, w_004_409, w_004_415, w_004_416, w_004_417, w_004_418, w_004_420, w_004_422, w_004_425, w_004_428, w_004_429, w_004_430, w_004_433, w_004_435, w_004_436, w_004_437, w_004_443, w_004_444, w_004_445, w_004_446, w_004_447, w_004_448, w_004_449, w_004_451, w_004_452, w_004_453, w_004_454, w_004_458, w_004_459, w_004_460, w_004_462, w_004_469, w_004_472, w_004_476, w_004_477, w_004_478, w_004_481, w_004_482, w_004_483, w_004_486, w_004_487, w_004_488, w_004_490, w_004_491, w_004_492, w_004_493, w_004_494, w_004_496, w_004_498, w_004_501, w_004_503, w_004_504, w_004_506, w_004_507, w_004_510, w_004_512, w_004_513, w_004_514, w_004_515, w_004_516, w_004_517, w_004_518, w_004_520, w_004_524, w_004_527, w_004_528, w_004_529, w_004_530, w_004_534, w_004_535, w_004_537, w_004_538, w_004_540, w_004_543, w_004_544, w_004_545, w_004_546, w_004_547, w_004_548, w_004_550, w_004_551, w_004_552, w_004_553, w_004_554, w_004_555, w_004_558, w_004_560, w_004_561, w_004_562, w_004_563, w_004_565, w_004_566, w_004_571, w_004_575, w_004_576, w_004_579, w_004_581, w_004_583, w_004_584, w_004_585, w_004_587, w_004_588, w_004_590, w_004_591, w_004_592, w_004_593, w_004_595, w_004_596, w_004_597, w_004_598, w_004_599, w_004_602, w_004_603, w_004_604, w_004_605, w_004_606, w_004_607, w_004_609, w_004_610, w_004_611, w_004_615, w_004_616, w_004_617, w_004_618, w_004_620, w_004_624, w_004_625, w_004_626, w_004_628, w_004_633, w_004_635, w_004_636, w_004_637, w_004_638, w_004_639, w_004_640, w_004_641, w_004_642, w_004_644, w_004_645, w_004_646, w_004_652, w_004_653, w_004_655, w_004_656, w_004_657, w_004_659, w_004_661, w_004_663, w_004_664, w_004_665, w_004_670, w_004_671, w_004_672, w_004_677, w_004_678, w_004_680, w_004_683, w_004_687, w_004_694, w_004_695, w_004_697, w_004_700, w_004_701, w_004_703, w_004_704, w_004_705, w_004_706, w_004_710, w_004_711, w_004_713, w_004_714, w_004_715, w_004_717, w_004_719, w_004_721, w_004_722, w_004_723, w_004_724, w_004_725, w_004_726, w_004_727, w_004_730, w_004_731, w_004_732, w_004_733, w_004_737, w_004_738, w_004_739, w_004_743, w_004_744, w_004_746, w_004_749, w_004_750, w_004_753, w_004_754, w_004_755, w_004_756, w_004_757, w_004_758, w_004_762, w_004_764, w_004_765, w_004_766, w_004_768, w_004_769, w_004_770, w_004_771, w_004_772, w_004_774, w_004_775, w_004_777, w_004_778, w_004_780, w_004_782, w_004_783, w_004_785, w_004_787, w_004_788, w_004_790, w_004_796, w_004_797, w_004_798, w_004_799, w_004_803, w_004_804, w_004_805, w_004_807, w_004_809, w_004_810, w_004_813, w_004_814, w_004_815, w_004_816, w_004_817, w_004_818, w_004_819, w_004_823, w_004_824, w_004_826, w_004_827, w_004_828, w_004_830, w_004_831, w_004_832, w_004_834, w_004_836, w_004_837, w_004_838, w_004_839, w_004_840, w_004_841, w_004_842, w_004_843, w_004_846, w_004_848, w_004_850, w_004_852, w_004_853, w_004_854, w_004_856, w_004_860, w_004_862, w_004_866, w_004_868, w_004_870, w_004_871, w_004_872, w_004_876, w_004_877, w_004_878, w_004_879, w_004_881, w_004_884, w_004_885, w_004_886, w_004_888, w_004_890, w_004_892, w_004_894, w_004_895, w_004_896, w_004_897, w_004_898, w_004_899, w_004_900, w_004_901, w_004_904, w_004_905, w_004_907, w_004_908, w_004_909, w_004_910, w_004_912, w_004_914, w_004_916, w_004_917, w_004_918, w_004_920, w_004_921, w_004_922, w_004_925, w_004_926, w_004_929, w_004_931, w_004_933, w_004_934, w_004_935, w_004_937, w_004_938, w_004_941, w_004_942, w_004_943, w_004_949, w_004_950, w_004_952, w_004_953, w_004_955, w_004_957, w_004_958, w_004_959, w_004_960, w_004_962, w_004_963, w_004_964, w_004_970, w_004_973, w_004_975, w_004_977, w_004_978, w_004_979, w_004_980, w_004_981, w_004_983, w_004_984, w_004_985, w_004_987, w_004_989, w_004_990, w_004_991, w_004_993, w_004_994, w_004_996, w_004_997, w_004_1001, w_004_1004, w_004_1008, w_004_1009, w_004_1011, w_004_1015, w_004_1016, w_004_1017, w_004_1020, w_004_1021, w_004_1023, w_004_1025, w_004_1027, w_004_1028, w_004_1029, w_004_1030, w_004_1033, w_004_1035, w_004_1037, w_004_1038, w_004_1039, w_004_1040, w_004_1043, w_004_1046, w_004_1047, w_004_1049, w_004_1050, w_004_1051, w_004_1053, w_004_1054, w_004_1056, w_004_1061, w_004_1062, w_004_1063, w_004_1065, w_004_1066, w_004_1069, w_004_1071, w_004_1073, w_004_1074, w_004_1076, w_004_1077, w_004_1078, w_004_1080, w_004_1082, w_004_1083, w_004_1085, w_004_1086, w_004_1089, w_004_1090, w_004_1091, w_004_1092, w_004_1093, w_004_1094, w_004_1095, w_004_1096, w_004_1097, w_004_1098, w_004_1100, w_004_1101, w_004_1102, w_004_1105, w_004_1107, w_004_1108, w_004_1109, w_004_1110, w_004_1111, w_004_1112, w_004_1114, w_004_1115, w_004_1116, w_004_1120, w_004_1121, w_004_1122, w_004_1123, w_004_1125, w_004_1127, w_004_1128, w_004_1130, w_004_1132, w_004_1133, w_004_1135, w_004_1136, w_004_1138, w_004_1140, w_004_1141, w_004_1149, w_004_1150, w_004_1151, w_004_1152, w_004_1153, w_004_1157, w_004_1158, w_004_1161, w_004_1164, w_004_1166, w_004_1169, w_004_1171, w_004_1174, w_004_1177, w_004_1179, w_004_1180, w_004_1181, w_004_1182, w_004_1184, w_004_1186, w_004_1187, w_004_1188, w_004_1189, w_004_1191, w_004_1194, w_004_1197, w_004_1200, w_004_1201, w_004_1202, w_004_1204, w_004_1206, w_004_1207, w_004_1208, w_004_1210, w_004_1211, w_004_1212, w_004_1215, w_004_1216, w_004_1217, w_004_1221, w_004_1222, w_004_1224, w_004_1226, w_004_1228, w_004_1229, w_004_1231, w_004_1232, w_004_1234, w_004_1235, w_004_1236, w_004_1239, w_004_1241, w_004_1243, w_004_1244, w_004_1248, w_004_1250, w_004_1254, w_004_1255, w_004_1259, w_004_1260, w_004_1263, w_004_1264, w_004_1265, w_004_1267, w_004_1268, w_004_1269, w_004_1270, w_004_1271, w_004_1272, w_004_1276, w_004_1278, w_004_1279, w_004_1280, w_004_1281, w_004_1283, w_004_1284, w_004_1287, w_004_1288, w_004_1289, w_004_1290, w_004_1291, w_004_1292, w_004_1293, w_004_1294, w_004_1295, w_004_1296, w_004_1298, w_004_1300, w_004_1301, w_004_1302, w_004_1305, w_004_1306, w_004_1310, w_004_1311, w_004_1312, w_004_1315, w_004_1319, w_004_1320, w_004_1321, w_004_1322, w_004_1324, w_004_1326, w_004_1328, w_004_1329, w_004_1330, w_004_1335, w_004_1337, w_004_1338, w_004_1340, w_004_1344, w_004_1348, w_004_1349, w_004_1352, w_004_1354, w_004_1356, w_004_1357, w_004_1358, w_004_1361, w_004_1362, w_004_1364, w_004_1365, w_004_1366, w_004_1374, w_004_1379, w_004_1380, w_004_1381, w_004_1382, w_004_1384, w_004_1388, w_004_1390, w_004_1393, w_004_1394, w_004_1398, w_004_1399, w_004_1401, w_004_1402, w_004_1404, w_004_1406, w_004_1409, w_004_1410, w_004_1412, w_004_1413, w_004_1414, w_004_1415, w_004_1417, w_004_1418, w_004_1420, w_004_1422, w_004_1423, w_004_1425, w_004_1427, w_004_1428, w_004_1430, w_004_1435, w_004_1436, w_004_1437, w_004_1442, w_004_1445, w_004_1446, w_004_1447, w_004_1448, w_004_1449, w_004_1453, w_004_1454, w_004_1455, w_004_1456, w_004_1458, w_004_1459, w_004_1460, w_004_1463, w_004_1466, w_004_1467, w_004_1468, w_004_1469, w_004_1470, w_004_1472, w_004_1474, w_004_1478, w_004_1480, w_004_1481, w_004_1484, w_004_1485, w_004_1487, w_004_1488, w_004_1492, w_004_1493, w_004_1494, w_004_1495, w_004_1501, w_004_1502, w_004_1508, w_004_1509, w_004_1511, w_004_1516, w_004_1517, w_004_1519, w_004_1521, w_004_1523, w_004_1524, w_004_1530, w_004_1532, w_004_1533, w_004_1534, w_004_1535, w_004_1537, w_004_1539, w_004_1540, w_004_1543, w_004_1544, w_004_1546, w_004_1547, w_004_1549, w_004_1552, w_004_1553, w_004_1554, w_004_1555, w_004_1558, w_004_1560, w_004_1562, w_004_1563, w_004_1565, w_004_1566, w_004_1568, w_004_1570, w_004_1572, w_004_1573, w_004_1575, w_004_1576, w_004_1578, w_004_1583, w_004_1589, w_004_1590, w_004_1592, w_004_1593, w_004_1594, w_004_1595, w_004_1596, w_004_1597, w_004_1599, w_004_1600, w_004_1601, w_004_1602, w_004_1603, w_004_1604, w_004_1605, w_004_1608, w_004_1610, w_004_1611, w_004_1612, w_004_1613, w_004_1614, w_004_1615, w_004_1616, w_004_1618, w_004_1619, w_004_1622, w_004_1624, w_004_1625, w_004_1626, w_004_1631, w_004_1633, w_004_1635, w_004_1636, w_004_1637, w_004_1638, w_004_1640, w_004_1641, w_004_1643, w_004_1645, w_004_1647, w_004_1648, w_004_1649, w_004_1652, w_004_1653, w_004_1655, w_004_1656, w_004_1659, w_004_1660, w_004_1661, w_004_1663, w_004_1664, w_004_1665, w_004_1667, w_004_1674, w_004_1675, w_004_1678, w_004_1679, w_004_1681, w_004_1682, w_004_1684, w_004_1686, w_004_1687, w_004_1689, w_004_1690, w_004_1692, w_004_1693, w_004_1694, w_004_1696, w_004_1698, w_004_1699, w_004_1702, w_004_1703, w_004_1706, w_004_1707, w_004_1708, w_004_1709, w_004_1711, w_004_1712, w_004_1714, w_004_1716, w_004_1718, w_004_1719, w_004_1720, w_004_1727, w_004_1731, w_004_1732, w_004_1733, w_004_1734, w_004_1737, w_004_1739, w_004_1740, w_004_1741, w_004_1742, w_004_1743, w_004_1744, w_004_1745, w_004_1746, w_004_1747, w_004_1748, w_004_1749, w_004_1750, w_004_1752, w_004_1753, w_004_1755, w_004_1756, w_004_1757, w_004_1760, w_004_1765, w_004_1767, w_004_1769, w_004_1770, w_004_1771, w_004_1773, w_004_1774, w_004_1776, w_004_1777, w_004_1778, w_004_1780, w_004_1781, w_004_1782, w_004_1784, w_004_1786, w_004_1787, w_004_1788, w_004_1791, w_004_1792, w_004_1793, w_004_1795, w_004_1797, w_004_1798, w_004_1799, w_004_1800, w_004_1801, w_004_1802, w_004_1805, w_004_1807, w_004_1809, w_004_1810, w_004_1811, w_004_1812, w_004_1814, w_004_1815, w_004_1817, w_004_1819, w_004_1821, w_004_1823, w_004_1827, w_004_1828, w_004_1829, w_004_1831, w_004_1832, w_004_1833, w_004_1834, w_004_1835, w_004_1836, w_004_1837, w_004_1839, w_004_1840, w_004_1841, w_004_1843, w_004_1845, w_004_1848, w_004_1849, w_004_1850, w_004_1851, w_004_1852, w_004_1855, w_004_1858, w_004_1860, w_004_1861, w_004_1863, w_004_1864, w_004_1865, w_004_1867, w_004_1868, w_004_1871, w_004_1872, w_004_1873, w_004_1874, w_004_1875, w_004_1882, w_004_1883, w_004_1884, w_004_1885, w_004_1886, w_004_1887, w_004_1888, w_004_1893, w_004_1894, w_004_1895, w_004_1896, w_004_1899, w_004_1900, w_004_1902, w_004_1905, w_004_1906, w_004_1907, w_004_1909, w_004_1910, w_004_1911;
  wire w_005_001, w_005_003, w_005_004, w_005_005, w_005_006, w_005_008, w_005_009, w_005_013, w_005_014, w_005_015, w_005_016, w_005_017, w_005_019, w_005_021, w_005_022, w_005_023, w_005_024, w_005_025, w_005_026, w_005_029, w_005_030, w_005_032, w_005_033, w_005_034, w_005_035, w_005_036, w_005_037, w_005_038, w_005_039, w_005_040, w_005_041, w_005_042, w_005_044, w_005_045, w_005_046, w_005_047, w_005_048, w_005_049, w_005_050, w_005_051, w_005_052, w_005_053, w_005_054, w_005_055, w_005_056, w_005_057, w_005_058, w_005_059, w_005_060, w_005_065, w_005_066, w_005_068, w_005_069, w_005_070, w_005_072, w_005_073, w_005_074, w_005_075, w_005_076, w_005_077, w_005_078, w_005_079, w_005_080, w_005_082, w_005_083, w_005_084, w_005_086, w_005_087, w_005_089, w_005_090, w_005_093, w_005_094, w_005_095, w_005_096, w_005_097, w_005_098, w_005_100, w_005_101, w_005_103, w_005_105, w_005_106, w_005_109, w_005_111, w_005_112, w_005_114, w_005_115, w_005_116, w_005_117, w_005_120, w_005_121, w_005_123, w_005_124, w_005_125, w_005_126, w_005_127, w_005_128, w_005_129, w_005_131, w_005_132, w_005_133, w_005_134, w_005_136, w_005_137, w_005_139, w_005_140, w_005_142, w_005_143, w_005_144, w_005_146, w_005_148, w_005_149, w_005_150, w_005_151, w_005_152, w_005_153, w_005_154, w_005_155, w_005_156, w_005_158, w_005_159, w_005_160, w_005_162, w_005_163, w_005_165, w_005_167, w_005_168, w_005_169, w_005_170, w_005_172, w_005_173, w_005_175, w_005_176, w_005_178, w_005_179, w_005_180, w_005_182, w_005_183, w_005_186, w_005_187, w_005_188, w_005_189, w_005_190, w_005_191, w_005_192, w_005_194, w_005_195, w_005_196, w_005_197, w_005_199, w_005_201, w_005_202, w_005_203, w_005_204, w_005_205, w_005_206, w_005_207, w_005_208, w_005_209, w_005_212, w_005_213, w_005_216, w_005_220, w_005_222, w_005_223, w_005_226, w_005_228, w_005_229, w_005_232, w_005_234, w_005_236, w_005_237, w_005_239, w_005_240, w_005_242, w_005_243, w_005_244, w_005_245, w_005_246, w_005_248, w_005_251, w_005_252, w_005_253, w_005_255, w_005_256, w_005_257, w_005_258, w_005_259, w_005_260, w_005_261, w_005_262, w_005_263, w_005_267, w_005_268, w_005_269, w_005_271, w_005_272, w_005_273, w_005_274, w_005_275, w_005_276, w_005_278, w_005_279, w_005_280, w_005_281, w_005_283, w_005_285, w_005_286, w_005_287, w_005_288, w_005_289, w_005_290, w_005_292, w_005_293, w_005_294, w_005_295, w_005_296, w_005_298, w_005_299, w_005_300, w_005_302, w_005_303, w_005_305, w_005_306, w_005_307, w_005_308, w_005_309, w_005_310, w_005_313, w_005_314, w_005_315, w_005_316, w_005_317, w_005_318, w_005_319, w_005_320, w_005_321, w_005_322, w_005_323, w_005_328, w_005_331, w_005_333, w_005_338, w_005_339, w_005_341, w_005_344, w_005_346, w_005_348, w_005_357, w_005_362, w_005_363, w_005_366, w_005_368, w_005_369, w_005_371, w_005_375, w_005_376, w_005_377, w_005_378, w_005_379, w_005_381, w_005_385, w_005_386, w_005_387, w_005_390, w_005_394, w_005_395, w_005_398, w_005_400, w_005_402, w_005_406, w_005_408, w_005_409, w_005_411, w_005_415, w_005_420, w_005_423, w_005_425, w_005_428, w_005_430, w_005_433, w_005_434, w_005_438, w_005_439, w_005_444, w_005_446, w_005_449, w_005_453, w_005_457, w_005_458, w_005_459, w_005_460, w_005_461, w_005_465, w_005_466, w_005_472, w_005_473, w_005_477, w_005_478, w_005_479, w_005_484, w_005_485, w_005_487, w_005_488, w_005_490, w_005_494, w_005_496, w_005_497, w_005_500, w_005_501, w_005_503, w_005_504, w_005_505, w_005_506, w_005_508, w_005_511, w_005_523, w_005_525, w_005_527, w_005_528, w_005_529, w_005_530, w_005_532, w_005_533, w_005_534, w_005_535, w_005_537, w_005_538, w_005_539, w_005_541, w_005_542, w_005_543, w_005_544, w_005_546, w_005_548, w_005_551, w_005_555, w_005_556, w_005_559, w_005_560, w_005_562, w_005_564, w_005_565, w_005_570, w_005_574, w_005_576, w_005_577, w_005_578, w_005_580, w_005_584, w_005_585, w_005_586, w_005_591, w_005_593, w_005_594, w_005_596, w_005_597, w_005_598, w_005_599, w_005_600, w_005_602, w_005_605, w_005_608, w_005_610, w_005_611, w_005_612, w_005_617, w_005_619, w_005_620, w_005_622, w_005_623, w_005_624, w_005_625, w_005_627, w_005_628, w_005_630, w_005_632, w_005_633, w_005_636, w_005_638, w_005_640, w_005_642, w_005_643, w_005_644, w_005_645, w_005_647, w_005_650, w_005_651, w_005_652, w_005_653, w_005_654, w_005_655, w_005_658, w_005_659, w_005_661, w_005_662, w_005_663, w_005_665, w_005_668, w_005_669, w_005_670, w_005_671, w_005_672, w_005_673, w_005_674, w_005_675, w_005_677, w_005_680, w_005_682, w_005_686, w_005_687, w_005_694, w_005_695, w_005_697, w_005_699, w_005_702, w_005_706, w_005_707, w_005_708, w_005_709, w_005_712, w_005_713, w_005_717, w_005_722, w_005_728, w_005_729, w_005_730, w_005_731, w_005_732, w_005_733, w_005_734, w_005_736, w_005_738, w_005_741, w_005_742, w_005_747, w_005_748, w_005_752, w_005_753, w_005_756, w_005_758, w_005_759, w_005_760, w_005_765, w_005_766, w_005_768, w_005_769, w_005_770, w_005_771, w_005_774, w_005_775, w_005_777, w_005_778, w_005_780, w_005_781, w_005_782, w_005_785, w_005_786, w_005_787, w_005_789, w_005_790, w_005_791, w_005_793, w_005_794, w_005_796, w_005_797, w_005_798, w_005_800, w_005_801, w_005_802, w_005_808, w_005_809, w_005_811, w_005_812, w_005_816, w_005_817, w_005_823, w_005_824, w_005_825, w_005_830, w_005_832, w_005_838, w_005_839, w_005_840, w_005_841, w_005_842, w_005_844, w_005_845, w_005_849, w_005_850, w_005_851, w_005_853, w_005_856, w_005_857, w_005_858, w_005_860, w_005_862, w_005_863, w_005_864, w_005_872, w_005_873, w_005_875, w_005_876, w_005_880, w_005_882, w_005_883, w_005_886, w_005_890, w_005_891, w_005_893, w_005_894, w_005_897, w_005_898, w_005_901, w_005_905, w_005_907, w_005_910, w_005_911, w_005_912, w_005_914, w_005_915, w_005_917, w_005_919, w_005_922, w_005_924, w_005_926, w_005_929, w_005_930, w_005_932, w_005_933, w_005_934, w_005_937, w_005_943, w_005_944, w_005_949, w_005_951, w_005_952, w_005_953, w_005_954, w_005_955, w_005_959, w_005_960, w_005_961, w_005_962, w_005_965, w_005_966, w_005_967, w_005_970, w_005_971, w_005_973, w_005_974, w_005_975, w_005_977, w_005_979, w_005_982, w_005_984, w_005_986, w_005_988, w_005_993, w_005_994, w_005_995, w_005_997, w_005_999, w_005_1002, w_005_1005, w_005_1006, w_005_1007, w_005_1010, w_005_1011, w_005_1015, w_005_1019, w_005_1022, w_005_1023, w_005_1025, w_005_1026, w_005_1027, w_005_1028, w_005_1033, w_005_1034, w_005_1035, w_005_1038, w_005_1041, w_005_1043, w_005_1044, w_005_1045, w_005_1047, w_005_1050, w_005_1052, w_005_1056, w_005_1057, w_005_1058, w_005_1059, w_005_1061, w_005_1065, w_005_1070, w_005_1074, w_005_1075, w_005_1076, w_005_1077, w_005_1078, w_005_1079, w_005_1080, w_005_1081, w_005_1082, w_005_1087, w_005_1088, w_005_1090, w_005_1092, w_005_1093, w_005_1094, w_005_1098, w_005_1099, w_005_1100, w_005_1101, w_005_1102, w_005_1103, w_005_1105, w_005_1106, w_005_1109, w_005_1112, w_005_1113, w_005_1114, w_005_1115, w_005_1116, w_005_1117, w_005_1118, w_005_1119, w_005_1121, w_005_1123, w_005_1125, w_005_1126, w_005_1129, w_005_1130, w_005_1132, w_005_1133, w_005_1134, w_005_1136, w_005_1137, w_005_1138, w_005_1139, w_005_1140, w_005_1141, w_005_1142, w_005_1143, w_005_1147, w_005_1149, w_005_1150, w_005_1151, w_005_1152, w_005_1153, w_005_1157, w_005_1158, w_005_1159, w_005_1160, w_005_1163, w_005_1165, w_005_1166, w_005_1167, w_005_1168, w_005_1171, w_005_1173, w_005_1175, w_005_1178, w_005_1180, w_005_1181, w_005_1182, w_005_1185, w_005_1186, w_005_1187, w_005_1189, w_005_1190, w_005_1197, w_005_1199, w_005_1205, w_005_1209, w_005_1211, w_005_1213, w_005_1216, w_005_1217, w_005_1218, w_005_1219, w_005_1220, w_005_1222, w_005_1223, w_005_1224, w_005_1228, w_005_1229, w_005_1233, w_005_1234, w_005_1235, w_005_1237, w_005_1239, w_005_1243, w_005_1251, w_005_1252, w_005_1254, w_005_1255, w_005_1257, w_005_1258, w_005_1259, w_005_1261, w_005_1264, w_005_1265, w_005_1266, w_005_1267, w_005_1268, w_005_1271, w_005_1274, w_005_1276, w_005_1278, w_005_1281, w_005_1283, w_005_1285, w_005_1286, w_005_1288, w_005_1289, w_005_1292, w_005_1293, w_005_1296, w_005_1297, w_005_1298, w_005_1300, w_005_1303, w_005_1304, w_005_1307, w_005_1308, w_005_1309, w_005_1310, w_005_1315, w_005_1317, w_005_1321, w_005_1322, w_005_1324, w_005_1328, w_005_1329, w_005_1330, w_005_1331, w_005_1336, w_005_1337, w_005_1346, w_005_1347, w_005_1348, w_005_1349, w_005_1353, w_005_1355, w_005_1357, w_005_1358, w_005_1360, w_005_1362, w_005_1364, w_005_1366, w_005_1368, w_005_1369, w_005_1370, w_005_1374, w_005_1376, w_005_1379, w_005_1380, w_005_1381, w_005_1384, w_005_1385, w_005_1392, w_005_1393, w_005_1394, w_005_1397, w_005_1398, w_005_1404, w_005_1408, w_005_1409, w_005_1410, w_005_1415, w_005_1418, w_005_1420, w_005_1421, w_005_1422, w_005_1424, w_005_1426, w_005_1428, w_005_1429, w_005_1430, w_005_1431, w_005_1436, w_005_1439, w_005_1440, w_005_1441, w_005_1443, w_005_1445, w_005_1446, w_005_1447, w_005_1448, w_005_1449, w_005_1450, w_005_1451, w_005_1461, w_005_1464, w_005_1467, w_005_1469, w_005_1470, w_005_1473, w_005_1478, w_005_1480, w_005_1485, w_005_1487, w_005_1491, w_005_1492, w_005_1493, w_005_1494, w_005_1495, w_005_1499, w_005_1501, w_005_1505, w_005_1511, w_005_1513, w_005_1519, w_005_1522, w_005_1523, w_005_1525, w_005_1526, w_005_1528, w_005_1529, w_005_1533, w_005_1534, w_005_1536, w_005_1538, w_005_1540, w_005_1542, w_005_1548, w_005_1549, w_005_1550, w_005_1551, w_005_1553, w_005_1554, w_005_1557, w_005_1558, w_005_1560, w_005_1561, w_005_1562, w_005_1566, w_005_1569, w_005_1572, w_005_1574, w_005_1575, w_005_1576, w_005_1577, w_005_1579, w_005_1580, w_005_1581, w_005_1582, w_005_1584, w_005_1587, w_005_1588, w_005_1591, w_005_1592, w_005_1593, w_005_1596, w_005_1597, w_005_1602, w_005_1603, w_005_1605, w_005_1609, w_005_1610, w_005_1612, w_005_1613, w_005_1616, w_005_1617, w_005_1619, w_005_1620, w_005_1622, w_005_1624, w_005_1626, w_005_1628, w_005_1631, w_005_1636, w_005_1637, w_005_1638, w_005_1639, w_005_1641, w_005_1645, w_005_1646, w_005_1650, w_005_1651, w_005_1652, w_005_1653, w_005_1656, w_005_1658, w_005_1662, w_005_1663, w_005_1664, w_005_1666, w_005_1667, w_005_1668, w_005_1669, w_005_1672, w_005_1674;
  wire w_006_000, w_006_001, w_006_002, w_006_003, w_006_004, w_006_005, w_006_006, w_006_007, w_006_008, w_006_009, w_006_010, w_006_011, w_006_012, w_006_013, w_006_014, w_006_015, w_006_017, w_006_018, w_006_019, w_006_020, w_006_021, w_006_022, w_006_023, w_006_024, w_006_025, w_006_026, w_006_027, w_006_028, w_006_029, w_006_030, w_006_031, w_006_032, w_006_033, w_006_034, w_006_035, w_006_036, w_006_038, w_006_039, w_006_040, w_006_041, w_006_042, w_006_043, w_006_044, w_006_045, w_006_046, w_006_047, w_006_048, w_006_049, w_006_050, w_006_051, w_006_052, w_006_053, w_006_054, w_006_055, w_006_056, w_006_057, w_006_058, w_006_059, w_006_060, w_006_061, w_006_062, w_006_063, w_006_064, w_006_065, w_006_066, w_006_067, w_006_068, w_006_069, w_006_070, w_006_071, w_006_072, w_006_073, w_006_074, w_006_075, w_006_076, w_006_077, w_006_078, w_006_079, w_006_080, w_006_081, w_006_082, w_006_083, w_006_084, w_006_085, w_006_086, w_006_087, w_006_088, w_006_089, w_006_090, w_006_091, w_006_092, w_006_093, w_006_094, w_006_095, w_006_096, w_006_097, w_006_098, w_006_099, w_006_100, w_006_101, w_006_102, w_006_103, w_006_104, w_006_105, w_006_106, w_006_107, w_006_108, w_006_109, w_006_110, w_006_111, w_006_112, w_006_113, w_006_114, w_006_115, w_006_116, w_006_117, w_006_118, w_006_119, w_006_120, w_006_121, w_006_122, w_006_123, w_006_124, w_006_125, w_006_126, w_006_127, w_006_128, w_006_129, w_006_130, w_006_131, w_006_132, w_006_133, w_006_134, w_006_135, w_006_137, w_006_138, w_006_139, w_006_140, w_006_141, w_006_142, w_006_143, w_006_144, w_006_145, w_006_146, w_006_147, w_006_148, w_006_149, w_006_150, w_006_151, w_006_152, w_006_153, w_006_154, w_006_155, w_006_156, w_006_157, w_006_158, w_006_159, w_006_160, w_006_161, w_006_162, w_006_163, w_006_164, w_006_165, w_006_166, w_006_167, w_006_168, w_006_169, w_006_170, w_006_171, w_006_172, w_006_173, w_006_174, w_006_175, w_006_176, w_006_177, w_006_178, w_006_179, w_006_180, w_006_182, w_006_183, w_006_184, w_006_185, w_006_186, w_006_187, w_006_188, w_006_189, w_006_190, w_006_191, w_006_192, w_006_193, w_006_194, w_006_195, w_006_196, w_006_197, w_006_198, w_006_199, w_006_200, w_006_201, w_006_202, w_006_203, w_006_204, w_006_205, w_006_206, w_006_207, w_006_208, w_006_209, w_006_210, w_006_211, w_006_212, w_006_214, w_006_215, w_006_216, w_006_217, w_006_218, w_006_219, w_006_220, w_006_221, w_006_222, w_006_223, w_006_224, w_006_225, w_006_226, w_006_227, w_006_228, w_006_229, w_006_230, w_006_231, w_006_232, w_006_233, w_006_234, w_006_235, w_006_236, w_006_237, w_006_238, w_006_239, w_006_240, w_006_241, w_006_242, w_006_243, w_006_244, w_006_245, w_006_246, w_006_247, w_006_248, w_006_249, w_006_250, w_006_251, w_006_252, w_006_253, w_006_254, w_006_255, w_006_256, w_006_257, w_006_258, w_006_259, w_006_260, w_006_261, w_006_262, w_006_263, w_006_264, w_006_265, w_006_266, w_006_267, w_006_268, w_006_269, w_006_270, w_006_271, w_006_272, w_006_273, w_006_274, w_006_275, w_006_276, w_006_277, w_006_278, w_006_279, w_006_280, w_006_281, w_006_282, w_006_283, w_006_284, w_006_285, w_006_286, w_006_287, w_006_288, w_006_289, w_006_290, w_006_291, w_006_292, w_006_293, w_006_294, w_006_295, w_006_296, w_006_297, w_006_298, w_006_299, w_006_300, w_006_301, w_006_302, w_006_303, w_006_304, w_006_305, w_006_306, w_006_307, w_006_308, w_006_309, w_006_310, w_006_311, w_006_312, w_006_313, w_006_314, w_006_315, w_006_316, w_006_317, w_006_318, w_006_319, w_006_320, w_006_321, w_006_322, w_006_323, w_006_324, w_006_325, w_006_326, w_006_327, w_006_328, w_006_329, w_006_330, w_006_331, w_006_332, w_006_333, w_006_334, w_006_335, w_006_336, w_006_337, w_006_338, w_006_339, w_006_340, w_006_341, w_006_342, w_006_343;
  wire w_007_000, w_007_001, w_007_002, w_007_003, w_007_005, w_007_009, w_007_013, w_007_014, w_007_015, w_007_017, w_007_018, w_007_019, w_007_020, w_007_021, w_007_022, w_007_023, w_007_024, w_007_025, w_007_026, w_007_027, w_007_028, w_007_030, w_007_031, w_007_032, w_007_033, w_007_034, w_007_035, w_007_036, w_007_037, w_007_038, w_007_039, w_007_042, w_007_043, w_007_044, w_007_045, w_007_046, w_007_048, w_007_049, w_007_051, w_007_053, w_007_054, w_007_055, w_007_057, w_007_058, w_007_059, w_007_060, w_007_061, w_007_062, w_007_063, w_007_064, w_007_066, w_007_068, w_007_069, w_007_071, w_007_072, w_007_074, w_007_077, w_007_079, w_007_080, w_007_081, w_007_082, w_007_084, w_007_085, w_007_088, w_007_090, w_007_091, w_007_092, w_007_095, w_007_097, w_007_098, w_007_101, w_007_102, w_007_103, w_007_104, w_007_105, w_007_106, w_007_107, w_007_108, w_007_109, w_007_110, w_007_111, w_007_113, w_007_114, w_007_115, w_007_118, w_007_119, w_007_120, w_007_121, w_007_124, w_007_125, w_007_126, w_007_127, w_007_128, w_007_130, w_007_131, w_007_132, w_007_135, w_007_136, w_007_137, w_007_138, w_007_141, w_007_144, w_007_146, w_007_147, w_007_148, w_007_149, w_007_151, w_007_152, w_007_154, w_007_155, w_007_157, w_007_158, w_007_159, w_007_162, w_007_164, w_007_166, w_007_168, w_007_170, w_007_171, w_007_174, w_007_175, w_007_176, w_007_181, w_007_182, w_007_183, w_007_186, w_007_187, w_007_188, w_007_189, w_007_190, w_007_193, w_007_194, w_007_199, w_007_200, w_007_202, w_007_203, w_007_205, w_007_206, w_007_207, w_007_208, w_007_209, w_007_210, w_007_211, w_007_212, w_007_213, w_007_214, w_007_215, w_007_216, w_007_218, w_007_221, w_007_222, w_007_223, w_007_224, w_007_225, w_007_228, w_007_229, w_007_230, w_007_232, w_007_233, w_007_235, w_007_236, w_007_237, w_007_238, w_007_241, w_007_243, w_007_244, w_007_245, w_007_247, w_007_251, w_007_252, w_007_253, w_007_255, w_007_257, w_007_258, w_007_261, w_007_264, w_007_266, w_007_267, w_007_268, w_007_269, w_007_270, w_007_271, w_007_272, w_007_275, w_007_277, w_007_278, w_007_279, w_007_280, w_007_283, w_007_285, w_007_288, w_007_289, w_007_290, w_007_292, w_007_293, w_007_294, w_007_295, w_007_298, w_007_299, w_007_304, w_007_305, w_007_306, w_007_307, w_007_309, w_007_311, w_007_313, w_007_314, w_007_315, w_007_316, w_007_317, w_007_318, w_007_320, w_007_322, w_007_325, w_007_327, w_007_329, w_007_330, w_007_337, w_007_338, w_007_340, w_007_342, w_007_346, w_007_348, w_007_349, w_007_351, w_007_353, w_007_354, w_007_357, w_007_358, w_007_359, w_007_360, w_007_364, w_007_366, w_007_367, w_007_368, w_007_370, w_007_373, w_007_377, w_007_378, w_007_379, w_007_380, w_007_381, w_007_382, w_007_384, w_007_388, w_007_391, w_007_393, w_007_398, w_007_399, w_007_401, w_007_402, w_007_405, w_007_406, w_007_411, w_007_415, w_007_417, w_007_418, w_007_421, w_007_423, w_007_434, w_007_436, w_007_438, w_007_439, w_007_441, w_007_442, w_007_443, w_007_444, w_007_446, w_007_447, w_007_449, w_007_451, w_007_453, w_007_458, w_007_463, w_007_466, w_007_475, w_007_477, w_007_478, w_007_479, w_007_482, w_007_483, w_007_484, w_007_485, w_007_490, w_007_491, w_007_498, w_007_503, w_007_509, w_007_515, w_007_517, w_007_518, w_007_520, w_007_523, w_007_524, w_007_525, w_007_526, w_007_531, w_007_532, w_007_534, w_007_539, w_007_540, w_007_543, w_007_544, w_007_546, w_007_547, w_007_549, w_007_550, w_007_555, w_007_559, w_007_561, w_007_563, w_007_564, w_007_567, w_007_568, w_007_569, w_007_573, w_007_576, w_007_577, w_007_579, w_007_580, w_007_583, w_007_586, w_007_589, w_007_590, w_007_592, w_007_597, w_007_598, w_007_599, w_007_601, w_007_603, w_007_604, w_007_605, w_007_609, w_007_610, w_007_612, w_007_613, w_007_618, w_007_622, w_007_623, w_007_624, w_007_627, w_007_628, w_007_632, w_007_634, w_007_636, w_007_637, w_007_638, w_007_639, w_007_640, w_007_646, w_007_652, w_007_654, w_007_655, w_007_656, w_007_657, w_007_660, w_007_663, w_007_664, w_007_666, w_007_673, w_007_676, w_007_680, w_007_682, w_007_687, w_007_689, w_007_691, w_007_697, w_007_698, w_007_699, w_007_701, w_007_703, w_007_704, w_007_712, w_007_713, w_007_714, w_007_715, w_007_720, w_007_722, w_007_725, w_007_726, w_007_729, w_007_732, w_007_734, w_007_738, w_007_740, w_007_741, w_007_742, w_007_744, w_007_746, w_007_747, w_007_750, w_007_752, w_007_755, w_007_756, w_007_757, w_007_761, w_007_763, w_007_768, w_007_769, w_007_772, w_007_774, w_007_778, w_007_779, w_007_781, w_007_782, w_007_784, w_007_785, w_007_786, w_007_790, w_007_793, w_007_796, w_007_798, w_007_800, w_007_802, w_007_803, w_007_804, w_007_805, w_007_808, w_007_811, w_007_814, w_007_816, w_007_817, w_007_822, w_007_823, w_007_828, w_007_829, w_007_834, w_007_837, w_007_838, w_007_839, w_007_840, w_007_847, w_007_849, w_007_850, w_007_851, w_007_855, w_007_858, w_007_860, w_007_862, w_007_863, w_007_865, w_007_869, w_007_871, w_007_873, w_007_874, w_007_875, w_007_879, w_007_880, w_007_881, w_007_883, w_007_884, w_007_887, w_007_889, w_007_891, w_007_892, w_007_894, w_007_900, w_007_903, w_007_904, w_007_905, w_007_907, w_007_915, w_007_916, w_007_920, w_007_921, w_007_924, w_007_925, w_007_927, w_007_928, w_007_929, w_007_931, w_007_934, w_007_935, w_007_941, w_007_944, w_007_945, w_007_946, w_007_947, w_007_948, w_007_951, w_007_953, w_007_954, w_007_957, w_007_961, w_007_963, w_007_964, w_007_966, w_007_967, w_007_969, w_007_975, w_007_977, w_007_979, w_007_980, w_007_981, w_007_987, w_007_996, w_007_997, w_007_999, w_007_1002, w_007_1003, w_007_1010, w_007_1020, w_007_1022, w_007_1026, w_007_1033, w_007_1036, w_007_1042, w_007_1043, w_007_1044, w_007_1045, w_007_1046, w_007_1047, w_007_1048, w_007_1049, w_007_1054, w_007_1060, w_007_1061, w_007_1063, w_007_1065, w_007_1068, w_007_1069, w_007_1077, w_007_1078, w_007_1080, w_007_1083, w_007_1084, w_007_1085, w_007_1086, w_007_1087, w_007_1089, w_007_1090, w_007_1094, w_007_1095, w_007_1097, w_007_1101, w_007_1103, w_007_1104, w_007_1110, w_007_1117, w_007_1118, w_007_1119, w_007_1120, w_007_1123, w_007_1127, w_007_1129, w_007_1130, w_007_1132, w_007_1134, w_007_1137, w_007_1138, w_007_1140, w_007_1141, w_007_1142, w_007_1148, w_007_1151, w_007_1153, w_007_1157, w_007_1159, w_007_1160, w_007_1161, w_007_1168, w_007_1173, w_007_1175, w_007_1176, w_007_1178, w_007_1179, w_007_1182, w_007_1184, w_007_1187, w_007_1189, w_007_1190, w_007_1194, w_007_1197, w_007_1198, w_007_1204, w_007_1206, w_007_1208, w_007_1209, w_007_1211, w_007_1214, w_007_1215, w_007_1219, w_007_1223, w_007_1227, w_007_1229, w_007_1230, w_007_1231, w_007_1233, w_007_1234, w_007_1235, w_007_1243, w_007_1244, w_007_1245, w_007_1246, w_007_1247, w_007_1248, w_007_1250, w_007_1251, w_007_1256, w_007_1257, w_007_1258, w_007_1259, w_007_1261, w_007_1263, w_007_1264, w_007_1269, w_007_1276, w_007_1279, w_007_1281, w_007_1284, w_007_1292, w_007_1294, w_007_1295, w_007_1298, w_007_1299, w_007_1302, w_007_1303, w_007_1304, w_007_1307, w_007_1310, w_007_1313, w_007_1315, w_007_1316, w_007_1318, w_007_1321, w_007_1323, w_007_1326, w_007_1328, w_007_1331, w_007_1333, w_007_1334, w_007_1337, w_007_1338, w_007_1340, w_007_1341, w_007_1343, w_007_1345, w_007_1347, w_007_1349, w_007_1350, w_007_1351, w_007_1353, w_007_1355, w_007_1358, w_007_1360, w_007_1365, w_007_1366, w_007_1368, w_007_1374, w_007_1377, w_007_1378, w_007_1379, w_007_1384, w_007_1388, w_007_1390, w_007_1393, w_007_1397, w_007_1402, w_007_1405, w_007_1406, w_007_1407, w_007_1412, w_007_1415, w_007_1420, w_007_1423, w_007_1435, w_007_1436, w_007_1442, w_007_1443, w_007_1444, w_007_1446, w_007_1449, w_007_1450, w_007_1451, w_007_1454, w_007_1455, w_007_1456, w_007_1458, w_007_1459, w_007_1460, w_007_1462, w_007_1465, w_007_1467, w_007_1468, w_007_1469, w_007_1470, w_007_1472, w_007_1473, w_007_1474, w_007_1477, w_007_1478, w_007_1479, w_007_1480, w_007_1481, w_007_1482, w_007_1484, w_007_1486, w_007_1487, w_007_1488, w_007_1492, w_007_1493, w_007_1494, w_007_1495, w_007_1497, w_007_1500, w_007_1502, w_007_1504, w_007_1506, w_007_1507, w_007_1508, w_007_1510, w_007_1511, w_007_1512, w_007_1513, w_007_1515, w_007_1519, w_007_1520, w_007_1522, w_007_1524, w_007_1527, w_007_1530, w_007_1531, w_007_1533, w_007_1536, w_007_1538, w_007_1543, w_007_1551, w_007_1554, w_007_1555, w_007_1562, w_007_1565, w_007_1566, w_007_1567, w_007_1570, w_007_1574, w_007_1579, w_007_1583, w_007_1584, w_007_1588, w_007_1590, w_007_1592, w_007_1593, w_007_1594, w_007_1595, w_007_1596, w_007_1597, w_007_1598, w_007_1599, w_007_1600, w_007_1601, w_007_1603, w_007_1605, w_007_1606, w_007_1615, w_007_1616, w_007_1617, w_007_1618, w_007_1619, w_007_1620;
  wire w_008_002, w_008_003, w_008_005, w_008_006, w_008_008, w_008_009, w_008_010, w_008_011, w_008_013, w_008_014, w_008_015, w_008_016, w_008_017, w_008_018, w_008_019, w_008_020, w_008_021, w_008_022, w_008_023, w_008_024, w_008_025, w_008_026, w_008_027, w_008_028, w_008_031, w_008_032, w_008_034, w_008_035, w_008_036, w_008_038, w_008_039, w_008_040, w_008_041, w_008_043, w_008_044, w_008_046, w_008_047, w_008_049, w_008_051, w_008_052, w_008_053, w_008_056, w_008_058, w_008_059, w_008_060, w_008_061, w_008_062, w_008_064, w_008_065, w_008_066, w_008_067, w_008_069, w_008_070, w_008_071, w_008_073, w_008_074, w_008_076, w_008_077, w_008_078, w_008_079, w_008_081, w_008_082, w_008_084, w_008_085, w_008_087, w_008_088, w_008_089, w_008_090, w_008_092, w_008_093, w_008_094, w_008_095, w_008_096, w_008_098, w_008_100, w_008_102, w_008_103, w_008_104, w_008_106, w_008_108, w_008_109, w_008_110, w_008_111, w_008_112, w_008_114, w_008_115, w_008_117, w_008_119, w_008_122, w_008_123, w_008_124, w_008_125, w_008_126, w_008_127, w_008_128, w_008_129, w_008_130, w_008_132, w_008_133, w_008_134, w_008_136, w_008_139, w_008_143, w_008_144, w_008_147, w_008_148, w_008_151, w_008_152, w_008_154, w_008_156, w_008_157, w_008_158, w_008_160, w_008_162, w_008_163, w_008_164, w_008_165, w_008_166, w_008_167, w_008_168, w_008_170, w_008_172, w_008_174, w_008_175, w_008_176, w_008_177, w_008_180, w_008_181, w_008_182, w_008_184, w_008_185, w_008_186, w_008_187, w_008_188, w_008_190, w_008_192, w_008_193, w_008_195, w_008_196, w_008_197, w_008_198, w_008_199, w_008_200, w_008_201, w_008_202, w_008_203, w_008_205, w_008_206, w_008_207, w_008_208, w_008_209, w_008_210, w_008_211, w_008_212, w_008_213, w_008_216, w_008_217, w_008_218, w_008_219, w_008_222, w_008_224, w_008_225, w_008_228, w_008_230, w_008_231, w_008_233, w_008_234, w_008_235, w_008_236, w_008_237, w_008_238, w_008_240, w_008_241, w_008_242, w_008_243, w_008_244, w_008_245, w_008_246, w_008_247, w_008_248, w_008_250, w_008_251, w_008_252, w_008_253, w_008_254, w_008_256, w_008_257, w_008_258, w_008_259, w_008_260, w_008_261, w_008_262, w_008_263, w_008_264, w_008_266, w_008_268, w_008_269, w_008_270, w_008_271, w_008_273, w_008_275, w_008_276, w_008_277, w_008_278, w_008_279, w_008_280, w_008_281, w_008_282, w_008_285, w_008_286, w_008_288, w_008_289, w_008_290, w_008_293, w_008_294, w_008_296, w_008_297, w_008_298, w_008_300, w_008_301, w_008_303, w_008_306, w_008_308, w_008_310, w_008_312, w_008_314, w_008_315, w_008_316, w_008_317, w_008_318, w_008_319, w_008_324, w_008_326, w_008_327, w_008_330, w_008_332, w_008_336, w_008_342, w_008_343, w_008_344, w_008_345, w_008_346, w_008_348, w_008_349, w_008_351, w_008_352, w_008_353, w_008_355, w_008_359, w_008_360, w_008_362, w_008_364, w_008_365, w_008_368, w_008_369, w_008_370, w_008_372, w_008_373, w_008_374, w_008_376, w_008_379, w_008_380, w_008_381, w_008_382, w_008_384, w_008_386, w_008_390, w_008_393, w_008_394, w_008_395, w_008_396, w_008_399, w_008_400, w_008_401, w_008_402, w_008_404, w_008_407, w_008_408, w_008_412, w_008_413, w_008_415, w_008_417, w_008_418, w_008_419, w_008_420, w_008_421, w_008_422, w_008_423, w_008_424, w_008_425, w_008_426, w_008_428, w_008_429, w_008_431, w_008_433, w_008_434, w_008_435, w_008_436, w_008_437, w_008_438, w_008_442, w_008_443, w_008_444, w_008_445, w_008_447, w_008_449, w_008_450, w_008_453, w_008_454, w_008_455, w_008_456, w_008_457, w_008_459, w_008_460, w_008_461, w_008_463, w_008_464, w_008_465, w_008_470, w_008_472, w_008_473, w_008_474, w_008_475, w_008_477, w_008_479, w_008_480, w_008_481, w_008_484, w_008_485, w_008_488, w_008_489, w_008_490, w_008_491, w_008_495, w_008_500, w_008_501, w_008_502, w_008_504, w_008_506, w_008_507, w_008_511, w_008_513, w_008_515, w_008_518, w_008_519, w_008_521, w_008_524, w_008_525, w_008_526, w_008_527, w_008_530, w_008_531, w_008_533, w_008_534, w_008_537, w_008_538, w_008_540, w_008_541, w_008_543, w_008_544, w_008_546, w_008_547, w_008_549, w_008_550, w_008_551, w_008_552, w_008_553, w_008_554, w_008_555, w_008_556, w_008_560, w_008_562, w_008_563, w_008_564, w_008_566, w_008_567, w_008_569, w_008_570, w_008_572, w_008_573, w_008_574, w_008_577, w_008_578, w_008_579, w_008_580, w_008_584, w_008_589, w_008_591, w_008_593, w_008_594, w_008_595, w_008_597, w_008_599, w_008_602, w_008_603, w_008_605, w_008_608, w_008_609, w_008_610, w_008_611, w_008_612, w_008_615, w_008_616, w_008_618, w_008_619, w_008_620, w_008_621, w_008_622, w_008_624, w_008_626, w_008_627, w_008_628, w_008_632, w_008_633, w_008_635, w_008_638, w_008_639, w_008_644, w_008_645, w_008_646, w_008_651, w_008_652, w_008_653, w_008_656, w_008_657, w_008_659, w_008_660, w_008_661, w_008_662, w_008_663, w_008_664, w_008_666, w_008_668, w_008_670, w_008_673, w_008_674, w_008_675, w_008_677, w_008_678, w_008_679, w_008_680, w_008_681, w_008_682, w_008_683, w_008_684, w_008_685, w_008_686, w_008_688, w_008_689, w_008_691, w_008_692, w_008_694, w_008_696, w_008_698, w_008_699, w_008_702, w_008_703, w_008_704, w_008_705, w_008_706, w_008_707, w_008_709, w_008_712, w_008_713, w_008_714, w_008_717, w_008_718, w_008_719, w_008_720, w_008_721, w_008_727, w_008_728, w_008_729, w_008_731, w_008_732, w_008_734, w_008_735, w_008_738, w_008_739, w_008_741, w_008_742, w_008_743, w_008_744, w_008_745, w_008_747, w_008_748, w_008_749, w_008_750, w_008_751, w_008_752, w_008_753, w_008_755, w_008_756, w_008_758, w_008_759, w_008_760, w_008_761, w_008_762, w_008_763, w_008_764, w_008_765, w_008_766, w_008_767, w_008_769, w_008_770, w_008_771, w_008_772, w_008_773, w_008_776, w_008_778, w_008_779, w_008_783, w_008_785, w_008_787, w_008_788, w_008_790, w_008_791, w_008_793, w_008_794, w_008_795, w_008_796, w_008_798, w_008_799, w_008_801, w_008_802, w_008_804, w_008_805, w_008_806, w_008_807, w_008_808, w_008_809, w_008_810, w_008_811, w_008_813, w_008_815, w_008_817, w_008_818, w_008_819, w_008_821, w_008_823, w_008_825, w_008_829, w_008_830, w_008_831, w_008_833, w_008_836, w_008_838, w_008_841, w_008_847, w_008_850, w_008_851, w_008_853, w_008_856, w_008_857, w_008_858, w_008_861, w_008_862;
  wire w_009_000, w_009_001, w_009_002, w_009_003, w_009_004, w_009_005, w_009_006, w_009_007, w_009_008, w_009_009, w_009_010, w_009_011, w_009_012, w_009_013, w_009_014, w_009_015, w_009_016, w_009_017, w_009_018, w_009_019, w_009_020, w_009_021, w_009_022, w_009_023, w_009_024, w_009_025, w_009_026, w_009_027, w_009_028, w_009_029, w_009_030, w_009_031, w_009_032, w_009_033, w_009_034, w_009_035, w_009_036, w_009_037, w_009_038, w_009_039, w_009_040, w_009_041, w_009_042, w_009_043, w_009_044, w_009_045, w_009_046, w_009_047, w_009_048, w_009_049, w_009_050, w_009_051, w_009_052, w_009_053, w_009_054, w_009_055, w_009_056, w_009_057, w_009_058, w_009_059, w_009_060, w_009_061, w_009_062, w_009_063, w_009_064, w_009_065, w_009_066, w_009_067, w_009_068, w_009_069, w_009_070, w_009_071, w_009_072, w_009_073, w_009_074, w_009_075, w_009_076, w_009_077, w_009_078, w_009_079, w_009_080, w_009_081, w_009_082, w_009_083, w_009_084, w_009_085, w_009_086, w_009_087, w_009_088, w_009_089, w_009_090, w_009_091, w_009_092, w_009_093, w_009_094, w_009_095, w_009_096, w_009_097, w_009_098, w_009_099, w_009_100, w_009_101, w_009_102, w_009_103, w_009_104, w_009_105, w_009_106, w_009_107, w_009_108, w_009_109, w_009_110, w_009_111, w_009_113, w_009_114, w_009_115, w_009_116, w_009_117, w_009_118, w_009_119, w_009_120, w_009_122, w_009_124, w_009_125, w_009_126, w_009_127, w_009_128, w_009_129, w_009_131;
  wire w_010_001, w_010_002, w_010_003, w_010_004, w_010_005, w_010_006, w_010_007, w_010_008, w_010_009, w_010_010, w_010_011, w_010_012, w_010_013, w_010_014, w_010_015, w_010_017, w_010_018, w_010_019, w_010_020, w_010_021, w_010_022, w_010_023, w_010_024, w_010_025, w_010_026, w_010_027, w_010_028, w_010_029, w_010_030, w_010_031, w_010_032, w_010_033, w_010_034, w_010_035, w_010_036, w_010_037, w_010_038, w_010_039, w_010_040, w_010_041, w_010_042, w_010_043, w_010_044, w_010_045, w_010_046, w_010_047, w_010_048, w_010_049, w_010_050, w_010_051, w_010_054, w_010_055, w_010_056, w_010_057, w_010_058, w_010_059, w_010_060, w_010_061, w_010_062, w_010_063, w_010_064, w_010_065, w_010_066, w_010_067, w_010_068, w_010_069, w_010_070, w_010_071, w_010_073, w_010_074, w_010_076, w_010_077, w_010_078, w_010_079, w_010_080, w_010_081, w_010_082, w_010_083, w_010_084, w_010_085, w_010_086, w_010_087, w_010_088, w_010_089, w_010_090, w_010_091, w_010_092, w_010_093, w_010_094, w_010_095, w_010_096, w_010_097, w_010_098, w_010_099, w_010_101, w_010_102, w_010_103, w_010_104, w_010_105, w_010_106, w_010_108, w_010_109, w_010_110, w_010_111, w_010_112, w_010_113, w_010_114, w_010_115, w_010_116, w_010_117, w_010_118, w_010_119, w_010_121, w_010_122, w_010_123, w_010_124, w_010_125, w_010_126, w_010_127, w_010_128, w_010_129, w_010_131, w_010_132, w_010_133, w_010_134, w_010_135, w_010_136, w_010_138, w_010_139, w_010_140, w_010_141, w_010_146, w_010_147, w_010_149, w_010_150, w_010_151, w_010_153, w_010_154, w_010_155, w_010_156, w_010_157, w_010_158, w_010_159, w_010_160, w_010_161, w_010_162, w_010_163, w_010_164, w_010_165, w_010_166, w_010_167, w_010_168, w_010_169, w_010_170, w_010_171, w_010_172, w_010_173, w_010_174, w_010_175, w_010_176, w_010_177, w_010_178, w_010_180, w_010_181, w_010_184, w_010_185, w_010_186, w_010_188, w_010_189, w_010_190, w_010_191, w_010_192, w_010_193, w_010_194, w_010_196, w_010_197, w_010_198, w_010_199, w_010_200, w_010_201, w_010_202, w_010_203, w_010_204, w_010_205, w_010_206, w_010_207, w_010_208, w_010_210, w_010_211, w_010_212, w_010_213, w_010_214, w_010_215, w_010_216, w_010_217, w_010_219, w_010_220, w_010_221, w_010_222, w_010_223, w_010_224, w_010_225, w_010_226, w_010_227, w_010_228, w_010_229, w_010_230, w_010_231, w_010_233, w_010_234, w_010_235, w_010_236, w_010_237, w_010_238, w_010_239, w_010_241, w_010_242, w_010_244, w_010_245, w_010_246, w_010_247, w_010_248, w_010_250, w_010_251, w_010_252, w_010_253, w_010_254, w_010_256, w_010_259, w_010_260, w_010_261, w_010_262, w_010_263, w_010_264, w_010_265, w_010_266, w_010_267, w_010_268, w_010_269, w_010_270, w_010_271, w_010_272, w_010_273, w_010_274, w_010_275, w_010_276, w_010_277, w_010_278, w_010_279, w_010_280, w_010_281, w_010_282, w_010_283, w_010_284, w_010_285, w_010_286, w_010_287, w_010_288, w_010_290, w_010_291, w_010_292, w_010_293, w_010_294, w_010_295, w_010_297, w_010_298, w_010_299, w_010_300, w_010_302, w_010_303, w_010_304, w_010_305, w_010_306, w_010_307, w_010_308, w_010_309, w_010_310, w_010_311, w_010_312, w_010_315, w_010_316, w_010_317, w_010_318, w_010_320, w_010_321, w_010_322, w_010_323, w_010_324, w_010_325, w_010_326, w_010_327, w_010_328, w_010_329, w_010_330, w_010_331, w_010_332, w_010_333, w_010_334, w_010_336, w_010_337, w_010_338, w_010_339, w_010_342, w_010_343, w_010_344, w_010_345, w_010_346, w_010_347, w_010_348, w_010_350, w_010_351, w_010_352, w_010_353, w_010_354, w_010_355, w_010_356, w_010_357, w_010_358, w_010_359, w_010_360, w_010_363, w_010_365, w_010_366, w_010_367, w_010_369, w_010_370, w_010_371, w_010_372, w_010_373, w_010_374, w_010_375, w_010_376, w_010_377, w_010_378, w_010_379, w_010_380, w_010_381, w_010_382, w_010_384, w_010_385, w_010_386, w_010_387, w_010_388, w_010_391, w_010_392, w_010_394, w_010_397, w_010_398, w_010_399, w_010_400, w_010_401, w_010_402, w_010_403, w_010_405, w_010_406, w_010_408, w_010_411, w_010_413, w_010_414, w_010_415, w_010_416, w_010_417, w_010_419, w_010_420;
  wire w_011_000, w_011_001, w_011_002, w_011_003, w_011_004, w_011_005, w_011_006, w_011_007, w_011_009, w_011_010, w_011_011, w_011_014, w_011_015, w_011_016, w_011_018, w_011_019, w_011_020, w_011_021, w_011_022, w_011_026, w_011_028, w_011_031, w_011_033, w_011_034, w_011_035, w_011_036, w_011_037, w_011_038, w_011_039, w_011_040, w_011_041, w_011_042, w_011_043, w_011_044, w_011_046, w_011_051, w_011_052, w_011_056, w_011_057, w_011_058, w_011_060, w_011_062, w_011_063, w_011_064, w_011_065, w_011_067, w_011_068, w_011_070, w_011_071, w_011_072, w_011_073, w_011_074, w_011_076, w_011_077, w_011_079, w_011_080, w_011_081, w_011_085, w_011_086, w_011_088, w_011_091, w_011_092, w_011_093, w_011_094, w_011_097, w_011_098, w_011_100, w_011_101, w_011_102, w_011_103, w_011_104, w_011_105, w_011_107, w_011_108, w_011_109, w_011_111, w_011_112, w_011_114, w_011_115, w_011_117, w_011_118, w_011_119, w_011_120, w_011_122, w_011_123, w_011_125, w_011_126, w_011_127, w_011_128, w_011_129, w_011_132, w_011_133, w_011_135, w_011_136, w_011_137, w_011_140, w_011_141, w_011_142, w_011_143, w_011_144, w_011_147, w_011_148, w_011_150, w_011_151, w_011_152, w_011_154, w_011_155, w_011_157, w_011_159, w_011_160, w_011_161, w_011_163, w_011_164, w_011_166, w_011_169, w_011_170, w_011_171, w_011_172, w_011_173, w_011_176, w_011_177, w_011_181, w_011_182, w_011_184, w_011_185, w_011_188, w_011_189, w_011_190, w_011_193, w_011_194, w_011_196, w_011_197, w_011_199, w_011_201, w_011_203, w_011_204, w_011_205, w_011_206, w_011_208, w_011_209, w_011_210, w_011_213, w_011_215, w_011_216, w_011_217, w_011_219, w_011_221, w_011_224, w_011_225, w_011_227, w_011_228, w_011_229, w_011_230, w_011_232, w_011_233, w_011_235, w_011_242, w_011_243, w_011_244, w_011_246, w_011_247, w_011_250, w_011_256, w_011_257, w_011_258, w_011_260, w_011_262, w_011_263, w_011_265, w_011_267, w_011_272, w_011_273, w_011_283, w_011_286, w_011_290, w_011_293, w_011_295, w_011_297, w_011_298, w_011_303, w_011_304, w_011_307, w_011_309, w_011_313, w_011_314, w_011_315, w_011_316, w_011_318, w_011_320, w_011_323, w_011_324, w_011_325, w_011_327, w_011_328, w_011_332, w_011_333, w_011_334, w_011_338, w_011_339, w_011_344, w_011_345, w_011_347, w_011_350, w_011_353, w_011_354, w_011_357, w_011_360, w_011_361, w_011_363, w_011_365, w_011_368, w_011_369, w_011_371, w_011_372, w_011_374, w_011_378, w_011_381, w_011_383, w_011_384, w_011_386, w_011_388, w_011_389, w_011_390, w_011_391, w_011_394, w_011_395, w_011_398, w_011_401, w_011_402, w_011_403, w_011_404, w_011_405, w_011_406, w_011_407, w_011_411, w_011_412, w_011_414, w_011_417, w_011_419, w_011_420, w_011_424, w_011_425, w_011_426, w_011_428, w_011_429, w_011_432, w_011_433, w_011_435, w_011_436, w_011_439, w_011_440, w_011_441, w_011_444, w_011_445, w_011_449, w_011_453, w_011_454, w_011_455, w_011_459, w_011_460, w_011_461, w_011_463, w_011_464, w_011_465, w_011_466, w_011_469, w_011_470, w_011_471, w_011_474, w_011_475, w_011_479, w_011_480, w_011_482, w_011_483, w_011_485, w_011_489, w_011_490, w_011_491, w_011_492, w_011_493, w_011_496, w_011_498, w_011_501, w_011_503, w_011_504, w_011_508, w_011_509, w_011_510, w_011_512, w_011_515, w_011_517, w_011_522, w_011_523, w_011_525, w_011_527, w_011_532, w_011_533, w_011_534, w_011_536, w_011_538, w_011_539, w_011_541, w_011_542, w_011_543, w_011_546, w_011_547, w_011_548, w_011_550, w_011_551, w_011_552, w_011_553, w_011_557, w_011_559, w_011_560, w_011_565, w_011_568, w_011_572, w_011_573, w_011_574, w_011_575, w_011_576, w_011_578, w_011_579, w_011_580, w_011_582, w_011_583, w_011_584, w_011_586, w_011_587, w_011_588, w_011_589, w_011_592, w_011_594, w_011_596, w_011_597, w_011_598, w_011_610, w_011_611, w_011_613, w_011_617, w_011_619, w_011_620, w_011_622, w_011_623, w_011_624, w_011_626, w_011_628, w_011_631, w_011_633, w_011_635, w_011_638, w_011_639, w_011_640, w_011_642, w_011_643, w_011_645, w_011_648, w_011_650, w_011_652, w_011_653, w_011_654, w_011_659, w_011_660, w_011_665, w_011_666, w_011_667, w_011_669, w_011_670, w_011_674, w_011_676, w_011_677, w_011_678, w_011_679, w_011_680, w_011_685, w_011_687, w_011_688, w_011_691, w_011_692, w_011_694, w_011_695, w_011_696, w_011_698, w_011_699, w_011_700, w_011_702, w_011_703, w_011_704, w_011_705, w_011_706, w_011_707, w_011_708, w_011_711, w_011_715, w_011_716, w_011_718, w_011_721, w_011_725, w_011_727, w_011_731, w_011_733, w_011_734, w_011_735, w_011_738, w_011_739, w_011_741, w_011_742, w_011_743, w_011_749, w_011_751, w_011_752, w_011_753, w_011_755, w_011_757, w_011_758, w_011_762, w_011_763, w_011_764, w_011_765, w_011_770, w_011_771, w_011_773, w_011_775, w_011_779, w_011_780, w_011_782, w_011_783, w_011_785, w_011_787, w_011_790, w_011_791, w_011_794, w_011_795, w_011_796, w_011_798, w_011_800, w_011_802, w_011_803, w_011_804, w_011_805, w_011_809, w_011_810, w_011_811, w_011_813, w_011_814, w_011_815, w_011_816, w_011_817, w_011_819, w_011_822, w_011_826, w_011_829, w_011_830, w_011_832, w_011_833, w_011_835, w_011_836, w_011_837, w_011_838, w_011_839, w_011_840, w_011_845, w_011_846, w_011_848, w_011_849, w_011_850, w_011_852, w_011_853, w_011_854, w_011_856, w_011_857, w_011_858, w_011_861, w_011_862, w_011_865, w_011_866, w_011_867, w_011_869, w_011_870, w_011_871, w_011_872, w_011_875, w_011_876, w_011_877, w_011_878, w_011_879, w_011_881, w_011_883;
  wire w_012_000, w_012_002, w_012_003, w_012_006, w_012_007, w_012_008, w_012_011, w_012_016, w_012_017, w_012_018, w_012_020, w_012_021, w_012_022, w_012_023, w_012_025, w_012_026, w_012_027, w_012_029, w_012_031, w_012_033, w_012_034, w_012_035, w_012_036, w_012_039, w_012_040, w_012_041, w_012_042, w_012_043, w_012_044, w_012_045, w_012_049, w_012_050, w_012_051, w_012_052, w_012_053, w_012_054, w_012_056, w_012_058, w_012_059, w_012_061, w_012_065, w_012_066, w_012_067, w_012_068, w_012_071, w_012_073, w_012_075, w_012_076, w_012_077, w_012_078, w_012_079, w_012_083, w_012_085, w_012_087, w_012_090, w_012_091, w_012_093, w_012_094, w_012_095, w_012_096, w_012_097, w_012_099, w_012_100, w_012_101, w_012_102, w_012_104, w_012_105, w_012_106, w_012_107, w_012_109, w_012_110, w_012_111, w_012_112, w_012_116, w_012_119, w_012_122, w_012_123, w_012_125, w_012_129, w_012_130, w_012_132, w_012_133, w_012_137, w_012_139, w_012_141, w_012_142, w_012_143, w_012_144, w_012_145, w_012_146, w_012_147, w_012_153, w_012_154, w_012_155, w_012_156, w_012_157, w_012_159, w_012_161, w_012_162, w_012_163, w_012_164, w_012_165, w_012_166, w_012_168, w_012_169, w_012_170, w_012_171, w_012_172, w_012_173, w_012_174, w_012_175, w_012_176, w_012_177, w_012_180, w_012_181, w_012_183, w_012_184, w_012_186, w_012_187, w_012_188, w_012_189, w_012_191, w_012_193, w_012_194, w_012_195, w_012_196, w_012_198, w_012_199, w_012_201, w_012_202, w_012_204, w_012_205, w_012_206, w_012_209, w_012_210, w_012_211, w_012_212, w_012_213, w_012_214, w_012_215, w_012_216, w_012_217, w_012_218, w_012_219, w_012_221, w_012_222, w_012_223, w_012_224, w_012_227, w_012_228, w_012_229, w_012_231, w_012_232, w_012_233, w_012_235, w_012_236, w_012_237, w_012_238, w_012_239, w_012_240, w_012_241, w_012_242, w_012_243, w_012_246, w_012_249, w_012_250, w_012_252, w_012_254, w_012_255, w_012_257, w_012_258, w_012_259, w_012_260, w_012_261, w_012_262, w_012_264, w_012_265, w_012_266, w_012_268, w_012_269, w_012_270, w_012_271, w_012_272, w_012_273, w_012_274, w_012_276, w_012_277, w_012_278, w_012_279, w_012_281, w_012_284, w_012_287, w_012_288, w_012_289, w_012_290, w_012_292, w_012_293, w_012_294, w_012_295, w_012_297, w_012_298, w_012_302, w_012_304, w_012_305, w_012_307, w_012_310, w_012_314, w_012_316, w_012_317, w_012_319, w_012_320, w_012_322, w_012_323, w_012_324, w_012_326, w_012_327, w_012_328, w_012_329, w_012_330, w_012_332, w_012_334, w_012_336, w_012_337, w_012_338, w_012_339, w_012_340, w_012_341, w_012_342, w_012_343, w_012_345, w_012_346, w_012_348, w_012_349, w_012_350, w_012_351, w_012_353, w_012_355, w_012_356, w_012_357, w_012_362, w_012_364, w_012_366, w_012_368, w_012_369, w_012_370, w_012_371, w_012_372, w_012_373, w_012_374, w_012_375, w_012_376, w_012_377, w_012_378, w_012_384, w_012_387, w_012_388, w_012_390, w_012_392, w_012_393, w_012_394, w_012_395, w_012_399, w_012_400, w_012_401, w_012_402, w_012_403, w_012_404, w_012_405, w_012_406, w_012_407, w_012_409, w_012_410, w_012_411, w_012_412, w_012_413, w_012_416, w_012_421, w_012_422, w_012_425, w_012_426, w_012_428, w_012_429, w_012_430, w_012_431, w_012_435, w_012_436, w_012_438, w_012_441, w_012_442, w_012_445, w_012_446, w_012_447, w_012_449, w_012_450, w_012_451, w_012_452, w_012_453, w_012_454, w_012_455, w_012_459, w_012_460, w_012_461, w_012_464, w_012_465, w_012_466, w_012_467, w_012_468, w_012_469, w_012_470, w_012_471, w_012_472, w_012_474, w_012_475, w_012_476, w_012_477, w_012_478, w_012_482, w_012_484, w_012_486, w_012_487, w_012_488, w_012_490, w_012_493, w_012_494, w_012_497, w_012_500, w_012_502, w_012_503, w_012_504, w_012_505, w_012_506, w_012_507, w_012_508, w_012_509, w_012_510, w_012_511, w_012_512, w_012_513, w_012_514, w_012_515, w_012_517, w_012_519, w_012_520, w_012_521, w_012_522, w_012_523, w_012_524, w_012_525, w_012_526, w_012_527, w_012_529, w_012_530, w_012_531, w_012_535, w_012_536, w_012_537, w_012_538, w_012_541, w_012_545, w_012_546, w_012_547, w_012_550, w_012_551, w_012_552, w_012_554, w_012_555, w_012_556, w_012_557, w_012_558, w_012_559, w_012_560, w_012_561, w_012_563, w_012_564, w_012_567, w_012_569, w_012_570, w_012_571, w_012_572, w_012_573, w_012_574, w_012_578, w_012_579, w_012_580, w_012_581, w_012_582, w_012_585, w_012_586, w_012_587, w_012_588, w_012_589, w_012_590, w_012_591, w_012_592, w_012_594, w_012_596, w_012_597, w_012_598, w_012_599, w_012_603, w_012_607, w_012_608, w_012_609, w_012_612, w_012_613, w_012_614, w_012_616, w_012_617, w_012_618, w_012_619, w_012_620, w_012_621, w_012_625, w_012_626, w_012_627, w_012_628, w_012_629, w_012_631, w_012_632, w_012_633, w_012_635, w_012_636, w_012_637, w_012_639, w_012_640, w_012_641, w_012_642, w_012_643, w_012_646, w_012_648, w_012_649, w_012_650, w_012_652, w_012_653, w_012_654, w_012_655, w_012_656, w_012_657, w_012_659, w_012_660, w_012_661, w_012_662, w_012_663, w_012_666, w_012_667;
  wire w_013_000, w_013_001, w_013_002, w_013_003, w_013_004, w_013_006, w_013_008, w_013_009, w_013_010, w_013_011, w_013_012, w_013_013, w_013_014, w_013_015, w_013_016, w_013_017, w_013_018, w_013_019, w_013_021, w_013_022, w_013_023, w_013_024, w_013_025, w_013_026, w_013_027, w_013_028, w_013_029, w_013_030, w_013_031, w_013_032, w_013_033, w_013_035, w_013_036, w_013_038, w_013_040, w_013_041, w_013_043, w_013_044, w_013_045, w_013_046, w_013_047, w_013_048, w_013_049, w_013_050, w_013_051, w_013_052, w_013_053, w_013_054, w_013_055, w_013_057, w_013_058, w_013_059, w_013_060, w_013_061, w_013_062, w_013_063, w_013_064, w_013_066, w_013_067, w_013_068, w_013_069, w_013_070, w_013_072, w_013_073, w_013_074, w_013_075, w_013_076, w_013_077, w_013_078, w_013_080, w_013_081, w_013_083, w_013_084, w_013_085, w_013_086, w_013_087, w_013_088, w_013_089, w_013_090, w_013_091, w_013_092, w_013_093, w_013_094, w_013_095, w_013_096, w_013_097, w_013_098, w_013_099, w_013_100, w_013_101, w_013_102, w_013_103, w_013_104, w_013_105, w_013_106, w_013_107, w_013_108, w_013_109, w_013_110, w_013_111, w_013_112, w_013_113, w_013_114, w_013_115, w_013_116, w_013_117, w_013_118, w_013_119, w_013_120, w_013_121, w_013_122, w_013_123, w_013_124, w_013_125, w_013_126, w_013_127, w_013_131, w_013_132, w_013_133, w_013_134, w_013_135, w_013_136, w_013_137, w_013_139, w_013_140, w_013_141, w_013_142, w_013_143, w_013_144, w_013_145, w_013_147, w_013_148, w_013_149, w_013_150, w_013_151, w_013_153, w_013_154, w_013_155, w_013_156, w_013_159, w_013_160, w_013_161, w_013_162, w_013_163, w_013_164, w_013_165, w_013_167, w_013_168, w_013_169, w_013_170, w_013_171, w_013_172, w_013_173, w_013_174, w_013_175, w_013_176, w_013_177, w_013_178, w_013_179, w_013_180, w_013_181, w_013_182, w_013_183, w_013_184, w_013_185, w_013_186, w_013_187, w_013_188, w_013_189, w_013_190, w_013_191, w_013_192, w_013_194, w_013_197, w_013_198, w_013_199, w_013_201, w_013_203, w_013_205, w_013_206, w_013_207, w_013_209, w_013_210, w_013_211, w_013_212, w_013_214, w_013_215, w_013_216, w_013_217, w_013_219, w_013_221, w_013_222, w_013_223, w_013_225, w_013_226, w_013_227, w_013_228, w_013_229, w_013_230, w_013_231, w_013_233, w_013_234, w_013_235, w_013_236, w_013_237, w_013_239, w_013_240, w_013_242, w_013_243, w_013_244, w_013_245, w_013_247, w_013_248, w_013_249, w_013_250, w_013_251, w_013_252, w_013_253, w_013_254, w_013_255, w_013_257, w_013_258, w_013_259, w_013_260, w_013_261, w_013_263, w_013_264, w_013_265, w_013_266, w_013_267, w_013_268, w_013_270, w_013_271, w_013_272, w_013_273, w_013_274, w_013_275, w_013_278, w_013_279, w_013_280, w_013_281, w_013_282, w_013_283, w_013_284, w_013_285, w_013_286, w_013_287, w_013_288, w_013_289, w_013_290, w_013_291, w_013_292, w_013_293, w_013_294, w_013_295, w_013_296, w_013_297, w_013_298, w_013_299, w_013_300, w_013_301, w_013_302, w_013_303, w_013_304, w_013_305, w_013_307, w_013_309, w_013_311, w_013_312, w_013_313, w_013_314, w_013_315, w_013_316, w_013_318, w_013_319, w_013_320, w_013_321, w_013_323, w_013_324, w_013_325, w_013_326, w_013_327, w_013_328, w_013_330, w_013_331, w_013_332, w_013_335, w_013_336, w_013_337, w_013_338;
  wire w_014_001, w_014_002, w_014_003, w_014_005, w_014_008, w_014_013, w_014_014, w_014_015, w_014_017, w_014_018, w_014_019, w_014_020, w_014_022, w_014_023, w_014_024, w_014_025, w_014_027, w_014_029, w_014_032, w_014_038, w_014_040, w_014_041, w_014_043, w_014_049, w_014_051, w_014_053, w_014_055, w_014_056, w_014_058, w_014_059, w_014_060, w_014_061, w_014_065, w_014_070, w_014_072, w_014_074, w_014_076, w_014_077, w_014_078, w_014_079, w_014_080, w_014_082, w_014_084, w_014_085, w_014_086, w_014_087, w_014_089, w_014_090, w_014_091, w_014_092, w_014_093, w_014_094, w_014_097, w_014_099, w_014_101, w_014_102, w_014_104, w_014_106, w_014_107, w_014_108, w_014_109, w_014_110, w_014_112, w_014_115, w_014_116, w_014_117, w_014_118, w_014_119, w_014_121, w_014_123, w_014_124, w_014_125, w_014_129, w_014_130, w_014_131, w_014_132, w_014_133, w_014_136, w_014_138, w_014_140, w_014_142, w_014_143, w_014_144, w_014_145, w_014_147, w_014_149, w_014_150, w_014_151, w_014_154, w_014_156, w_014_157, w_014_158, w_014_159, w_014_160, w_014_161, w_014_163, w_014_164, w_014_165, w_014_167, w_014_168, w_014_169, w_014_171, w_014_172, w_014_177, w_014_178, w_014_179, w_014_181, w_014_184, w_014_189, w_014_191, w_014_193, w_014_194, w_014_195, w_014_196, w_014_197, w_014_199, w_014_203, w_014_204, w_014_205, w_014_208, w_014_209, w_014_210, w_014_211, w_014_212, w_014_213, w_014_214, w_014_218, w_014_219, w_014_221, w_014_223, w_014_225, w_014_226, w_014_229, w_014_232, w_014_234, w_014_235, w_014_237, w_014_239, w_014_242, w_014_243, w_014_246, w_014_247, w_014_248, w_014_249, w_014_251, w_014_252, w_014_255, w_014_256, w_014_257, w_014_258, w_014_261, w_014_262, w_014_263, w_014_264, w_014_266, w_014_268, w_014_270, w_014_271, w_014_272, w_014_273, w_014_274, w_014_276, w_014_277, w_014_278, w_014_279, w_014_280, w_014_286, w_014_288, w_014_290, w_014_291, w_014_293, w_014_295, w_014_296, w_014_299, w_014_300, w_014_304, w_014_308, w_014_309, w_014_310, w_014_311, w_014_312, w_014_313, w_014_314, w_014_315, w_014_316, w_014_318, w_014_319, w_014_320, w_014_321, w_014_322, w_014_323, w_014_324, w_014_326, w_014_327, w_014_329, w_014_330, w_014_333, w_014_334, w_014_335, w_014_337, w_014_340, w_014_341, w_014_342, w_014_344, w_014_345, w_014_349, w_014_352, w_014_353, w_014_359, w_014_360, w_014_361, w_014_362, w_014_365, w_014_366, w_014_370, w_014_372, w_014_375, w_014_376, w_014_380, w_014_383, w_014_384, w_014_385, w_014_387, w_014_390, w_014_392, w_014_393, w_014_397, w_014_398, w_014_402, w_014_403, w_014_405, w_014_406, w_014_411, w_014_412, w_014_416, w_014_417, w_014_420, w_014_422, w_014_426, w_014_427, w_014_430, w_014_432, w_014_433, w_014_434, w_014_436, w_014_437, w_014_438, w_014_439, w_014_442, w_014_443, w_014_445, w_014_447, w_014_451, w_014_453, w_014_454, w_014_457, w_014_459, w_014_461, w_014_465, w_014_467, w_014_469, w_014_470, w_014_473, w_014_475, w_014_477, w_014_478, w_014_481, w_014_483, w_014_486, w_014_487, w_014_489, w_014_491, w_014_492, w_014_495, w_014_500, w_014_502, w_014_504, w_014_505, w_014_506, w_014_508, w_014_509, w_014_512, w_014_516, w_014_517, w_014_518, w_014_519, w_014_520, w_014_523, w_014_524, w_014_525, w_014_526, w_014_528, w_014_529, w_014_532, w_014_533, w_014_534, w_014_537, w_014_540, w_014_543, w_014_544, w_014_545, w_014_547, w_014_551, w_014_556, w_014_560, w_014_561, w_014_565, w_014_567, w_014_569, w_014_573, w_014_574, w_014_576, w_014_577, w_014_578, w_014_579, w_014_581, w_014_582, w_014_583, w_014_586, w_014_588, w_014_590, w_014_598, w_014_599, w_014_601, w_014_604, w_014_606, w_014_607, w_014_609, w_014_611, w_014_613, w_014_614, w_014_617, w_014_619, w_014_623, w_014_624, w_014_626, w_014_629, w_014_632, w_014_636, w_014_639, w_014_640, w_014_641, w_014_643, w_014_644, w_014_646, w_014_648, w_014_649, w_014_650, w_014_651, w_014_652, w_014_653, w_014_654, w_014_659, w_014_661, w_014_662, w_014_663, w_014_664, w_014_666, w_014_668, w_014_672, w_014_673, w_014_677, w_014_685, w_014_686, w_014_688, w_014_690, w_014_691, w_014_692, w_014_696, w_014_702, w_014_703, w_014_704, w_014_707, w_014_708, w_014_709, w_014_711, w_014_713, w_014_716, w_014_717, w_014_719, w_014_721, w_014_722, w_014_723, w_014_726, w_014_728, w_014_729, w_014_732, w_014_734, w_014_736, w_014_738, w_014_740, w_014_745, w_014_746, w_014_752, w_014_755, w_014_757, w_014_767, w_014_768, w_014_772, w_014_777, w_014_780, w_014_784, w_014_787, w_014_793, w_014_795, w_014_796, w_014_798, w_014_801, w_014_805, w_014_806, w_014_807, w_014_808, w_014_809, w_014_810, w_014_814, w_014_815, w_014_819, w_014_821, w_014_822, w_014_823, w_014_824, w_014_825, w_014_826, w_014_829, w_014_830, w_014_831;
  wire w_015_000, w_015_001, w_015_002, w_015_003, w_015_004, w_015_005, w_015_006, w_015_007, w_015_008, w_015_010, w_015_011, w_015_012, w_015_013, w_015_014, w_015_015, w_015_016, w_015_017, w_015_019, w_015_020, w_015_021, w_015_022, w_015_023, w_015_024, w_015_025, w_015_026, w_015_027, w_015_030, w_015_031, w_015_032, w_015_033, w_015_034, w_015_035, w_015_036, w_015_038, w_015_039, w_015_040, w_015_041, w_015_042, w_015_043, w_015_044, w_015_045, w_015_046, w_015_047, w_015_048, w_015_049, w_015_050, w_015_052, w_015_053, w_015_055, w_015_056, w_015_057, w_015_058, w_015_059, w_015_060, w_015_061, w_015_062, w_015_064, w_015_065, w_015_066, w_015_067, w_015_068, w_015_069, w_015_070, w_015_071, w_015_073, w_015_074, w_015_075, w_015_076, w_015_077, w_015_078, w_015_079, w_015_080, w_015_081, w_015_082, w_015_083, w_015_084, w_015_086, w_015_087, w_015_088, w_015_089, w_015_090, w_015_091, w_015_093, w_015_094, w_015_097, w_015_099, w_015_100, w_015_101, w_015_103, w_015_104, w_015_105, w_015_106, w_015_108, w_015_110, w_015_112, w_015_113, w_015_115, w_015_116, w_015_117, w_015_118, w_015_119, w_015_120, w_015_122, w_015_124, w_015_125, w_015_126, w_015_127, w_015_128, w_015_129, w_015_130, w_015_131, w_015_133, w_015_134, w_015_135, w_015_136, w_015_137, w_015_138, w_015_140, w_015_141, w_015_142, w_015_143, w_015_144, w_015_146, w_015_147, w_015_149, w_015_150, w_015_151, w_015_152, w_015_153, w_015_154, w_015_155, w_015_157, w_015_158, w_015_159, w_015_160, w_015_161, w_015_162, w_015_163, w_015_164, w_015_165, w_015_166, w_015_168, w_015_169, w_015_170, w_015_171, w_015_172, w_015_173, w_015_174, w_015_176, w_015_177, w_015_178, w_015_181, w_015_183, w_015_184, w_015_185, w_015_186, w_015_187, w_015_188, w_015_189, w_015_190, w_015_191, w_015_192, w_015_193, w_015_194, w_015_195, w_015_196, w_015_198, w_015_199, w_015_200, w_015_201, w_015_203, w_015_204, w_015_205, w_015_206, w_015_207, w_015_208, w_015_209, w_015_210, w_015_211, w_015_212, w_015_213, w_015_214, w_015_216, w_015_217, w_015_218, w_015_219, w_015_220, w_015_221, w_015_222, w_015_223, w_015_224, w_015_225, w_015_226, w_015_227, w_015_228, w_015_229, w_015_230, w_015_232, w_015_234, w_015_235, w_015_236, w_015_237, w_015_238, w_015_240, w_015_241, w_015_242, w_015_243, w_015_244, w_015_245, w_015_246, w_015_247, w_015_248, w_015_249, w_015_250, w_015_251, w_015_252, w_015_253, w_015_254, w_015_255, w_015_256, w_015_257, w_015_258, w_015_259, w_015_260, w_015_261, w_015_262, w_015_264, w_015_265, w_015_266, w_015_267, w_015_268, w_015_270, w_015_271, w_015_273, w_015_274, w_015_275, w_015_276, w_015_277, w_015_278, w_015_279, w_015_280, w_015_281, w_015_282, w_015_283, w_015_285, w_015_286, w_015_287, w_015_288, w_015_289, w_015_290, w_015_291, w_015_293;
  wire w_016_000, w_016_001, w_016_002, w_016_003, w_016_004, w_016_005, w_016_006, w_016_007, w_016_008, w_016_009, w_016_010, w_016_011, w_016_012, w_016_013, w_016_014, w_016_015, w_016_016, w_016_017, w_016_018, w_016_019, w_016_020, w_016_021, w_016_022, w_016_023, w_016_024, w_016_025, w_016_026, w_016_027, w_016_028, w_016_029, w_016_030, w_016_031, w_016_032, w_016_033, w_016_034, w_016_035, w_016_036, w_016_037, w_016_038;
  wire w_017_002, w_017_003, w_017_005, w_017_006, w_017_007, w_017_010, w_017_012, w_017_013, w_017_014, w_017_016, w_017_017, w_017_018, w_017_019, w_017_020, w_017_022, w_017_023, w_017_029, w_017_032, w_017_033, w_017_034, w_017_036, w_017_038, w_017_040, w_017_044, w_017_045, w_017_046, w_017_047, w_017_052, w_017_057, w_017_059, w_017_075, w_017_077, w_017_084, w_017_085, w_017_087, w_017_088, w_017_089, w_017_100, w_017_102, w_017_106, w_017_117, w_017_124, w_017_133, w_017_141, w_017_142, w_017_143, w_017_150, w_017_155, w_017_158, w_017_159, w_017_162, w_017_171, w_017_174, w_017_179, w_017_183, w_017_194, w_017_197, w_017_198, w_017_203, w_017_205, w_017_211, w_017_214, w_017_218, w_017_225, w_017_229, w_017_234, w_017_236, w_017_240, w_017_244, w_017_251, w_017_253, w_017_254, w_017_264, w_017_269, w_017_282, w_017_288, w_017_299, w_017_300, w_017_303, w_017_305, w_017_307, w_017_315, w_017_317, w_017_322, w_017_324, w_017_325, w_017_326, w_017_333, w_017_334, w_017_335, w_017_346, w_017_352, w_017_360, w_017_366, w_017_368, w_017_373, w_017_381, w_017_384, w_017_385, w_017_386, w_017_390, w_017_393, w_017_396, w_017_397, w_017_398, w_017_404, w_017_408, w_017_411, w_017_413, w_017_417, w_017_427, w_017_428, w_017_429, w_017_432, w_017_434, w_017_436, w_017_442, w_017_446, w_017_450, w_017_457, w_017_459, w_017_468, w_017_471, w_017_472, w_017_476, w_017_478, w_017_479, w_017_482, w_017_485, w_017_491, w_017_502, w_017_507, w_017_508, w_017_513, w_017_524, w_017_525, w_017_528, w_017_534, w_017_539, w_017_540, w_017_549, w_017_551, w_017_556, w_017_558, w_017_562, w_017_589, w_017_595, w_017_602, w_017_605, w_017_615, w_017_616, w_017_619, w_017_622, w_017_623, w_017_624, w_017_631, w_017_633, w_017_644, w_017_647, w_017_649, w_017_664, w_017_665, w_017_666, w_017_673, w_017_675, w_017_677, w_017_678, w_017_681, w_017_684, w_017_685, w_017_687, w_017_691, w_017_694, w_017_697, w_017_702, w_017_703, w_017_704, w_017_707, w_017_713, w_017_722, w_017_723, w_017_730, w_017_732, w_017_734, w_017_736, w_017_740, w_017_742, w_017_743, w_017_744, w_017_748, w_017_753, w_017_773, w_017_774, w_017_777, w_017_779, w_017_781, w_017_798, w_017_804, w_017_805, w_017_809, w_017_812, w_017_813, w_017_821, w_017_838, w_017_841, w_017_845, w_017_846, w_017_847, w_017_851, w_017_858, w_017_863, w_017_864, w_017_867, w_017_871, w_017_873, w_017_875, w_017_885, w_017_891, w_017_895, w_017_896, w_017_899, w_017_902, w_017_903, w_017_905, w_017_914, w_017_917, w_017_921, w_017_929, w_017_932, w_017_933, w_017_935, w_017_944, w_017_947, w_017_950, w_017_953, w_017_956, w_017_960, w_017_967, w_017_975, w_017_977, w_017_982, w_017_984, w_017_985, w_017_990, w_017_998, w_017_1000, w_017_1001, w_017_1005, w_017_1006, w_017_1008, w_017_1014, w_017_1020, w_017_1023, w_017_1026, w_017_1031, w_017_1036, w_017_1041, w_017_1043, w_017_1047, w_017_1049, w_017_1051, w_017_1058, w_017_1059, w_017_1060, w_017_1065, w_017_1067, w_017_1070, w_017_1071, w_017_1074, w_017_1077, w_017_1079, w_017_1092, w_017_1098, w_017_1101, w_017_1103, w_017_1104, w_017_1109, w_017_1111, w_017_1113, w_017_1116, w_017_1123, w_017_1126, w_017_1128, w_017_1129, w_017_1131, w_017_1133, w_017_1135, w_017_1139, w_017_1140, w_017_1143, w_017_1145, w_017_1153, w_017_1163, w_017_1165, w_017_1179, w_017_1182, w_017_1195, w_017_1201, w_017_1206, w_017_1207, w_017_1214, w_017_1216, w_017_1218, w_017_1220, w_017_1223, w_017_1224, w_017_1226, w_017_1227, w_017_1231, w_017_1232, w_017_1237, w_017_1238, w_017_1240, w_017_1241, w_017_1242, w_017_1244, w_017_1246, w_017_1250, w_017_1262, w_017_1269, w_017_1271, w_017_1280, w_017_1284, w_017_1288, w_017_1301, w_017_1308, w_017_1310, w_017_1312, w_017_1322, w_017_1325, w_017_1327, w_017_1333, w_017_1336, w_017_1340, w_017_1348, w_017_1351, w_017_1354, w_017_1357, w_017_1365, w_017_1366, w_017_1369, w_017_1370, w_017_1372, w_017_1373, w_017_1374, w_017_1379, w_017_1380, w_017_1381, w_017_1383, w_017_1388, w_017_1391, w_017_1392, w_017_1393, w_017_1396, w_017_1397, w_017_1400, w_017_1402, w_017_1407, w_017_1410, w_017_1416, w_017_1419, w_017_1421, w_017_1422, w_017_1423, w_017_1430, w_017_1439, w_017_1443, w_017_1445, w_017_1448, w_017_1449, w_017_1453, w_017_1457, w_017_1460, w_017_1464, w_017_1469, w_017_1480, w_017_1497, w_017_1504, w_017_1505, w_017_1517, w_017_1530, w_017_1531, w_017_1533, w_017_1534, w_017_1541, w_017_1550, w_017_1552, w_017_1556, w_017_1557, w_017_1563, w_017_1575, w_017_1576, w_017_1578, w_017_1583, w_017_1586, w_017_1588, w_017_1591, w_017_1595, w_017_1598, w_017_1606, w_017_1607, w_017_1612, w_017_1622, w_017_1626, w_017_1630, w_017_1633, w_017_1636, w_017_1639, w_017_1640, w_017_1645, w_017_1646, w_017_1654, w_017_1655, w_017_1656, w_017_1658, w_017_1665, w_017_1666, w_017_1670, w_017_1671, w_017_1672, w_017_1679, w_017_1686, w_017_1689, w_017_1694, w_017_1706, w_017_1707, w_017_1710, w_017_1715, w_017_1718, w_017_1727, w_017_1729, w_017_1732, w_017_1738, w_017_1743, w_017_1750, w_017_1753, w_017_1763, w_017_1768, w_017_1778, w_017_1792, w_017_1797, w_017_1802, w_017_1809, w_017_1814, w_017_1816, w_017_1818, w_017_1822, w_017_1823, w_017_1828, w_017_1831, w_017_1839, w_017_1852, w_017_1857, w_017_1860, w_017_1866, w_017_1870, w_017_1871, w_017_1873, w_017_1877, w_017_1878, w_017_1881, w_017_1882, w_017_1885, w_017_1888, w_017_1893, w_017_1895, w_017_1900, w_017_1903, w_017_1910, w_017_1911, w_017_1913, w_017_1923, w_017_1924, w_017_1935, w_017_1937, w_017_1945, w_017_1947;
  wire w_018_003, w_018_004, w_018_005, w_018_006, w_018_007, w_018_008, w_018_009, w_018_010, w_018_011, w_018_012, w_018_013, w_018_014, w_018_015, w_018_016, w_018_017, w_018_018, w_018_019, w_018_021, w_018_022, w_018_024, w_018_025, w_018_026, w_018_027, w_018_028, w_018_029, w_018_030, w_018_031, w_018_032, w_018_033, w_018_035, w_018_036, w_018_037, w_018_038, w_018_039, w_018_040, w_018_041, w_018_043, w_018_044, w_018_045, w_018_046, w_018_047, w_018_048, w_018_049, w_018_050, w_018_052, w_018_054, w_018_055, w_018_056, w_018_057, w_018_059, w_018_061, w_018_063, w_018_064, w_018_065, w_018_066, w_018_067, w_018_068, w_018_069, w_018_070, w_018_071, w_018_072, w_018_073, w_018_075, w_018_077, w_018_078, w_018_079, w_018_080, w_018_081, w_018_082, w_018_084, w_018_085, w_018_086, w_018_087, w_018_088, w_018_089, w_018_090, w_018_091, w_018_092, w_018_094, w_018_097, w_018_098, w_018_100, w_018_101, w_018_102, w_018_103, w_018_104, w_018_105, w_018_107, w_018_108, w_018_109, w_018_110, w_018_111, w_018_112, w_018_113, w_018_114, w_018_115, w_018_117, w_018_118, w_018_119, w_018_120, w_018_121, w_018_122, w_018_124, w_018_125, w_018_127, w_018_128, w_018_129, w_018_131, w_018_132, w_018_133, w_018_134, w_018_135, w_018_136, w_018_137, w_018_138, w_018_139, w_018_140, w_018_141, w_018_142, w_018_143, w_018_144, w_018_145, w_018_146, w_018_147, w_018_148, w_018_149, w_018_150, w_018_151, w_018_152, w_018_153, w_018_155, w_018_156, w_018_157, w_018_158, w_018_159, w_018_160, w_018_161, w_018_162, w_018_163, w_018_165, w_018_167, w_018_168, w_018_170, w_018_171, w_018_172, w_018_175, w_018_176, w_018_178, w_018_180, w_018_181, w_018_182, w_018_183, w_018_184, w_018_186, w_018_187, w_018_189, w_018_190, w_018_191, w_018_192, w_018_193, w_018_194, w_018_195, w_018_196, w_018_197, w_018_198, w_018_200, w_018_201, w_018_202, w_018_203, w_018_204, w_018_205, w_018_206, w_018_207, w_018_209, w_018_210, w_018_211, w_018_212, w_018_213, w_018_214, w_018_215, w_018_216, w_018_218, w_018_219, w_018_220, w_018_221, w_018_222, w_018_223, w_018_224, w_018_225, w_018_226, w_018_227, w_018_228, w_018_229, w_018_230, w_018_231, w_018_232, w_018_233, w_018_234, w_018_235, w_018_236, w_018_237, w_018_239, w_018_240, w_018_241, w_018_242, w_018_243, w_018_244, w_018_245, w_018_246, w_018_248, w_018_249, w_018_250, w_018_251, w_018_252, w_018_253, w_018_254, w_018_255, w_018_256, w_018_257, w_018_258, w_018_259, w_018_260, w_018_261, w_018_262, w_018_263, w_018_264, w_018_265, w_018_266, w_018_267, w_018_268, w_018_269, w_018_271, w_018_272, w_018_273, w_018_274, w_018_275, w_018_276, w_018_278, w_018_279, w_018_280, w_018_281, w_018_282;
  wire w_019_000, w_019_001, w_019_002, w_019_005, w_019_010, w_019_011, w_019_014, w_019_019, w_019_020, w_019_021, w_019_023, w_019_024, w_019_025, w_019_027, w_019_028, w_019_030, w_019_031, w_019_032, w_019_040, w_019_055, w_019_058, w_019_062, w_019_071, w_019_074, w_019_077, w_019_080, w_019_081, w_019_082, w_019_083, w_019_085, w_019_089, w_019_090, w_019_091, w_019_092, w_019_097, w_019_099, w_019_101, w_019_105, w_019_106, w_019_110, w_019_113, w_019_115, w_019_122, w_019_123, w_019_124, w_019_127, w_019_128, w_019_130, w_019_132, w_019_133, w_019_135, w_019_139, w_019_141, w_019_142, w_019_144, w_019_145, w_019_150, w_019_151, w_019_152, w_019_153, w_019_161, w_019_164, w_019_165, w_019_167, w_019_176, w_019_183, w_019_188, w_019_189, w_019_190, w_019_191, w_019_192, w_019_201, w_019_202, w_019_204, w_019_205, w_019_206, w_019_209, w_019_212, w_019_213, w_019_216, w_019_219, w_019_220, w_019_222, w_019_225, w_019_229, w_019_230, w_019_232, w_019_234, w_019_237, w_019_239, w_019_240, w_019_244, w_019_246, w_019_250, w_019_252, w_019_253, w_019_257, w_019_259, w_019_262, w_019_269, w_019_273, w_019_277, w_019_278, w_019_279, w_019_284, w_019_287, w_019_288, w_019_289, w_019_290, w_019_292, w_019_294, w_019_296, w_019_297, w_019_298, w_019_302, w_019_303, w_019_304, w_019_305, w_019_310, w_019_317, w_019_326, w_019_328, w_019_329, w_019_331, w_019_338, w_019_339, w_019_340, w_019_342, w_019_343, w_019_344, w_019_347, w_019_350, w_019_353, w_019_358, w_019_359, w_019_360, w_019_361, w_019_365, w_019_368, w_019_369, w_019_374, w_019_377, w_019_383, w_019_385, w_019_386, w_019_387, w_019_389, w_019_391, w_019_395, w_019_397, w_019_401, w_019_402, w_019_404, w_019_405, w_019_406, w_019_407, w_019_409, w_019_411, w_019_415, w_019_416, w_019_417, w_019_419, w_019_420, w_019_423, w_019_428, w_019_430, w_019_436, w_019_437, w_019_438, w_019_439, w_019_441, w_019_445, w_019_449, w_019_450, w_019_451, w_019_459, w_019_463, w_019_465, w_019_467, w_019_470, w_019_474, w_019_476, w_019_478, w_019_480, w_019_481, w_019_482, w_019_485, w_019_486, w_019_487, w_019_488, w_019_491, w_019_494, w_019_499, w_019_500, w_019_504, w_019_505, w_019_507, w_019_512, w_019_514, w_019_516, w_019_519, w_019_521, w_019_524, w_019_525, w_019_526, w_019_527, w_019_530, w_019_537, w_019_538, w_019_543, w_019_544, w_019_545, w_019_547, w_019_551, w_019_552, w_019_553, w_019_556, w_019_558, w_019_559, w_019_560, w_019_563, w_019_568, w_019_569, w_019_571, w_019_573, w_019_575, w_019_577, w_019_580, w_019_583, w_019_585, w_019_586, w_019_590, w_019_593, w_019_595, w_019_596, w_019_597, w_019_598, w_019_599, w_019_601, w_019_604, w_019_608, w_019_610, w_019_613, w_019_614, w_019_615, w_019_617, w_019_618, w_019_619, w_019_625, w_019_627, w_019_629, w_019_631, w_019_632, w_019_633, w_019_637, w_019_643, w_019_647, w_019_648, w_019_655, w_019_656, w_019_657, w_019_659, w_019_665, w_019_666, w_019_668, w_019_671, w_019_673, w_019_675, w_019_682, w_019_689, w_019_691, w_019_692, w_019_695, w_019_699, w_019_700, w_019_701, w_019_702, w_019_705, w_019_706, w_019_707, w_019_709, w_019_710, w_019_717, w_019_718, w_019_721, w_019_722, w_019_723, w_019_724, w_019_726, w_019_729, w_019_732, w_019_745, w_019_748, w_019_753, w_019_754, w_019_755, w_019_756, w_019_757, w_019_761, w_019_763, w_019_766, w_019_770, w_019_771, w_019_772, w_019_773, w_019_775, w_019_776, w_019_778, w_019_782, w_019_783, w_019_784, w_019_786, w_019_790, w_019_791, w_019_797, w_019_800, w_019_808, w_019_812, w_019_814, w_019_815, w_019_817, w_019_819, w_019_825, w_019_831, w_019_834, w_019_836, w_019_842, w_019_843, w_019_844, w_019_845, w_019_849, w_019_858, w_019_859, w_019_860, w_019_864, w_019_865, w_019_866, w_019_868, w_019_876, w_019_877, w_019_879, w_019_881, w_019_882, w_019_888, w_019_890, w_019_893, w_019_894, w_019_897, w_019_898, w_019_900, w_019_905, w_019_908, w_019_909, w_019_917, w_019_918, w_019_920, w_019_926, w_019_951, w_019_953, w_019_958, w_019_960, w_019_962, w_019_965, w_019_968, w_019_975, w_019_978, w_019_980, w_019_994, w_019_1007, w_019_1008, w_019_1017, w_019_1019, w_019_1021, w_019_1022, w_019_1026, w_019_1029, w_019_1031, w_019_1036, w_019_1037, w_019_1040, w_019_1048, w_019_1057, w_019_1059, w_019_1060, w_019_1070, w_019_1073, w_019_1074, w_019_1082, w_019_1084, w_019_1085, w_019_1086, w_019_1089, w_019_1097;
  wire w_020_007, w_020_014, w_020_015, w_020_017, w_020_020, w_020_028, w_020_029, w_020_030, w_020_032, w_020_039, w_020_041, w_020_045, w_020_063, w_020_064, w_020_068, w_020_074, w_020_075, w_020_085, w_020_092, w_020_093, w_020_096, w_020_106, w_020_107, w_020_111, w_020_112, w_020_114, w_020_116, w_020_117, w_020_121, w_020_123, w_020_133, w_020_134, w_020_135, w_020_138, w_020_139, w_020_151, w_020_152, w_020_154, w_020_160, w_020_162, w_020_164, w_020_171, w_020_174, w_020_176, w_020_178, w_020_182, w_020_183, w_020_191, w_020_193, w_020_196, w_020_201, w_020_203, w_020_204, w_020_209, w_020_210, w_020_217, w_020_219, w_020_220, w_020_227, w_020_228, w_020_229, w_020_231, w_020_239, w_020_240, w_020_243, w_020_244, w_020_249, w_020_250, w_020_252, w_020_256, w_020_265, w_020_269, w_020_274, w_020_277, w_020_278, w_020_286, w_020_288, w_020_289, w_020_290, w_020_292, w_020_293, w_020_295, w_020_296, w_020_298, w_020_301, w_020_304, w_020_305, w_020_308, w_020_312, w_020_314, w_020_315, w_020_317, w_020_323, w_020_325, w_020_327, w_020_330, w_020_332, w_020_333, w_020_338, w_020_342, w_020_343, w_020_348, w_020_350, w_020_351, w_020_354, w_020_355, w_020_358, w_020_359, w_020_360, w_020_366, w_020_369, w_020_371, w_020_373, w_020_375, w_020_376, w_020_377, w_020_379, w_020_381, w_020_383, w_020_385, w_020_387, w_020_388, w_020_395, w_020_397, w_020_399, w_020_401, w_020_404, w_020_405, w_020_416, w_020_422, w_020_423, w_020_430, w_020_431, w_020_439, w_020_440, w_020_441, w_020_445, w_020_448, w_020_449, w_020_452, w_020_453, w_020_456, w_020_457, w_020_460, w_020_464, w_020_465, w_020_466, w_020_469, w_020_473, w_020_476, w_020_478, w_020_480, w_020_483, w_020_485, w_020_487, w_020_488, w_020_490, w_020_493, w_020_494, w_020_498, w_020_500, w_020_503, w_020_507, w_020_510, w_020_516, w_020_517, w_020_518, w_020_519, w_020_520, w_020_521, w_020_525, w_020_527, w_020_528, w_020_538, w_020_539, w_020_544, w_020_545, w_020_546, w_020_549, w_020_551, w_020_557, w_020_559, w_020_569, w_020_572, w_020_573, w_020_579, w_020_581, w_020_582, w_020_583, w_020_585, w_020_589, w_020_591, w_020_593, w_020_597, w_020_598, w_020_599, w_020_603, w_020_606, w_020_611, w_020_612, w_020_614, w_020_620, w_020_622, w_020_628, w_020_629, w_020_630, w_020_631, w_020_643, w_020_648, w_020_649, w_020_650, w_020_651, w_020_652, w_020_658, w_020_659, w_020_662, w_020_663, w_020_664, w_020_667, w_020_668, w_020_671, w_020_673, w_020_674, w_020_676, w_020_677, w_020_685, w_020_687, w_020_692, w_020_694, w_020_696, w_020_701, w_020_714, w_020_717, w_020_720, w_020_722, w_020_727, w_020_730, w_020_734, w_020_742, w_020_745, w_020_746, w_020_750, w_020_752, w_020_753, w_020_755, w_020_764, w_020_766, w_020_772, w_020_776, w_020_777, w_020_784, w_020_792, w_020_793, w_020_794, w_020_796, w_020_806, w_020_808, w_020_811, w_020_821, w_020_830, w_020_839, w_020_842, w_020_843, w_020_846, w_020_857, w_020_858, w_020_860, w_020_867, w_020_869, w_020_870, w_020_875, w_020_880, w_020_886, w_020_887, w_020_892, w_020_895, w_020_897, w_020_905, w_020_915, w_020_922, w_020_923, w_020_924, w_020_929, w_020_934, w_020_937, w_020_939, w_020_941, w_020_946, w_020_949, w_020_951, w_020_961, w_020_976, w_020_979, w_020_981, w_020_983, w_020_986, w_020_989, w_020_991, w_020_993, w_020_994, w_020_995, w_020_1001, w_020_1017, w_020_1020, w_020_1021, w_020_1030, w_020_1038, w_020_1040, w_020_1043, w_020_1053, w_020_1060, w_020_1062, w_020_1063, w_020_1068, w_020_1072, w_020_1084, w_020_1085, w_020_1091, w_020_1095, w_020_1097, w_020_1108, w_020_1115, w_020_1120, w_020_1121, w_020_1125, w_020_1129, w_020_1131, w_020_1139, w_020_1143, w_020_1144, w_020_1147, w_020_1151, w_020_1155, w_020_1163, w_020_1166, w_020_1176, w_020_1189, w_020_1191, w_020_1194, w_020_1196, w_020_1198, w_020_1202, w_020_1215, w_020_1219, w_020_1222, w_020_1225, w_020_1235, w_020_1245, w_020_1255, w_020_1258, w_020_1263, w_020_1265;
  wire w_021_000, w_021_001, w_021_002, w_021_003, w_021_005, w_021_006, w_021_007, w_021_009, w_021_010, w_021_011, w_021_013, w_021_015, w_021_016, w_021_018, w_021_019, w_021_020, w_021_021, w_021_022, w_021_023, w_021_024, w_021_025, w_021_026, w_021_027, w_021_028, w_021_033, w_021_034, w_021_035, w_021_036, w_021_037, w_021_041, w_021_042, w_021_044, w_021_045, w_021_046, w_021_047, w_021_048, w_021_049, w_021_050, w_021_051, w_021_053, w_021_054, w_021_055, w_021_057, w_021_058, w_021_060, w_021_061, w_021_063, w_021_064, w_021_065, w_021_066, w_021_068, w_021_069, w_021_071, w_021_072, w_021_073, w_021_074, w_021_075, w_021_076, w_021_077, w_021_078, w_021_079, w_021_080, w_021_081, w_021_082, w_021_083, w_021_084, w_021_085, w_021_086, w_021_087, w_021_088, w_021_089, w_021_090, w_021_091, w_021_092, w_021_093, w_021_094, w_021_095, w_021_096, w_021_097, w_021_099, w_021_100, w_021_101, w_021_102, w_021_103, w_021_104, w_021_105, w_021_107, w_021_111, w_021_112, w_021_115, w_021_116, w_021_117, w_021_118, w_021_119, w_021_120, w_021_122, w_021_123, w_021_124, w_021_126, w_021_128, w_021_129, w_021_130, w_021_132, w_021_134, w_021_135, w_021_136, w_021_137, w_021_138, w_021_139, w_021_140, w_021_141, w_021_142, w_021_143, w_021_144, w_021_145, w_021_147, w_021_148, w_021_149, w_021_150, w_021_151, w_021_153, w_021_154, w_021_155, w_021_156, w_021_157, w_021_158, w_021_159, w_021_161, w_021_162, w_021_163, w_021_166, w_021_167, w_021_169, w_021_171, w_021_172, w_021_174, w_021_177, w_021_179, w_021_180, w_021_182, w_021_184, w_021_185, w_021_186, w_021_187, w_021_189, w_021_191, w_021_193, w_021_194, w_021_195, w_021_198, w_021_199, w_021_201, w_021_202, w_021_203, w_021_204, w_021_205, w_021_207, w_021_208, w_021_210, w_021_211, w_021_212, w_021_214, w_021_216, w_021_218, w_021_220, w_021_221, w_021_223, w_021_224, w_021_225, w_021_226, w_021_227, w_021_228, w_021_229, w_021_231, w_021_232, w_021_233, w_021_234, w_021_235, w_021_236, w_021_237, w_021_238, w_021_239, w_021_240, w_021_241, w_021_242, w_021_244, w_021_245, w_021_246, w_021_248, w_021_249, w_021_250, w_021_251, w_021_253, w_021_254, w_021_255, w_021_256, w_021_257, w_021_258, w_021_259, w_021_260, w_021_261, w_021_262, w_021_263, w_021_264, w_021_265, w_021_266, w_021_268, w_021_269, w_021_270, w_021_271, w_021_272, w_021_273, w_021_274, w_021_275, w_021_276, w_021_277;
  wire w_022_000, w_022_001, w_022_002, w_022_003, w_022_004, w_022_005, w_022_007, w_022_008, w_022_009, w_022_010, w_022_011, w_022_012, w_022_013, w_022_015, w_022_016, w_022_018, w_022_023, w_022_025, w_022_026, w_022_027, w_022_028, w_022_029, w_022_030, w_022_031, w_022_032, w_022_033, w_022_036, w_022_037, w_022_038, w_022_039, w_022_041, w_022_042, w_022_043, w_022_045, w_022_046, w_022_047, w_022_051, w_022_053, w_022_054, w_022_055, w_022_056, w_022_057, w_022_058, w_022_059, w_022_060, w_022_061, w_022_062, w_022_064, w_022_066, w_022_067, w_022_068, w_022_069, w_022_070, w_022_072, w_022_074, w_022_075, w_022_076, w_022_078, w_022_079, w_022_081, w_022_083, w_022_084, w_022_085, w_022_088, w_022_089, w_022_090, w_022_093, w_022_094, w_022_096, w_022_097, w_022_098, w_022_099, w_022_101, w_022_103, w_022_104, w_022_105, w_022_107, w_022_108, w_022_109, w_022_111, w_022_113, w_022_114, w_022_116, w_022_118, w_022_120, w_022_122, w_022_123, w_022_128, w_022_129, w_022_131, w_022_132, w_022_133, w_022_135, w_022_136, w_022_137, w_022_139, w_022_140, w_022_141, w_022_142, w_022_143, w_022_144, w_022_146, w_022_148, w_022_149, w_022_150, w_022_152, w_022_153, w_022_155, w_022_156, w_022_159, w_022_161, w_022_163, w_022_166, w_022_168, w_022_169, w_022_171, w_022_172, w_022_173, w_022_175, w_022_177, w_022_178, w_022_179, w_022_181, w_022_182, w_022_184, w_022_185, w_022_186, w_022_188, w_022_194, w_022_195, w_022_196, w_022_197, w_022_200, w_022_201, w_022_202, w_022_203, w_022_204, w_022_206, w_022_208, w_022_210, w_022_212, w_022_213, w_022_217, w_022_219, w_022_222, w_022_223, w_022_224, w_022_225, w_022_227, w_022_230, w_022_231, w_022_232, w_022_233, w_022_234, w_022_235, w_022_236, w_022_238, w_022_244, w_022_246, w_022_248, w_022_249, w_022_251, w_022_254, w_022_262, w_022_265, w_022_266, w_022_267, w_022_268, w_022_275, w_022_277, w_022_278, w_022_279, w_022_280, w_022_281, w_022_283, w_022_286, w_022_287, w_022_289, w_022_290, w_022_293, w_022_294, w_022_295, w_022_296, w_022_297, w_022_298, w_022_300, w_022_302, w_022_304, w_022_305, w_022_306, w_022_307, w_022_308, w_022_309, w_022_310, w_022_311, w_022_312, w_022_316, w_022_320, w_022_321, w_022_322, w_022_323, w_022_324, w_022_325, w_022_327, w_022_329, w_022_331, w_022_332, w_022_335, w_022_338, w_022_339, w_022_340, w_022_341, w_022_342, w_022_343, w_022_344, w_022_346, w_022_347, w_022_348, w_022_349, w_022_353, w_022_354, w_022_356, w_022_362, w_022_365, w_022_367, w_022_368, w_022_369, w_022_370, w_022_371, w_022_373, w_022_374, w_022_376, w_022_377, w_022_381, w_022_382, w_022_383, w_022_385, w_022_386, w_022_388, w_022_390, w_022_391, w_022_392, w_022_393, w_022_395, w_022_397, w_022_398, w_022_399, w_022_400, w_022_401, w_022_402, w_022_403, w_022_404, w_022_405, w_022_407, w_022_408, w_022_409, w_022_410, w_022_412, w_022_413, w_022_414, w_022_416, w_022_417, w_022_418, w_022_420, w_022_428, w_022_430, w_022_440, w_022_441, w_022_442, w_022_443, w_022_444, w_022_445, w_022_446, w_022_447, w_022_451, w_022_452, w_022_453, w_022_454, w_022_455, w_022_456, w_022_457, w_022_458, w_022_459;
  wire w_023_003, w_023_004, w_023_009, w_023_010, w_023_012, w_023_013, w_023_019, w_023_020, w_023_023, w_023_026, w_023_029, w_023_039, w_023_040, w_023_043, w_023_045, w_023_046, w_023_049, w_023_060, w_023_061, w_023_062, w_023_064, w_023_065, w_023_066, w_023_070, w_023_071, w_023_072, w_023_076, w_023_077, w_023_088, w_023_091, w_023_093, w_023_097, w_023_100, w_023_101, w_023_111, w_023_114, w_023_117, w_023_123, w_023_126, w_023_135, w_023_136, w_023_142, w_023_147, w_023_154, w_023_156, w_023_157, w_023_158, w_023_161, w_023_169, w_023_176, w_023_180, w_023_181, w_023_187, w_023_190, w_023_191, w_023_198, w_023_199, w_023_204, w_023_205, w_023_206, w_023_211, w_023_212, w_023_213, w_023_216, w_023_219, w_023_227, w_023_232, w_023_235, w_023_236, w_023_237, w_023_238, w_023_243, w_023_245, w_023_250, w_023_253, w_023_255, w_023_256, w_023_257, w_023_261, w_023_262, w_023_265, w_023_266, w_023_269, w_023_277, w_023_278, w_023_280, w_023_282, w_023_283, w_023_289, w_023_290, w_023_291, w_023_293, w_023_294, w_023_299, w_023_300, w_023_301, w_023_311, w_023_318, w_023_319, w_023_321, w_023_328, w_023_329, w_023_331, w_023_333, w_023_334, w_023_335, w_023_336, w_023_338, w_023_339, w_023_342, w_023_345, w_023_347, w_023_348, w_023_349, w_023_353, w_023_355, w_023_357, w_023_359, w_023_364, w_023_367, w_023_379, w_023_380, w_023_412, w_023_414, w_023_447, w_023_448, w_023_449, w_023_450, w_023_459, w_023_474, w_023_476, w_023_479, w_023_487, w_023_491, w_023_496, w_023_498, w_023_502, w_023_514, w_023_515, w_023_527, w_023_533, w_023_538, w_023_546, w_023_553, w_023_558, w_023_577, w_023_585, w_023_589, w_023_596, w_023_614, w_023_622, w_023_624, w_023_625, w_023_632, w_023_635, w_023_640, w_023_642, w_023_646, w_023_648, w_023_650, w_023_654, w_023_656, w_023_666, w_023_667, w_023_679, w_023_682, w_023_702, w_023_708, w_023_710, w_023_718, w_023_720, w_023_726, w_023_732, w_023_733, w_023_736, w_023_748, w_023_758, w_023_759, w_023_764, w_023_769, w_023_775, w_023_776, w_023_780, w_023_785, w_023_787, w_023_791, w_023_811, w_023_818, w_023_820, w_023_822, w_023_824, w_023_826, w_023_829, w_023_834, w_023_836, w_023_848, w_023_849, w_023_852, w_023_864, w_023_878, w_023_880, w_023_882, w_023_885, w_023_902, w_023_903, w_023_906, w_023_914, w_023_915, w_023_921, w_023_929, w_023_934, w_023_937, w_023_939, w_023_956, w_023_969, w_023_974, w_023_986, w_023_994, w_023_996, w_023_1004, w_023_1006, w_023_1007, w_023_1013, w_023_1019, w_023_1023, w_023_1026, w_023_1031, w_023_1037, w_023_1043, w_023_1046, w_023_1065, w_023_1068, w_023_1090, w_023_1098, w_023_1105, w_023_1114, w_023_1115, w_023_1116, w_023_1132, w_023_1140, w_023_1141, w_023_1153, w_023_1156, w_023_1163, w_023_1166, w_023_1168, w_023_1179, w_023_1180, w_023_1182, w_023_1194, w_023_1196, w_023_1199, w_023_1200, w_023_1208, w_023_1216, w_023_1218, w_023_1219, w_023_1225, w_023_1226, w_023_1259, w_023_1262, w_023_1265, w_023_1266, w_023_1273, w_023_1275, w_023_1283, w_023_1284, w_023_1292, w_023_1294, w_023_1298, w_023_1313, w_023_1318, w_023_1327, w_023_1336, w_023_1348, w_023_1357, w_023_1363, w_023_1364, w_023_1369, w_023_1371, w_023_1380, w_023_1391, w_023_1396, w_023_1398, w_023_1410, w_023_1412, w_023_1421, w_023_1431, w_023_1439, w_023_1452, w_023_1455, w_023_1460, w_023_1474, w_023_1484, w_023_1494, w_023_1502, w_023_1503, w_023_1507, w_023_1543, w_023_1544, w_023_1545, w_023_1553, w_023_1560, w_023_1567, w_023_1569, w_023_1572, w_023_1573, w_023_1580, w_023_1585, w_023_1594, w_023_1595, w_023_1596, w_023_1598, w_023_1604, w_023_1607, w_023_1608, w_023_1612;
  wire w_024_000, w_024_002, w_024_003, w_024_004, w_024_009, w_024_011, w_024_016, w_024_017, w_024_018, w_024_022, w_024_028, w_024_029, w_024_031, w_024_032, w_024_035, w_024_038, w_024_043, w_024_044, w_024_047, w_024_054, w_024_055, w_024_059, w_024_061, w_024_062, w_024_064, w_024_065, w_024_066, w_024_071, w_024_072, w_024_075, w_024_077, w_024_081, w_024_082, w_024_084, w_024_087, w_024_088, w_024_089, w_024_091, w_024_092, w_024_095, w_024_098, w_024_103, w_024_107, w_024_111, w_024_114, w_024_120, w_024_121, w_024_125, w_024_126, w_024_127, w_024_132, w_024_134, w_024_143, w_024_145, w_024_146, w_024_148, w_024_153, w_024_163, w_024_164, w_024_165, w_024_166, w_024_168, w_024_173, w_024_177, w_024_178, w_024_179, w_024_182, w_024_186, w_024_189, w_024_194, w_024_195, w_024_197, w_024_199, w_024_200, w_024_201, w_024_208, w_024_211, w_024_212, w_024_217, w_024_218, w_024_220, w_024_221, w_024_222, w_024_243, w_024_245, w_024_247, w_024_250, w_024_252, w_024_260, w_024_262, w_024_263, w_024_265, w_024_269, w_024_274, w_024_277, w_024_282, w_024_284, w_024_285, w_024_288, w_024_289, w_024_290, w_024_292, w_024_293, w_024_297, w_024_299, w_024_301, w_024_303, w_024_304, w_024_308, w_024_309, w_024_310, w_024_311, w_024_313, w_024_316, w_024_318, w_024_323, w_024_335, w_024_336, w_024_337, w_024_342, w_024_345, w_024_346, w_024_347, w_024_348, w_024_349, w_024_351, w_024_355, w_024_366, w_024_380, w_024_403, w_024_415, w_024_425, w_024_430, w_024_435, w_024_439, w_024_444, w_024_453, w_024_460, w_024_462, w_024_468, w_024_471, w_024_473, w_024_480, w_024_488, w_024_503, w_024_506, w_024_509, w_024_514, w_024_524, w_024_528, w_024_533, w_024_539, w_024_542, w_024_559, w_024_563, w_024_577, w_024_585, w_024_593, w_024_596, w_024_606, w_024_610, w_024_616, w_024_617, w_024_621, w_024_647, w_024_677, w_024_679, w_024_682, w_024_683, w_024_685, w_024_686, w_024_688, w_024_692, w_024_700, w_024_723, w_024_735, w_024_736, w_024_741, w_024_757, w_024_761, w_024_772, w_024_777, w_024_778, w_024_781, w_024_785, w_024_790, w_024_791, w_024_800, w_024_812, w_024_823, w_024_827, w_024_830, w_024_840, w_024_842, w_024_844, w_024_857, w_024_869, w_024_874, w_024_880, w_024_882, w_024_887, w_024_888, w_024_895, w_024_899, w_024_905, w_024_915, w_024_917, w_024_918, w_024_924, w_024_927, w_024_929, w_024_933, w_024_934, w_024_939, w_024_940, w_024_944, w_024_949, w_024_964, w_024_965, w_024_972, w_024_976, w_024_977, w_024_986, w_024_995, w_024_998, w_024_1001, w_024_1003, w_024_1006, w_024_1009, w_024_1010, w_024_1032, w_024_1050, w_024_1053, w_024_1055, w_024_1059, w_024_1066, w_024_1076, w_024_1079, w_024_1085, w_024_1089, w_024_1094, w_024_1098, w_024_1105, w_024_1121, w_024_1133, w_024_1137, w_024_1164, w_024_1187, w_024_1188, w_024_1190, w_024_1193, w_024_1203, w_024_1221, w_024_1225, w_024_1226, w_024_1230, w_024_1235, w_024_1241, w_024_1244, w_024_1248, w_024_1250, w_024_1261, w_024_1269, w_024_1276, w_024_1297, w_024_1320, w_024_1327, w_024_1341, w_024_1362, w_024_1377, w_024_1383, w_024_1385, w_024_1393, w_024_1399, w_024_1401, w_024_1404, w_024_1408, w_024_1422, w_024_1424, w_024_1430, w_024_1431, w_024_1438, w_024_1465, w_024_1466, w_024_1473, w_024_1478, w_024_1489, w_024_1495, w_024_1498, w_024_1504, w_024_1522, w_024_1523, w_024_1539, w_024_1544, w_024_1545, w_024_1555, w_024_1557, w_024_1561, w_024_1563, w_024_1568, w_024_1569, w_024_1570, w_024_1572, w_024_1576, w_024_1579, w_024_1583, w_024_1590, w_024_1591, w_024_1607, w_024_1615, w_024_1617, w_024_1622, w_024_1623, w_024_1624, w_024_1638, w_024_1640, w_024_1642, w_024_1645, w_024_1649;
  wire w_025_000, w_025_006, w_025_007, w_025_008, w_025_013, w_025_014, w_025_015, w_025_016, w_025_017, w_025_021, w_025_022, w_025_029, w_025_031, w_025_032, w_025_034, w_025_035, w_025_036, w_025_059, w_025_061, w_025_064, w_025_070, w_025_080, w_025_081, w_025_082, w_025_088, w_025_092, w_025_097, w_025_099, w_025_100, w_025_101, w_025_102, w_025_106, w_025_111, w_025_116, w_025_119, w_025_137, w_025_142, w_025_145, w_025_150, w_025_165, w_025_171, w_025_172, w_025_173, w_025_177, w_025_178, w_025_179, w_025_180, w_025_182, w_025_186, w_025_198, w_025_202, w_025_206, w_025_208, w_025_209, w_025_216, w_025_221, w_025_230, w_025_232, w_025_235, w_025_240, w_025_243, w_025_244, w_025_247, w_025_253, w_025_255, w_025_259, w_025_262, w_025_267, w_025_287, w_025_289, w_025_290, w_025_298, w_025_300, w_025_307, w_025_311, w_025_314, w_025_327, w_025_328, w_025_335, w_025_337, w_025_342, w_025_352, w_025_355, w_025_358, w_025_374, w_025_377, w_025_389, w_025_390, w_025_396, w_025_414, w_025_416, w_025_420, w_025_422, w_025_434, w_025_435, w_025_437, w_025_451, w_025_455, w_025_456, w_025_458, w_025_479, w_025_481, w_025_491, w_025_492, w_025_502, w_025_515, w_025_518, w_025_521, w_025_527, w_025_547, w_025_548, w_025_552, w_025_553, w_025_556, w_025_565, w_025_570, w_025_573, w_025_579, w_025_580, w_025_592, w_025_593, w_025_596, w_025_601, w_025_604, w_025_617, w_025_629, w_025_630, w_025_639, w_025_647, w_025_649, w_025_657, w_025_661, w_025_668, w_025_679, w_025_683, w_025_688, w_025_695, w_025_697, w_025_699, w_025_704, w_025_705, w_025_707, w_025_711, w_025_712, w_025_718, w_025_719, w_025_725, w_025_730, w_025_734, w_025_738, w_025_739, w_025_747, w_025_759, w_025_766, w_025_768, w_025_775, w_025_777, w_025_779, w_025_780, w_025_782, w_025_783, w_025_788, w_025_795, w_025_810, w_025_815, w_025_817, w_025_823, w_025_824, w_025_825, w_025_837, w_025_839, w_025_842, w_025_848, w_025_877, w_025_888, w_025_897, w_025_911, w_025_913, w_025_914, w_025_938, w_025_941, w_025_953, w_025_959, w_025_961, w_025_976, w_025_982, w_025_983, w_025_988, w_025_992, w_025_999, w_025_1002, w_025_1004, w_025_1006, w_025_1007, w_025_1025, w_025_1028, w_025_1036, w_025_1037, w_025_1041, w_025_1042, w_025_1047, w_025_1048, w_025_1051, w_025_1053, w_025_1065, w_025_1070, w_025_1079, w_025_1083, w_025_1084, w_025_1085, w_025_1094, w_025_1097, w_025_1120, w_025_1124, w_025_1125, w_025_1126, w_025_1134, w_025_1161, w_025_1164, w_025_1169, w_025_1170, w_025_1174, w_025_1192, w_025_1211, w_025_1222, w_025_1241, w_025_1242, w_025_1243, w_025_1249, w_025_1251, w_025_1258, w_025_1265, w_025_1273, w_025_1280, w_025_1287, w_025_1295, w_025_1304, w_025_1309, w_025_1317, w_025_1321, w_025_1338, w_025_1341, w_025_1350, w_025_1351, w_025_1357, w_025_1374, w_025_1375, w_025_1379, w_025_1391, w_025_1399, w_025_1401, w_025_1406, w_025_1407, w_025_1408, w_025_1412, w_025_1425, w_025_1426, w_025_1432, w_025_1433, w_025_1434, w_025_1441, w_025_1442, w_025_1452, w_025_1456, w_025_1469, w_025_1472, w_025_1476, w_025_1483, w_025_1484, w_025_1495, w_025_1498, w_025_1508, w_025_1520, w_025_1524, w_025_1529, w_025_1533, w_025_1537, w_025_1538, w_025_1540, w_025_1543, w_025_1544, w_025_1549, w_025_1550, w_025_1564, w_025_1572, w_025_1575, w_025_1597, w_025_1611, w_025_1615, w_025_1622, w_025_1626, w_025_1629, w_025_1633, w_025_1651, w_025_1655, w_025_1661, w_025_1668, w_025_1671, w_025_1674, w_025_1675, w_025_1678, w_025_1698, w_025_1703;
  wire w_026_001, w_026_005, w_026_007, w_026_010, w_026_011, w_026_020, w_026_022, w_026_024, w_026_027, w_026_045, w_026_048, w_026_055, w_026_056, w_026_058, w_026_060, w_026_065, w_026_068, w_026_069, w_026_073, w_026_074, w_026_075, w_026_079, w_026_090, w_026_097, w_026_099, w_026_103, w_026_106, w_026_108, w_026_110, w_026_117, w_026_119, w_026_123, w_026_125, w_026_127, w_026_134, w_026_136, w_026_144, w_026_148, w_026_152, w_026_153, w_026_154, w_026_155, w_026_156, w_026_159, w_026_161, w_026_170, w_026_172, w_026_175, w_026_189, w_026_190, w_026_192, w_026_195, w_026_201, w_026_203, w_026_216, w_026_218, w_026_219, w_026_224, w_026_227, w_026_230, w_026_233, w_026_234, w_026_236, w_026_238, w_026_257, w_026_258, w_026_262, w_026_265, w_026_266, w_026_267, w_026_268, w_026_275, w_026_276, w_026_287, w_026_288, w_026_291, w_026_295, w_026_300, w_026_311, w_026_317, w_026_318, w_026_324, w_026_325, w_026_330, w_026_331, w_026_337, w_026_341, w_026_345, w_026_352, w_026_354, w_026_360, w_026_366, w_026_374, w_026_376, w_026_378, w_026_379, w_026_382, w_026_388, w_026_394, w_026_396, w_026_404, w_026_416, w_026_419, w_026_423, w_026_431, w_026_435, w_026_439, w_026_440, w_026_443, w_026_446, w_026_449, w_026_450, w_026_451, w_026_453, w_026_457, w_026_466, w_026_467, w_026_468, w_026_480, w_026_481, w_026_491, w_026_510, w_026_515, w_026_521, w_026_533, w_026_545, w_026_567, w_026_570, w_026_572, w_026_577, w_026_588, w_026_595, w_026_597, w_026_601, w_026_602, w_026_609, w_026_610, w_026_620, w_026_622, w_026_639, w_026_650, w_026_654, w_026_658, w_026_660, w_026_661, w_026_665, w_026_666, w_026_671, w_026_691, w_026_695, w_026_699, w_026_717, w_026_723, w_026_725, w_026_741, w_026_750, w_026_751, w_026_763, w_026_771, w_026_772, w_026_777, w_026_785, w_026_790, w_026_797, w_026_813, w_026_815, w_026_817, w_026_820, w_026_830, w_026_838, w_026_843, w_026_844, w_026_846, w_026_860, w_026_871, w_026_874, w_026_879, w_026_882, w_026_884, w_026_901, w_026_905, w_026_909, w_026_937, w_026_949, w_026_952, w_026_955, w_026_984, w_026_987, w_026_991, w_026_993, w_026_994, w_026_995, w_026_997, w_026_998, w_026_1002, w_026_1006, w_026_1008, w_026_1012, w_026_1016, w_026_1026, w_026_1027, w_026_1028, w_026_1029, w_026_1031, w_026_1035, w_026_1043, w_026_1044, w_026_1048, w_026_1070, w_026_1071, w_026_1072, w_026_1080, w_026_1084, w_026_1094, w_026_1097, w_026_1105, w_026_1107, w_026_1109, w_026_1111, w_026_1112, w_026_1113, w_026_1116, w_026_1123, w_026_1126, w_026_1135, w_026_1136, w_026_1155, w_026_1158, w_026_1159, w_026_1169, w_026_1177, w_026_1178, w_026_1182, w_026_1186, w_026_1201, w_026_1202, w_026_1221, w_026_1223, w_026_1226, w_026_1240, w_026_1243, w_026_1244, w_026_1253, w_026_1257, w_026_1260, w_026_1268, w_026_1274, w_026_1277, w_026_1287, w_026_1289, w_026_1296, w_026_1297, w_026_1304, w_026_1305, w_026_1316, w_026_1325, w_026_1336, w_026_1347, w_026_1356, w_026_1357, w_026_1359, w_026_1365, w_026_1366, w_026_1371, w_026_1376, w_026_1407, w_026_1415, w_026_1418, w_026_1424, w_026_1427, w_026_1429, w_026_1436, w_026_1443, w_026_1448, w_026_1455, w_026_1456, w_026_1463, w_026_1467, w_026_1470, w_026_1483, w_026_1489, w_026_1491, w_026_1507, w_026_1512, w_026_1520;
  wire w_027_001, w_027_003, w_027_006, w_027_007, w_027_008, w_027_011, w_027_012, w_027_013, w_027_014, w_027_016, w_027_017, w_027_018, w_027_019, w_027_028, w_027_029, w_027_032, w_027_033, w_027_038, w_027_040, w_027_041, w_027_043, w_027_044, w_027_048, w_027_052, w_027_054, w_027_057, w_027_059, w_027_061, w_027_062, w_027_063, w_027_065, w_027_067, w_027_069, w_027_074, w_027_076, w_027_077, w_027_079, w_027_081, w_027_082, w_027_091, w_027_093, w_027_097, w_027_102, w_027_105, w_027_107, w_027_108, w_027_109, w_027_110, w_027_114, w_027_117, w_027_120, w_027_122, w_027_129, w_027_130, w_027_132, w_027_143, w_027_144, w_027_145, w_027_146, w_027_147, w_027_149, w_027_150, w_027_155, w_027_157, w_027_158, w_027_159, w_027_160, w_027_161, w_027_163, w_027_167, w_027_172, w_027_174, w_027_175, w_027_176, w_027_178, w_027_180, w_027_182, w_027_183, w_027_184, w_027_186, w_027_187, w_027_190, w_027_198, w_027_199, w_027_201, w_027_203, w_027_204, w_027_207, w_027_209, w_027_210, w_027_211, w_027_214, w_027_215, w_027_218, w_027_219, w_027_220, w_027_226, w_027_229, w_027_231, w_027_236, w_027_237, w_027_242, w_027_243, w_027_246, w_027_247, w_027_249, w_027_258, w_027_261, w_027_272, w_027_276, w_027_277, w_027_279, w_027_280, w_027_286, w_027_287, w_027_288, w_027_297, w_027_301, w_027_303, w_027_308, w_027_318, w_027_319, w_027_322, w_027_323, w_027_326, w_027_328, w_027_334, w_027_335, w_027_344, w_027_345, w_027_347, w_027_348, w_027_351, w_027_356, w_027_362, w_027_364, w_027_366, w_027_370, w_027_371, w_027_374, w_027_376, w_027_380, w_027_383, w_027_384, w_027_387, w_027_389, w_027_393, w_027_394, w_027_395, w_027_396, w_027_397, w_027_398, w_027_403, w_027_407, w_027_408, w_027_409, w_027_411, w_027_413, w_027_414, w_027_417, w_027_419, w_027_421, w_027_422, w_027_427, w_027_429, w_027_430, w_027_436, w_027_437, w_027_440, w_027_443, w_027_444, w_027_447, w_027_451, w_027_456, w_027_458, w_027_459, w_027_460, w_027_461, w_027_465, w_027_467, w_027_469, w_027_470, w_027_472, w_027_475, w_027_476, w_027_481, w_027_482, w_027_493, w_027_496, w_027_498, w_027_507, w_027_509, w_027_512, w_027_513, w_027_516, w_027_521, w_027_523, w_027_524, w_027_529, w_027_530, w_027_531, w_027_533, w_027_536, w_027_543, w_027_547, w_027_550, w_027_552, w_027_553, w_027_556, w_027_558, w_027_560, w_027_563, w_027_564, w_027_565, w_027_567, w_027_571, w_027_572, w_027_574, w_027_575, w_027_578, w_027_579, w_027_580, w_027_583, w_027_584, w_027_585, w_027_587, w_027_588, w_027_590, w_027_591;
  wire w_028_000, w_028_001, w_028_002, w_028_004, w_028_007, w_028_010, w_028_018, w_028_022, w_028_024, w_028_025, w_028_026, w_028_028, w_028_029, w_028_035, w_028_038, w_028_041, w_028_046, w_028_049, w_028_051, w_028_054, w_028_056, w_028_061, w_028_062, w_028_064, w_028_066, w_028_067, w_028_070, w_028_071, w_028_076, w_028_077, w_028_079, w_028_082, w_028_083, w_028_084, w_028_087, w_028_088, w_028_092, w_028_094, w_028_095, w_028_097, w_028_098, w_028_102, w_028_106, w_028_108, w_028_111, w_028_112, w_028_114, w_028_116, w_028_118, w_028_119, w_028_120, w_028_124, w_028_126, w_028_130, w_028_132, w_028_135, w_028_137, w_028_140, w_028_145, w_028_146, w_028_149, w_028_150, w_028_152, w_028_155, w_028_157, w_028_158, w_028_159, w_028_160, w_028_169, w_028_170, w_028_172, w_028_175, w_028_177, w_028_181, w_028_189, w_028_191, w_028_194, w_028_195, w_028_197, w_028_204, w_028_209, w_028_217, w_028_219, w_028_223, w_028_231, w_028_236, w_028_237, w_028_243, w_028_244, w_028_247, w_028_251, w_028_253, w_028_256, w_028_257, w_028_258, w_028_266, w_028_267, w_028_275, w_028_277, w_028_279, w_028_280, w_028_285, w_028_287, w_028_292, w_028_298, w_028_300, w_028_301, w_028_311, w_028_313, w_028_317, w_028_319, w_028_323, w_028_325, w_028_335, w_028_340, w_028_342, w_028_346, w_028_353, w_028_355, w_028_365, w_028_373, w_028_380, w_028_381, w_028_384, w_028_397, w_028_399, w_028_404, w_028_409, w_028_414, w_028_418, w_028_420, w_028_426, w_028_430, w_028_435, w_028_453, w_028_454, w_028_461, w_028_463, w_028_465, w_028_469, w_028_470, w_028_472, w_028_473, w_028_479, w_028_480, w_028_485, w_028_491, w_028_495, w_028_513, w_028_516, w_028_526, w_028_528, w_028_529, w_028_530, w_028_541, w_028_546, w_028_549, w_028_552, w_028_553, w_028_557, w_028_565, w_028_566, w_028_568, w_028_580, w_028_581, w_028_583, w_028_586, w_028_589, w_028_592, w_028_595, w_028_610, w_028_619, w_028_622, w_028_623, w_028_624, w_028_626, w_028_630, w_028_633, w_028_636, w_028_638, w_028_639, w_028_641, w_028_647, w_028_648, w_028_653, w_028_655, w_028_664, w_028_666, w_028_668, w_028_670, w_028_671, w_028_674, w_028_678, w_028_680, w_028_683, w_028_690, w_028_698, w_028_704, w_028_705, w_028_706, w_028_714, w_028_716, w_028_719, w_028_721, w_028_722, w_028_725, w_028_727, w_028_731, w_028_735, w_028_748, w_028_757, w_028_760, w_028_763, w_028_764, w_028_766, w_028_767, w_028_768, w_028_777, w_028_780, w_028_783, w_028_795, w_028_798, w_028_801, w_028_805, w_028_809, w_028_813, w_028_814, w_028_823, w_028_826, w_028_829, w_028_832, w_028_847, w_028_851, w_028_852, w_028_853, w_028_855, w_028_863, w_028_866, w_028_871, w_028_873, w_028_874, w_028_876, w_028_880, w_028_889, w_028_907;
  wire w_029_003, w_029_004, w_029_005, w_029_014, w_029_017, w_029_020, w_029_022, w_029_032, w_029_033, w_029_036, w_029_039, w_029_040, w_029_042, w_029_047, w_029_051, w_029_053, w_029_061, w_029_070, w_029_072, w_029_073, w_029_077, w_029_083, w_029_084, w_029_085, w_029_088, w_029_090, w_029_092, w_029_095, w_029_098, w_029_105, w_029_106, w_029_110, w_029_113, w_029_119, w_029_125, w_029_129, w_029_130, w_029_132, w_029_133, w_029_135, w_029_136, w_029_142, w_029_143, w_029_146, w_029_148, w_029_149, w_029_151, w_029_163, w_029_164, w_029_165, w_029_166, w_029_178, w_029_180, w_029_187, w_029_188, w_029_193, w_029_202, w_029_206, w_029_210, w_029_211, w_029_213, w_029_215, w_029_220, w_029_227, w_029_233, w_029_242, w_029_243, w_029_244, w_029_245, w_029_250, w_029_251, w_029_256, w_029_258, w_029_263, w_029_273, w_029_274, w_029_277, w_029_281, w_029_283, w_029_291, w_029_296, w_029_300, w_029_305, w_029_307, w_029_308, w_029_311, w_029_319, w_029_328, w_029_329, w_029_332, w_029_347, w_029_354, w_029_365, w_029_367, w_029_377, w_029_383, w_029_387, w_029_389, w_029_391, w_029_394, w_029_399, w_029_402, w_029_414, w_029_416, w_029_429, w_029_440, w_029_444, w_029_450, w_029_453, w_029_468, w_029_470, w_029_471, w_029_474, w_029_475, w_029_476, w_029_477, w_029_486, w_029_490, w_029_494, w_029_496, w_029_502, w_029_504, w_029_507, w_029_509, w_029_511, w_029_516, w_029_524, w_029_529, w_029_532, w_029_533, w_029_538, w_029_539, w_029_541, w_029_547, w_029_548, w_029_550, w_029_552, w_029_553, w_029_554, w_029_557, w_029_565, w_029_567, w_029_568, w_029_579, w_029_582, w_029_583, w_029_584, w_029_586, w_029_589, w_029_594, w_029_603, w_029_611, w_029_613, w_029_614, w_029_615, w_029_622, w_029_626, w_029_628, w_029_631, w_029_632, w_029_637, w_029_638, w_029_644, w_029_650, w_029_661, w_029_679, w_029_685, w_029_692, w_029_693, w_029_694, w_029_709, w_029_715, w_029_718, w_029_719, w_029_720, w_029_731, w_029_739, w_029_740, w_029_747, w_029_754, w_029_755, w_029_756, w_029_766, w_029_782, w_029_792, w_029_802, w_029_810, w_029_836, w_029_837, w_029_849, w_029_856, w_029_887, w_029_892, w_029_899, w_029_901, w_029_904, w_029_911, w_029_921, w_029_934, w_029_935, w_029_943, w_029_945, w_029_962, w_029_970, w_029_976, w_029_982, w_029_985, w_029_987, w_029_998, w_029_999, w_029_1002, w_029_1003, w_029_1005, w_029_1006, w_029_1053, w_029_1057, w_029_1059, w_029_1074, w_029_1077, w_029_1087, w_029_1091, w_029_1092, w_029_1106, w_029_1109, w_029_1118, w_029_1124, w_029_1126, w_029_1127, w_029_1129, w_029_1135, w_029_1141, w_029_1142, w_029_1155, w_029_1159, w_029_1170, w_029_1171, w_029_1172, w_029_1176, w_029_1193, w_029_1207, w_029_1210, w_029_1236, w_029_1240, w_029_1244, w_029_1245, w_029_1272, w_029_1276, w_029_1281, w_029_1296, w_029_1328, w_029_1337;
  wire w_030_000, w_030_003, w_030_007, w_030_012, w_030_016, w_030_017, w_030_019, w_030_020, w_030_025, w_030_038, w_030_042, w_030_048, w_030_050, w_030_055, w_030_059, w_030_065, w_030_067, w_030_069, w_030_070, w_030_071, w_030_072, w_030_073, w_030_078, w_030_079, w_030_082, w_030_083, w_030_098, w_030_102, w_030_105, w_030_110, w_030_112, w_030_124, w_030_126, w_030_127, w_030_134, w_030_140, w_030_146, w_030_147, w_030_150, w_030_154, w_030_159, w_030_161, w_030_167, w_030_169, w_030_170, w_030_172, w_030_173, w_030_174, w_030_175, w_030_179, w_030_181, w_030_182, w_030_183, w_030_184, w_030_185, w_030_186, w_030_191, w_030_196, w_030_206, w_030_207, w_030_208, w_030_214, w_030_218, w_030_220, w_030_222, w_030_224, w_030_225, w_030_227, w_030_228, w_030_229, w_030_239, w_030_240, w_030_245, w_030_248, w_030_250, w_030_253, w_030_261, w_030_262, w_030_264, w_030_266, w_030_273, w_030_302, w_030_305, w_030_306, w_030_309, w_030_313, w_030_314, w_030_315, w_030_317, w_030_318, w_030_334, w_030_339, w_030_344, w_030_345, w_030_348, w_030_349, w_030_354, w_030_362, w_030_364, w_030_368, w_030_380, w_030_382, w_030_385, w_030_392, w_030_396, w_030_411, w_030_412, w_030_422, w_030_424, w_030_426, w_030_430, w_030_434, w_030_435, w_030_444, w_030_447, w_030_454, w_030_459, w_030_467, w_030_470, w_030_471, w_030_477, w_030_491, w_030_496, w_030_502, w_030_503, w_030_504, w_030_523, w_030_525, w_030_533, w_030_534, w_030_542, w_030_548, w_030_549, w_030_557, w_030_559, w_030_561, w_030_565, w_030_570, w_030_571, w_030_572, w_030_578, w_030_591, w_030_592, w_030_613, w_030_614, w_030_615, w_030_620, w_030_623, w_030_625, w_030_626, w_030_630, w_030_633, w_030_634, w_030_635, w_030_636, w_030_638, w_030_641, w_030_648, w_030_653, w_030_658, w_030_663, w_030_664, w_030_667, w_030_670, w_030_677, w_030_679, w_030_695, w_030_696, w_030_699, w_030_705, w_030_706, w_030_710, w_030_715, w_030_716, w_030_723, w_030_727, w_030_732, w_030_737, w_030_742, w_030_745, w_030_747, w_030_753, w_030_757, w_030_766, w_030_767, w_030_769, w_030_774, w_030_776, w_030_777, w_030_780, w_030_781, w_030_783, w_030_789, w_030_795, w_030_799, w_030_804, w_030_811, w_030_816, w_030_826, w_030_830, w_030_837, w_030_840, w_030_845, w_030_852;
  wire w_031_003, w_031_004, w_031_012, w_031_016, w_031_021, w_031_027, w_031_037, w_031_038, w_031_039, w_031_040, w_031_050, w_031_051, w_031_052, w_031_054, w_031_057, w_031_061, w_031_062, w_031_076, w_031_078, w_031_087, w_031_091, w_031_092, w_031_100, w_031_102, w_031_111, w_031_113, w_031_116, w_031_117, w_031_123, w_031_134, w_031_136, w_031_137, w_031_145, w_031_150, w_031_152, w_031_153, w_031_159, w_031_184, w_031_194, w_031_201, w_031_210, w_031_217, w_031_226, w_031_228, w_031_229, w_031_246, w_031_248, w_031_250, w_031_252, w_031_256, w_031_260, w_031_265, w_031_270, w_031_274, w_031_279, w_031_284, w_031_287, w_031_289, w_031_292, w_031_296, w_031_300, w_031_306, w_031_308, w_031_312, w_031_315, w_031_330, w_031_333, w_031_337, w_031_340, w_031_341, w_031_343, w_031_349, w_031_350, w_031_351, w_031_356, w_031_357, w_031_359, w_031_366, w_031_370, w_031_378, w_031_384, w_031_385, w_031_387, w_031_389, w_031_394, w_031_395, w_031_398, w_031_404, w_031_409, w_031_422, w_031_425, w_031_429, w_031_449, w_031_456, w_031_457, w_031_465, w_031_468, w_031_476, w_031_480, w_031_485, w_031_492, w_031_495, w_031_500, w_031_502, w_031_509, w_031_510, w_031_511, w_031_513, w_031_515, w_031_517, w_031_521, w_031_529, w_031_536, w_031_546, w_031_564, w_031_575, w_031_576, w_031_587, w_031_594, w_031_597, w_031_609, w_031_610, w_031_611, w_031_617, w_031_619, w_031_620, w_031_625, w_031_631, w_031_634, w_031_635, w_031_643, w_031_645, w_031_647, w_031_658, w_031_662, w_031_674, w_031_676, w_031_684, w_031_697, w_031_704, w_031_712, w_031_713, w_031_715, w_031_718, w_031_724, w_031_726, w_031_733, w_031_743, w_031_744, w_031_750, w_031_752, w_031_753, w_031_762, w_031_766, w_031_770, w_031_777, w_031_778, w_031_781, w_031_786, w_031_789, w_031_814, w_031_815, w_031_819, w_031_820, w_031_825, w_031_827, w_031_828, w_031_842, w_031_847, w_031_848, w_031_852, w_031_853, w_031_861, w_031_864, w_031_874, w_031_917, w_031_925, w_031_934, w_031_937, w_031_949, w_031_963, w_031_974, w_031_981, w_031_983, w_031_985, w_031_988, w_031_990, w_031_1001, w_031_1006, w_031_1019, w_031_1021, w_031_1025, w_031_1026, w_031_1027, w_031_1037, w_031_1045, w_031_1052, w_031_1054, w_031_1065, w_031_1109, w_031_1110, w_031_1126, w_031_1129, w_031_1130;
  wire w_032_000, w_032_001, w_032_002, w_032_003, w_032_004, w_032_005, w_032_009, w_032_011, w_032_012, w_032_013, w_032_015, w_032_018, w_032_019, w_032_020, w_032_021, w_032_023, w_032_025, w_032_026, w_032_027, w_032_028, w_032_029, w_032_030, w_032_031, w_032_032, w_032_035, w_032_036, w_032_037, w_032_038, w_032_039, w_032_042, w_032_043, w_032_045, w_032_046, w_032_048, w_032_050, w_032_051, w_032_052, w_032_053, w_032_054, w_032_056, w_032_057, w_032_058, w_032_059, w_032_061, w_032_065, w_032_066, w_032_067, w_032_068, w_032_069, w_032_072, w_032_073, w_032_075, w_032_077, w_032_080, w_032_081, w_032_084, w_032_086, w_032_087, w_032_089, w_032_090, w_032_091, w_032_092, w_032_095, w_032_098, w_032_099, w_032_101, w_032_102, w_032_103, w_032_105, w_032_106, w_032_108, w_032_111, w_032_112, w_032_116, w_032_118, w_032_119, w_032_122, w_032_126, w_032_127, w_032_130, w_032_131, w_032_132, w_032_134, w_032_135, w_032_138, w_032_140, w_032_141, w_032_142, w_032_144, w_032_146, w_032_147, w_032_148, w_032_150, w_032_152, w_032_153, w_032_154, w_032_155, w_032_156, w_032_158, w_032_160, w_032_163, w_032_164, w_032_165, w_032_167, w_032_169, w_032_170, w_032_173, w_032_175, w_032_176, w_032_179, w_032_180, w_032_182, w_032_185, w_032_187, w_032_190, w_032_193, w_032_194, w_032_195, w_032_196, w_032_197, w_032_199, w_032_201, w_032_202, w_032_206, w_032_208, w_032_210, w_032_211, w_032_212, w_032_215, w_032_216, w_032_218, w_032_222, w_032_223, w_032_224, w_032_225, w_032_227, w_032_231, w_032_232, w_032_233, w_032_234, w_032_235, w_032_236, w_032_237, w_032_239, w_032_241, w_032_244;
  wire w_033_001, w_033_004, w_033_012, w_033_016, w_033_018, w_033_022, w_033_033, w_033_040, w_033_053, w_033_055, w_033_058, w_033_064, w_033_067, w_033_069, w_033_081, w_033_082, w_033_083, w_033_086, w_033_087, w_033_090, w_033_093, w_033_099, w_033_103, w_033_107, w_033_109, w_033_112, w_033_113, w_033_114, w_033_115, w_033_117, w_033_121, w_033_123, w_033_127, w_033_137, w_033_138, w_033_139, w_033_168, w_033_175, w_033_191, w_033_195, w_033_210, w_033_218, w_033_221, w_033_222, w_033_232, w_033_234, w_033_244, w_033_245, w_033_248, w_033_249, w_033_260, w_033_276, w_033_283, w_033_284, w_033_294, w_033_307, w_033_314, w_033_320, w_033_322, w_033_323, w_033_326, w_033_332, w_033_341, w_033_347, w_033_355, w_033_361, w_033_370, w_033_373, w_033_390, w_033_391, w_033_393, w_033_397, w_033_413, w_033_423, w_033_453, w_033_457, w_033_476, w_033_478, w_033_482, w_033_485, w_033_498, w_033_501, w_033_523, w_033_528, w_033_539, w_033_550, w_033_563, w_033_574, w_033_595, w_033_600, w_033_602, w_033_605, w_033_629, w_033_631, w_033_634, w_033_638, w_033_643, w_033_649, w_033_655, w_033_660, w_033_672, w_033_682, w_033_697, w_033_708, w_033_713, w_033_722, w_033_730, w_033_752, w_033_755, w_033_801, w_033_803, w_033_805, w_033_845, w_033_847, w_033_869, w_033_876, w_033_895, w_033_923, w_033_927, w_033_944, w_033_949, w_033_970, w_033_979, w_033_987, w_033_999, w_033_1001, w_033_1015, w_033_1018, w_033_1032, w_033_1033, w_033_1044, w_033_1049, w_033_1060, w_033_1068, w_033_1076, w_033_1077, w_033_1098, w_033_1099, w_033_1104, w_033_1112, w_033_1116, w_033_1136, w_033_1142, w_033_1156, w_033_1187, w_033_1193, w_033_1205, w_033_1210, w_033_1214, w_033_1235, w_033_1239, w_033_1243, w_033_1249, w_033_1268, w_033_1277, w_033_1280, w_033_1284, w_033_1291, w_033_1295, w_033_1305, w_033_1307, w_033_1318, w_033_1324, w_033_1357, w_033_1375, w_033_1376, w_033_1405, w_033_1406, w_033_1409, w_033_1411, w_033_1417, w_033_1421, w_033_1429, w_033_1436, w_033_1438, w_033_1444, w_033_1448, w_033_1461, w_033_1489, w_033_1498, w_033_1507, w_033_1512, w_033_1523, w_033_1524, w_033_1551, w_033_1577, w_033_1605, w_033_1619, w_033_1624, w_033_1634, w_033_1635, w_033_1638, w_033_1643, w_033_1647, w_033_1650;
  wire w_034_006, w_034_007, w_034_009, w_034_011, w_034_016, w_034_022, w_034_031, w_034_034, w_034_044, w_034_057, w_034_061, w_034_066, w_034_067, w_034_072, w_034_074, w_034_079, w_034_083, w_034_089, w_034_090, w_034_099, w_034_104, w_034_109, w_034_114, w_034_115, w_034_116, w_034_121, w_034_122, w_034_125, w_034_130, w_034_133, w_034_134, w_034_140, w_034_144, w_034_145, w_034_161, w_034_166, w_034_178, w_034_182, w_034_185, w_034_189, w_034_196, w_034_199, w_034_201, w_034_203, w_034_204, w_034_205, w_034_213, w_034_214, w_034_216, w_034_225, w_034_226, w_034_227, w_034_241, w_034_245, w_034_248, w_034_252, w_034_254, w_034_268, w_034_269, w_034_273, w_034_274, w_034_276, w_034_281, w_034_289, w_034_292, w_034_297, w_034_300, w_034_305, w_034_308, w_034_309, w_034_314, w_034_315, w_034_316, w_034_322, w_034_323, w_034_328, w_034_329, w_034_330, w_034_336, w_034_339, w_034_345, w_034_347, w_034_350, w_034_351, w_034_354, w_034_358, w_034_363, w_034_368, w_034_369, w_034_371, w_034_372, w_034_376, w_034_377, w_034_378, w_034_379, w_034_382, w_034_391, w_034_398, w_034_400, w_034_403, w_034_404, w_034_405, w_034_406, w_034_407, w_034_410, w_034_412, w_034_415, w_034_416, w_034_418, w_034_419, w_034_420, w_034_422, w_034_424, w_034_430, w_034_433, w_034_434, w_034_439, w_034_441, w_034_442, w_034_452, w_034_459, w_034_460, w_034_462, w_034_463, w_034_471, w_034_475, w_034_476, w_034_486, w_034_488, w_034_494, w_034_498, w_034_500, w_034_504, w_034_506, w_034_511, w_034_513, w_034_521, w_034_526, w_034_527, w_034_528, w_034_545, w_034_551, w_034_555, w_034_557, w_034_558, w_034_559, w_034_563, w_034_564, w_034_566, w_034_568, w_034_569, w_034_570, w_034_575, w_034_577, w_034_578, w_034_582, w_034_583, w_034_584, w_034_585, w_034_590, w_034_592, w_034_595, w_034_599, w_034_607, w_034_608, w_034_610, w_034_612, w_034_613, w_034_620, w_034_621, w_034_630, w_034_649, w_034_653, w_034_657, w_034_664, w_034_665, w_034_669, w_034_674, w_034_677, w_034_680, w_034_686, w_034_690;
  wire w_035_003, w_035_004, w_035_026, w_035_028, w_035_029, w_035_036, w_035_037, w_035_050, w_035_051, w_035_052, w_035_061, w_035_064, w_035_066, w_035_076, w_035_077, w_035_083, w_035_084, w_035_087, w_035_088, w_035_091, w_035_095, w_035_096, w_035_101, w_035_102, w_035_103, w_035_104, w_035_109, w_035_111, w_035_116, w_035_117, w_035_130, w_035_134, w_035_136, w_035_138, w_035_139, w_035_144, w_035_149, w_035_152, w_035_160, w_035_167, w_035_168, w_035_175, w_035_188, w_035_194, w_035_203, w_035_208, w_035_209, w_035_212, w_035_213, w_035_217, w_035_225, w_035_228, w_035_235, w_035_238, w_035_240, w_035_255, w_035_263, w_035_274, w_035_276, w_035_301, w_035_323, w_035_328, w_035_343, w_035_349, w_035_350, w_035_351, w_035_352, w_035_358, w_035_397, w_035_433, w_035_440, w_035_446, w_035_460, w_035_467, w_035_516, w_035_520, w_035_546, w_035_574, w_035_600, w_035_608, w_035_626, w_035_637, w_035_640, w_035_642, w_035_643, w_035_644, w_035_647, w_035_657, w_035_671, w_035_678, w_035_712, w_035_722, w_035_760, w_035_772, w_035_777, w_035_804, w_035_805, w_035_815, w_035_818, w_035_832, w_035_840, w_035_844, w_035_848, w_035_861, w_035_866, w_035_894, w_035_908, w_035_921, w_035_936, w_035_938, w_035_941, w_035_976, w_035_987, w_035_991, w_035_996, w_035_997, w_035_998, w_035_999, w_035_1010, w_035_1016, w_035_1017, w_035_1023, w_035_1037, w_035_1040, w_035_1041, w_035_1053, w_035_1054, w_035_1079, w_035_1098, w_035_1102, w_035_1107, w_035_1112, w_035_1119, w_035_1125, w_035_1135, w_035_1146, w_035_1147, w_035_1176, w_035_1198, w_035_1203, w_035_1226, w_035_1227, w_035_1234, w_035_1255, w_035_1267, w_035_1273, w_035_1281, w_035_1303, w_035_1335, w_035_1357, w_035_1371, w_035_1391, w_035_1397, w_035_1425, w_035_1428, w_035_1431, w_035_1437, w_035_1450, w_035_1464, w_035_1471, w_035_1475, w_035_1484, w_035_1485, w_035_1487, w_035_1502, w_035_1506, w_035_1510, w_035_1513, w_035_1518, w_035_1527, w_035_1530, w_035_1546, w_035_1585, w_035_1596, w_035_1601, w_035_1619, w_035_1621, w_035_1646, w_035_1664, w_035_1671, w_035_1673, w_035_1685, w_035_1707, w_035_1713, w_035_1720;
  wire w_036_018, w_036_025, w_036_029, w_036_032, w_036_033, w_036_037, w_036_045, w_036_047, w_036_049, w_036_056, w_036_071, w_036_079, w_036_085, w_036_101, w_036_107, w_036_114, w_036_123, w_036_124, w_036_133, w_036_137, w_036_143, w_036_147, w_036_148, w_036_149, w_036_151, w_036_161, w_036_166, w_036_169, w_036_170, w_036_173, w_036_179, w_036_180, w_036_194, w_036_196, w_036_199, w_036_200, w_036_206, w_036_207, w_036_218, w_036_222, w_036_226, w_036_238, w_036_252, w_036_255, w_036_256, w_036_258, w_036_272, w_036_273, w_036_281, w_036_282, w_036_283, w_036_297, w_036_310, w_036_319, w_036_322, w_036_323, w_036_337, w_036_353, w_036_355, w_036_361, w_036_369, w_036_374, w_036_375, w_036_379, w_036_390, w_036_398, w_036_405, w_036_408, w_036_435, w_036_441, w_036_450, w_036_451, w_036_452, w_036_454, w_036_456, w_036_481, w_036_482, w_036_486, w_036_488, w_036_492, w_036_493, w_036_495, w_036_496, w_036_505, w_036_513, w_036_525, w_036_538, w_036_543, w_036_577, w_036_580, w_036_585, w_036_589, w_036_594, w_036_596, w_036_650, w_036_652, w_036_657, w_036_692, w_036_696, w_036_697, w_036_702, w_036_712, w_036_713, w_036_723, w_036_728, w_036_764, w_036_778, w_036_781, w_036_786, w_036_790, w_036_803, w_036_813, w_036_815, w_036_826, w_036_837, w_036_842, w_036_850, w_036_866, w_036_875, w_036_880, w_036_895, w_036_914, w_036_924, w_036_937, w_036_939, w_036_953, w_036_965, w_036_972, w_036_978, w_036_982, w_036_992, w_036_1005, w_036_1014, w_036_1023, w_036_1034, w_036_1043, w_036_1049, w_036_1071, w_036_1076, w_036_1104, w_036_1107, w_036_1114, w_036_1115, w_036_1129, w_036_1139, w_036_1140, w_036_1149, w_036_1150, w_036_1153, w_036_1174, w_036_1210, w_036_1217, w_036_1218, w_036_1220, w_036_1222, w_036_1226, w_036_1227, w_036_1234, w_036_1237, w_036_1239, w_036_1273, w_036_1289, w_036_1294, w_036_1306, w_036_1309, w_036_1320, w_036_1325, w_036_1336, w_036_1339, w_036_1341, w_036_1346, w_036_1356, w_036_1366, w_036_1373, w_036_1379, w_036_1397, w_036_1399, w_036_1406, w_036_1426, w_036_1438, w_036_1440, w_036_1454, w_036_1457, w_036_1464, w_036_1473, w_036_1475, w_036_1481, w_036_1493;
  wire w_037_001, w_037_007, w_037_028, w_037_046, w_037_055, w_037_072, w_037_076, w_037_081, w_037_085, w_037_090, w_037_098, w_037_111, w_037_114, w_037_119, w_037_137, w_037_143, w_037_145, w_037_155, w_037_156, w_037_157, w_037_160, w_037_161, w_037_175, w_037_188, w_037_190, w_037_193, w_037_197, w_037_201, w_037_210, w_037_219, w_037_222, w_037_226, w_037_262, w_037_303, w_037_324, w_037_328, w_037_352, w_037_355, w_037_363, w_037_372, w_037_387, w_037_407, w_037_438, w_037_446, w_037_496, w_037_502, w_037_508, w_037_510, w_037_517, w_037_519, w_037_535, w_037_541, w_037_547, w_037_553, w_037_563, w_037_567, w_037_594, w_037_604, w_037_607, w_037_627, w_037_629, w_037_633, w_037_649, w_037_669, w_037_670, w_037_674, w_037_675, w_037_679, w_037_684, w_037_690, w_037_702, w_037_705, w_037_706, w_037_713, w_037_741, w_037_745, w_037_765, w_037_774, w_037_777, w_037_778, w_037_793, w_037_804, w_037_807, w_037_812, w_037_849, w_037_876, w_037_879, w_037_884, w_037_900, w_037_901, w_037_906, w_037_923, w_037_939, w_037_942, w_037_949, w_037_953, w_037_982, w_037_998, w_037_999, w_037_1000, w_037_1035, w_037_1050, w_037_1054, w_037_1076, w_037_1081, w_037_1083, w_037_1084, w_037_1088, w_037_1103, w_037_1106, w_037_1108, w_037_1128, w_037_1132, w_037_1140, w_037_1149, w_037_1177, w_037_1186, w_037_1194, w_037_1210, w_037_1211, w_037_1234, w_037_1238, w_037_1254, w_037_1259, w_037_1278, w_037_1290, w_037_1292, w_037_1307, w_037_1309, w_037_1320, w_037_1329, w_037_1339, w_037_1340, w_037_1343, w_037_1344, w_037_1349, w_037_1357, w_037_1389, w_037_1406, w_037_1421, w_037_1422, w_037_1432, w_037_1441, w_037_1451, w_037_1461, w_037_1462, w_037_1488, w_037_1489, w_037_1494, w_037_1500, w_037_1520, w_037_1528, w_037_1531, w_037_1532, w_037_1541, w_037_1554, w_037_1602, w_037_1625, w_037_1637, w_037_1646, w_037_1656, w_037_1659, w_037_1674, w_037_1676, w_037_1678, w_037_1679, w_037_1689, w_037_1694, w_037_1711, w_037_1730;
  wire w_038_002, w_038_006, w_038_007, w_038_012, w_038_015, w_038_019, w_038_021, w_038_022, w_038_027, w_038_028, w_038_031, w_038_034, w_038_039, w_038_043, w_038_045, w_038_048, w_038_049, w_038_052, w_038_055, w_038_058, w_038_061, w_038_063, w_038_065, w_038_068, w_038_073, w_038_076, w_038_077, w_038_081, w_038_084, w_038_100, w_038_108, w_038_109, w_038_111, w_038_112, w_038_113, w_038_118, w_038_122, w_038_130, w_038_134, w_038_136, w_038_141, w_038_144, w_038_148, w_038_150, w_038_152, w_038_153, w_038_155, w_038_158, w_038_160, w_038_161, w_038_170, w_038_173, w_038_175, w_038_178, w_038_181, w_038_183, w_038_186, w_038_192, w_038_196, w_038_198, w_038_200, w_038_201, w_038_207, w_038_208, w_038_211, w_038_221, w_038_224, w_038_227, w_038_233, w_038_235, w_038_236, w_038_239, w_038_255, w_038_256, w_038_258, w_038_260, w_038_263, w_038_265, w_038_269, w_038_276, w_038_281, w_038_287, w_038_290, w_038_299, w_038_300, w_038_302, w_038_304, w_038_308, w_038_317, w_038_319, w_038_320, w_038_325, w_038_327, w_038_331, w_038_332, w_038_333, w_038_335, w_038_337, w_038_338, w_038_339, w_038_345, w_038_348, w_038_353, w_038_362, w_038_364, w_038_366, w_038_367, w_038_368, w_038_372, w_038_378, w_038_382, w_038_384, w_038_385, w_038_387, w_038_390, w_038_391, w_038_392, w_038_395, w_038_397, w_038_400, w_038_401, w_038_402, w_038_404, w_038_405, w_038_410, w_038_412, w_038_413, w_038_429, w_038_438, w_038_439, w_038_448, w_038_451, w_038_454, w_038_457, w_038_458, w_038_459, w_038_464, w_038_473, w_038_475, w_038_479, w_038_480, w_038_484, w_038_485, w_038_486;
  wire w_039_007, w_039_018, w_039_024, w_039_025, w_039_027, w_039_033, w_039_065, w_039_075, w_039_087, w_039_092, w_039_100, w_039_113, w_039_133, w_039_135, w_039_142, w_039_167, w_039_178, w_039_198, w_039_199, w_039_204, w_039_250, w_039_252, w_039_259, w_039_260, w_039_266, w_039_272, w_039_289, w_039_306, w_039_310, w_039_313, w_039_347, w_039_351, w_039_415, w_039_429, w_039_466, w_039_470, w_039_477, w_039_482, w_039_490, w_039_501, w_039_507, w_039_516, w_039_526, w_039_530, w_039_533, w_039_558, w_039_568, w_039_595, w_039_597, w_039_599, w_039_610, w_039_612, w_039_614, w_039_618, w_039_629, w_039_631, w_039_648, w_039_650, w_039_665, w_039_676, w_039_687, w_039_707, w_039_714, w_039_721, w_039_726, w_039_752, w_039_759, w_039_775, w_039_782, w_039_788, w_039_793, w_039_805, w_039_834, w_039_835, w_039_842, w_039_847, w_039_879, w_039_881, w_039_895, w_039_910, w_039_915, w_039_932, w_039_933, w_039_936, w_039_938, w_039_969, w_039_977, w_039_1009, w_039_1059, w_039_1065, w_039_1078, w_039_1097, w_039_1126, w_039_1145, w_039_1151, w_039_1162, w_039_1213, w_039_1227, w_039_1232, w_039_1235, w_039_1273, w_039_1280, w_039_1295, w_039_1297, w_039_1308, w_039_1311, w_039_1335, w_039_1361, w_039_1362, w_039_1372, w_039_1392, w_039_1407, w_039_1446, w_039_1457, w_039_1470, w_039_1496, w_039_1509, w_039_1530, w_039_1548, w_039_1551, w_039_1577, w_039_1582, w_039_1588, w_039_1597, w_039_1600, w_039_1605, w_039_1611, w_039_1634, w_039_1643, w_039_1654, w_039_1699, w_039_1726, w_039_1731, w_039_1753, w_039_1768, w_039_1770, w_039_1788, w_039_1835, w_039_1836, w_039_1856, w_039_1869, w_039_1890, w_039_1891, w_039_1906, w_039_1907, w_039_1919, w_039_1932;
  wire w_040_011, w_040_015, w_040_016, w_040_019, w_040_020, w_040_024, w_040_030, w_040_037, w_040_044, w_040_048, w_040_052, w_040_055, w_040_056, w_040_059, w_040_060, w_040_061, w_040_068, w_040_075, w_040_080, w_040_086, w_040_093, w_040_096, w_040_102, w_040_121, w_040_127, w_040_134, w_040_148, w_040_165, w_040_172, w_040_183, w_040_189, w_040_203, w_040_208, w_040_210, w_040_212, w_040_220, w_040_225, w_040_226, w_040_227, w_040_239, w_040_255, w_040_260, w_040_272, w_040_273, w_040_278, w_040_294, w_040_297, w_040_306, w_040_307, w_040_312, w_040_314, w_040_315, w_040_320, w_040_323, w_040_324, w_040_325, w_040_333, w_040_353, w_040_356, w_040_364, w_040_365, w_040_380, w_040_387, w_040_390, w_040_407, w_040_411, w_040_423, w_040_427, w_040_436, w_040_447, w_040_461, w_040_462, w_040_463, w_040_468, w_040_472, w_040_473, w_040_482, w_040_489, w_040_495, w_040_512, w_040_521, w_040_526, w_040_527, w_040_539, w_040_568, w_040_577, w_040_583, w_040_585, w_040_590, w_040_593, w_040_632, w_040_663, w_040_667, w_040_673, w_040_679, w_040_683, w_040_695, w_040_700, w_040_724, w_040_729, w_040_737, w_040_754, w_040_757, w_040_759, w_040_764, w_040_766, w_040_770, w_040_771, w_040_791, w_040_813, w_040_823, w_040_832, w_040_848, w_040_852, w_040_854, w_040_856, w_040_869, w_040_904, w_040_911, w_040_914, w_040_938, w_040_959, w_040_978, w_040_979, w_040_981, w_040_984, w_040_987, w_040_1003, w_040_1005, w_040_1013, w_040_1028, w_040_1038, w_040_1046, w_040_1076, w_040_1082, w_040_1084, w_040_1102, w_040_1119, w_040_1125, w_040_1134, w_040_1138, w_040_1156, w_040_1178, w_040_1195, w_040_1213, w_040_1232, w_040_1237, w_040_1263, w_040_1276, w_040_1286, w_040_1291, w_040_1294, w_040_1304, w_040_1314, w_040_1320, w_040_1327, w_040_1350, w_040_1352, w_040_1383;
  wire w_041_002, w_041_004, w_041_007, w_041_008, w_041_010, w_041_012, w_041_017, w_041_018, w_041_021, w_041_022, w_041_025, w_041_026, w_041_035, w_041_037, w_041_042, w_041_043, w_041_044, w_041_045, w_041_049, w_041_052, w_041_053, w_041_055, w_041_059, w_041_062, w_041_063, w_041_064, w_041_065, w_041_066, w_041_069, w_041_071, w_041_073, w_041_074, w_041_077, w_041_081, w_041_082, w_041_084, w_041_085, w_041_087, w_041_090, w_041_091, w_041_092, w_041_096, w_041_098, w_041_107, w_041_108, w_041_110, w_041_111, w_041_113, w_041_114, w_041_115, w_041_118, w_041_121, w_041_122, w_041_124, w_041_126, w_041_127, w_041_128, w_041_131, w_041_132, w_041_134, w_041_140, w_041_146, w_041_149, w_041_150, w_041_152, w_041_154, w_041_155, w_041_156, w_041_157, w_041_158, w_041_161, w_041_169, w_041_171, w_041_178, w_041_180, w_041_181, w_041_183, w_041_186, w_041_187, w_041_188, w_041_191, w_041_193, w_041_194, w_041_197, w_041_198, w_041_199, w_041_200, w_041_201, w_041_202, w_041_204, w_041_205, w_041_206, w_041_207, w_041_208, w_041_211, w_041_212, w_041_217, w_041_219, w_041_229, w_041_230, w_041_231, w_041_232, w_041_235, w_041_237, w_041_245, w_041_246, w_041_247, w_041_248, w_041_249, w_041_250, w_041_253, w_041_254, w_041_257, w_041_258, w_041_264, w_041_265, w_041_267, w_041_268, w_041_271, w_041_273, w_041_275, w_041_278, w_041_279, w_041_282, w_041_285, w_041_288, w_041_289, w_041_294;
  wire w_042_000, w_042_001, w_042_002, w_042_003, w_042_007, w_042_008, w_042_009, w_042_014, w_042_016, w_042_017, w_042_018, w_042_019, w_042_021, w_042_022, w_042_023, w_042_025, w_042_026, w_042_027, w_042_028, w_042_029, w_042_030, w_042_031, w_042_034, w_042_035, w_042_036, w_042_037, w_042_040, w_042_041, w_042_044, w_042_046, w_042_047, w_042_048, w_042_051, w_042_052, w_042_053, w_042_054, w_042_055, w_042_058, w_042_060, w_042_062, w_042_063, w_042_064, w_042_065, w_042_068, w_042_072, w_042_073, w_042_074, w_042_076, w_042_077, w_042_079, w_042_081, w_042_084, w_042_085, w_042_086, w_042_088, w_042_089, w_042_093, w_042_094, w_042_095, w_042_096, w_042_097, w_042_100, w_042_102, w_042_103, w_042_104, w_042_105, w_042_107, w_042_109, w_042_110, w_042_111, w_042_112, w_042_113, w_042_115, w_042_117, w_042_118, w_042_119, w_042_121, w_042_122, w_042_124, w_042_125, w_042_127, w_042_128, w_042_129, w_042_130, w_042_132, w_042_134, w_042_135, w_042_137, w_042_139, w_042_140, w_042_141, w_042_142;
  wire w_043_000, w_043_001, w_043_004, w_043_005, w_043_006, w_043_010, w_043_011, w_043_012, w_043_013, w_043_014, w_043_015, w_043_016, w_043_019, w_043_020, w_043_021, w_043_022, w_043_023, w_043_024, w_043_025, w_043_026, w_043_027, w_043_028, w_043_029, w_043_030, w_043_031, w_043_032, w_043_034, w_043_035, w_043_036, w_043_037, w_043_039, w_043_040, w_043_041, w_043_042, w_043_043, w_043_046, w_043_048, w_043_049, w_043_050, w_043_051, w_043_052, w_043_053, w_043_054, w_043_055, w_043_056, w_043_057, w_043_058, w_043_059, w_043_060, w_043_062, w_043_063, w_043_064, w_043_065, w_043_066, w_043_067, w_043_068, w_043_070, w_043_071, w_043_073, w_043_075, w_043_077, w_043_078, w_043_079, w_043_081, w_043_082, w_043_083, w_043_084, w_043_085, w_043_088, w_043_089, w_043_091, w_043_092, w_043_093, w_043_094, w_043_095, w_043_096, w_043_097, w_043_098, w_043_099, w_043_100, w_043_101, w_043_102, w_043_103, w_043_105;
  wire w_044_018, w_044_022, w_044_030, w_044_033, w_044_035, w_044_047, w_044_056, w_044_074, w_044_087, w_044_107, w_044_112, w_044_115, w_044_129, w_044_132, w_044_134, w_044_137, w_044_142, w_044_147, w_044_156, w_044_166, w_044_175, w_044_176, w_044_184, w_044_189, w_044_196, w_044_199, w_044_201, w_044_226, w_044_264, w_044_308, w_044_309, w_044_314, w_044_324, w_044_342, w_044_355, w_044_357, w_044_374, w_044_390, w_044_393, w_044_414, w_044_443, w_044_462, w_044_465, w_044_466, w_044_475, w_044_538, w_044_541, w_044_542, w_044_569, w_044_607, w_044_613, w_044_618, w_044_665, w_044_675, w_044_682, w_044_697, w_044_718, w_044_724, w_044_764, w_044_777, w_044_778, w_044_784, w_044_788, w_044_790, w_044_791, w_044_794, w_044_795, w_044_831, w_044_870, w_044_897, w_044_907, w_044_908, w_044_913, w_044_914, w_044_931, w_044_951, w_044_954, w_044_963, w_044_972, w_044_990, w_044_1077, w_044_1093, w_044_1095, w_044_1108, w_044_1116, w_044_1117, w_044_1134, w_044_1139, w_044_1141, w_044_1146, w_044_1152, w_044_1176, w_044_1197, w_044_1209, w_044_1217, w_044_1224, w_044_1230, w_044_1251, w_044_1261, w_044_1268, w_044_1274, w_044_1327, w_044_1330, w_044_1342, w_044_1344, w_044_1377, w_044_1379, w_044_1383, w_044_1386, w_044_1405, w_044_1417, w_044_1426, w_044_1427, w_044_1446, w_044_1447, w_044_1459, w_044_1465, w_044_1481, w_044_1505, w_044_1523, w_044_1550, w_044_1566, w_044_1580, w_044_1614, w_044_1616, w_044_1629, w_044_1630, w_044_1635, w_044_1639, w_044_1684, w_044_1690, w_044_1695, w_044_1723, w_044_1750, w_044_1751, w_044_1752, w_044_1769, w_044_1781, w_044_1783, w_044_1792;
  wire w_045_005, w_045_009, w_045_023, w_045_041, w_045_065, w_045_066, w_045_070, w_045_072, w_045_077, w_045_082, w_045_093, w_045_110, w_045_163, w_045_170, w_045_171, w_045_199, w_045_209, w_045_213, w_045_224, w_045_226, w_045_251, w_045_255, w_045_266, w_045_288, w_045_290, w_045_303, w_045_310, w_045_331, w_045_335, w_045_338, w_045_344, w_045_346, w_045_365, w_045_398, w_045_405, w_045_424, w_045_437, w_045_452, w_045_475, w_045_483, w_045_490, w_045_495, w_045_524, w_045_547, w_045_548, w_045_574, w_045_578, w_045_580, w_045_583, w_045_588, w_045_599, w_045_607, w_045_617, w_045_635, w_045_662, w_045_666, w_045_710, w_045_711, w_045_721, w_045_731, w_045_747, w_045_752, w_045_766, w_045_786, w_045_796, w_045_802, w_045_805, w_045_830, w_045_874, w_045_937, w_045_957, w_045_962, w_045_1002, w_045_1015, w_045_1052, w_045_1064, w_045_1066, w_045_1071, w_045_1086, w_045_1102, w_045_1104, w_045_1139, w_045_1153, w_045_1161, w_045_1181, w_045_1189, w_045_1203, w_045_1229, w_045_1231, w_045_1242, w_045_1264, w_045_1313, w_045_1328, w_045_1333, w_045_1349, w_045_1414, w_045_1467, w_045_1486, w_045_1488, w_045_1489, w_045_1507, w_045_1538, w_045_1551, w_045_1561, w_045_1590, w_045_1596, w_045_1599, w_045_1622, w_045_1646, w_045_1650, w_045_1653, w_045_1659, w_045_1677, w_045_1693, w_045_1704, w_045_1715, w_045_1718, w_045_1738, w_045_1756, w_045_1806, w_045_1824, w_045_1830, w_045_1833, w_045_1878;
  wire w_046_005, w_046_008, w_046_011, w_046_012, w_046_014, w_046_017, w_046_018, w_046_020, w_046_028, w_046_029, w_046_030, w_046_034, w_046_040, w_046_042, w_046_045, w_046_048, w_046_049, w_046_052, w_046_054, w_046_056, w_046_060, w_046_062, w_046_066, w_046_070, w_046_072, w_046_074, w_046_075, w_046_076, w_046_077, w_046_078, w_046_079, w_046_082, w_046_083, w_046_087, w_046_090, w_046_098, w_046_099, w_046_105, w_046_109, w_046_114, w_046_118, w_046_119, w_046_120, w_046_121, w_046_122, w_046_123, w_046_124, w_046_127, w_046_128, w_046_130, w_046_131, w_046_133, w_046_134, w_046_136, w_046_138, w_046_139, w_046_140, w_046_145, w_046_147, w_046_148, w_046_149, w_046_156, w_046_159, w_046_168, w_046_170, w_046_171, w_046_173, w_046_174, w_046_178, w_046_180, w_046_181, w_046_191, w_046_192, w_046_193, w_046_195, w_046_198, w_046_202, w_046_203, w_046_207, w_046_208, w_046_213, w_046_215, w_046_216, w_046_218, w_046_219, w_046_220, w_046_223, w_046_225, w_046_226, w_046_228, w_046_230, w_046_231, w_046_232, w_046_233, w_046_236, w_046_237, w_046_238, w_046_247, w_046_248, w_046_250, w_046_251, w_046_252, w_046_254, w_046_255, w_046_258, w_046_259, w_046_266, w_046_267, w_046_270, w_046_274, w_046_276, w_046_277, w_046_278, w_046_279, w_046_280, w_046_282;
  wire w_047_000, w_047_007, w_047_013, w_047_015, w_047_019, w_047_022, w_047_028, w_047_031, w_047_046, w_047_054, w_047_056, w_047_057, w_047_059, w_047_060, w_047_062, w_047_065, w_047_073, w_047_074, w_047_100, w_047_103, w_047_107, w_047_115, w_047_119, w_047_129, w_047_139, w_047_140, w_047_141, w_047_149, w_047_174, w_047_175, w_047_190, w_047_194, w_047_195, w_047_196, w_047_224, w_047_226, w_047_230, w_047_231, w_047_233, w_047_235, w_047_241, w_047_251, w_047_253, w_047_259, w_047_262, w_047_280, w_047_283, w_047_288, w_047_291, w_047_301, w_047_303, w_047_319, w_047_320, w_047_329, w_047_331, w_047_332, w_047_335, w_047_338, w_047_340, w_047_341, w_047_345, w_047_362, w_047_363, w_047_372, w_047_375, w_047_384, w_047_386, w_047_387, w_047_391, w_047_400, w_047_404, w_047_415, w_047_418, w_047_419, w_047_425, w_047_428, w_047_434, w_047_441, w_047_442, w_047_462, w_047_465, w_047_475, w_047_480, w_047_489, w_047_491, w_047_496, w_047_500, w_047_501, w_047_503, w_047_518, w_047_524, w_047_532, w_047_537, w_047_543, w_047_545, w_047_548, w_047_550, w_047_552, w_047_558, w_047_562, w_047_568, w_047_569, w_047_570, w_047_573, w_047_577, w_047_579, w_047_585, w_047_594, w_047_595, w_047_599, w_047_606, w_047_632, w_047_639, w_047_640, w_047_641, w_047_653, w_047_675, w_047_692, w_047_698;
  wire w_048_000, w_048_007, w_048_010, w_048_018, w_048_021, w_048_033, w_048_053, w_048_054, w_048_057, w_048_072, w_048_073, w_048_077, w_048_090, w_048_092, w_048_098, w_048_117, w_048_132, w_048_134, w_048_135, w_048_142, w_048_148, w_048_159, w_048_162, w_048_171, w_048_194, w_048_202, w_048_204, w_048_209, w_048_213, w_048_229, w_048_230, w_048_236, w_048_243, w_048_250, w_048_253, w_048_276, w_048_312, w_048_317, w_048_326, w_048_328, w_048_345, w_048_348, w_048_354, w_048_358, w_048_373, w_048_383, w_048_405, w_048_406, w_048_409, w_048_415, w_048_416, w_048_421, w_048_431, w_048_432, w_048_436, w_048_439, w_048_440, w_048_446, w_048_447, w_048_472, w_048_473, w_048_479, w_048_487, w_048_520, w_048_527, w_048_536, w_048_546, w_048_548, w_048_551, w_048_553, w_048_554, w_048_560, w_048_561, w_048_564, w_048_567, w_048_583, w_048_584, w_048_588, w_048_593, w_048_597, w_048_598, w_048_622, w_048_623, w_048_627, w_048_629, w_048_637, w_048_649, w_048_651, w_048_652, w_048_668, w_048_671, w_048_672, w_048_676, w_048_677, w_048_694, w_048_705, w_048_713, w_048_724, w_048_742, w_048_746, w_048_751, w_048_752, w_048_758, w_048_762, w_048_770, w_048_777, w_048_781, w_048_783, w_048_787, w_048_792, w_048_797, w_048_799, w_048_802, w_048_824, w_048_827, w_048_849, w_048_850, w_048_881, w_048_884, w_048_897, w_048_901, w_048_904, w_048_908, w_048_909, w_048_918, w_048_963, w_048_966, w_048_974;
  wire w_049_008, w_049_013, w_049_020, w_049_031, w_049_043, w_049_047, w_049_055, w_049_076, w_049_077, w_049_080, w_049_087, w_049_095, w_049_099, w_049_110, w_049_112, w_049_132, w_049_157, w_049_169, w_049_190, w_049_206, w_049_213, w_049_220, w_049_241, w_049_252, w_049_253, w_049_255, w_049_260, w_049_272, w_049_275, w_049_277, w_049_282, w_049_289, w_049_300, w_049_306, w_049_309, w_049_311, w_049_315, w_049_327, w_049_335, w_049_336, w_049_345, w_049_347, w_049_370, w_049_377, w_049_378, w_049_393, w_049_403, w_049_404, w_049_429, w_049_433, w_049_447, w_049_454, w_049_457, w_049_488, w_049_489, w_049_494, w_049_515, w_049_519, w_049_521, w_049_529, w_049_530, w_049_537, w_049_541, w_049_542, w_049_543, w_049_548, w_049_554, w_049_571, w_049_584, w_049_594, w_049_595, w_049_601, w_049_606, w_049_616, w_049_620, w_049_634, w_049_651, w_049_700, w_049_710, w_049_738, w_049_786, w_049_803, w_049_813, w_049_869, w_049_871, w_049_882, w_049_909, w_049_929, w_049_962, w_049_971, w_049_999, w_049_1001, w_049_1006, w_049_1033, w_049_1041, w_049_1057, w_049_1058, w_049_1067, w_049_1075, w_049_1111, w_049_1129, w_049_1136, w_049_1140, w_049_1143, w_049_1157, w_049_1165, w_049_1167, w_049_1169, w_049_1207, w_049_1221, w_049_1227, w_049_1243, w_049_1303, w_049_1320, w_049_1359;
  wire w_050_010, w_050_015, w_050_016, w_050_020, w_050_032, w_050_033, w_050_038, w_050_041, w_050_044, w_050_045, w_050_052, w_050_066, w_050_069, w_050_071, w_050_079, w_050_090, w_050_097, w_050_101, w_050_102, w_050_105, w_050_154, w_050_155, w_050_161, w_050_162, w_050_169, w_050_174, w_050_175, w_050_176, w_050_181, w_050_185, w_050_190, w_050_191, w_050_193, w_050_197, w_050_217, w_050_220, w_050_225, w_050_257, w_050_266, w_050_275, w_050_276, w_050_314, w_050_321, w_050_322, w_050_326, w_050_342, w_050_352, w_050_353, w_050_354, w_050_362, w_050_367, w_050_368, w_050_370, w_050_380, w_050_382, w_050_383, w_050_393, w_050_395, w_050_406, w_050_418, w_050_420, w_050_435, w_050_438, w_050_448, w_050_462, w_050_468, w_050_499, w_050_502, w_050_552, w_050_556, w_050_562, w_050_565, w_050_597, w_050_610, w_050_614, w_050_671, w_050_683, w_050_686, w_050_715, w_050_718, w_050_731, w_050_749, w_050_751, w_050_760, w_050_764, w_050_802, w_050_814, w_050_819, w_050_855, w_050_875, w_050_897, w_050_961, w_050_967, w_050_972, w_050_994, w_050_1020, w_050_1023, w_050_1045, w_050_1052, w_050_1057, w_050_1082, w_050_1088, w_050_1119, w_050_1147, w_050_1148, w_050_1158, w_050_1164, w_050_1200, w_050_1218, w_050_1224, w_050_1231, w_050_1239, w_050_1244, w_050_1293, w_050_1319, w_050_1344, w_050_1369, w_050_1374, w_050_1379, w_050_1383, w_050_1390, w_050_1394, w_050_1397, w_050_1398, w_050_1405, w_050_1433, w_050_1435, w_050_1452, w_050_1469, w_050_1499, w_050_1537;
  wire w_051_020, w_051_022, w_051_023, w_051_026, w_051_027, w_051_046, w_051_074, w_051_108, w_051_121, w_051_126, w_051_127, w_051_143, w_051_149, w_051_184, w_051_190, w_051_198, w_051_202, w_051_209, w_051_210, w_051_230, w_051_246, w_051_252, w_051_265, w_051_268, w_051_273, w_051_274, w_051_285, w_051_290, w_051_291, w_051_292, w_051_294, w_051_310, w_051_347, w_051_382, w_051_407, w_051_422, w_051_425, w_051_431, w_051_440, w_051_455, w_051_469, w_051_480, w_051_501, w_051_559, w_051_563, w_051_571, w_051_576, w_051_580, w_051_581, w_051_582, w_051_595, w_051_621, w_051_628, w_051_633, w_051_638, w_051_640, w_051_643, w_051_649, w_051_653, w_051_670, w_051_673, w_051_675, w_051_701, w_051_702, w_051_703, w_051_710, w_051_714, w_051_735, w_051_768, w_051_773, w_051_777, w_051_783, w_051_804, w_051_812, w_051_828, w_051_837, w_051_847, w_051_849, w_051_853, w_051_868, w_051_881, w_051_891, w_051_939, w_051_947, w_051_958, w_051_960, w_051_982, w_051_992, w_051_996, w_051_1001, w_051_1012, w_051_1015, w_051_1022, w_051_1023, w_051_1044, w_051_1064, w_051_1068, w_051_1073, w_051_1092;
  wire w_052_011, w_052_016, w_052_017, w_052_031, w_052_034, w_052_037, w_052_042, w_052_047, w_052_058, w_052_059, w_052_061, w_052_145, w_052_166, w_052_173, w_052_185, w_052_198, w_052_205, w_052_218, w_052_242, w_052_266, w_052_309, w_052_338, w_052_382, w_052_388, w_052_391, w_052_392, w_052_405, w_052_432, w_052_440, w_052_461, w_052_465, w_052_498, w_052_503, w_052_547, w_052_566, w_052_574, w_052_587, w_052_640, w_052_667, w_052_711, w_052_715, w_052_731, w_052_733, w_052_743, w_052_817, w_052_825, w_052_844, w_052_853, w_052_857, w_052_877, w_052_904, w_052_925, w_052_947, w_052_952, w_052_965, w_052_981, w_052_987, w_052_1001, w_052_1038, w_052_1058, w_052_1072, w_052_1104, w_052_1110, w_052_1126, w_052_1133, w_052_1203, w_052_1220, w_052_1247, w_052_1248, w_052_1264, w_052_1284, w_052_1289, w_052_1295, w_052_1299, w_052_1301, w_052_1304, w_052_1323, w_052_1331, w_052_1340, w_052_1341, w_052_1364, w_052_1375, w_052_1379, w_052_1394, w_052_1396, w_052_1437, w_052_1458, w_052_1482, w_052_1525, w_052_1549, w_052_1554, w_052_1564, w_052_1566, w_052_1573, w_052_1588, w_052_1598, w_052_1601, w_052_1621, w_052_1682, w_052_1690, w_052_1709, w_052_1721, w_052_1771, w_052_1783, w_052_1785, w_052_1792, w_052_1801, w_052_1844, w_052_1856, w_052_1875, w_052_1907, w_052_1918;
  wire w_053_000, w_053_001, w_053_003, w_053_004, w_053_005, w_053_007, w_053_011, w_053_012, w_053_013, w_053_014, w_053_016, w_053_017, w_053_018, w_053_019, w_053_023, w_053_024, w_053_028, w_053_029, w_053_031, w_053_032, w_053_033, w_053_034, w_053_035, w_053_036, w_053_040, w_053_042, w_053_043, w_053_044, w_053_045, w_053_047, w_053_048, w_053_049, w_053_050, w_053_053, w_053_060, w_053_063, w_053_064, w_053_068, w_053_069, w_053_071, w_053_073, w_053_076, w_053_077, w_053_080, w_053_083, w_053_084, w_053_085, w_053_087, w_053_089, w_053_091, w_053_092, w_053_095, w_053_096, w_053_098, w_053_103, w_053_104, w_053_105, w_053_106, w_053_107, w_053_108, w_053_109, w_053_110, w_053_114, w_053_116, w_053_117, w_053_118, w_053_120, w_053_121;
  wire w_054_003, w_054_007, w_054_016, w_054_036, w_054_042, w_054_052, w_054_057, w_054_060, w_054_065, w_054_073, w_054_079, w_054_086, w_054_095, w_054_102, w_054_103, w_054_117, w_054_158, w_054_166, w_054_170, w_054_172, w_054_180, w_054_186, w_054_188, w_054_193, w_054_204, w_054_220, w_054_233, w_054_238, w_054_251, w_054_269, w_054_275, w_054_286, w_054_299, w_054_300, w_054_303, w_054_308, w_054_313, w_054_315, w_054_320, w_054_332, w_054_334, w_054_343, w_054_352, w_054_353, w_054_355, w_054_365, w_054_366, w_054_382, w_054_390, w_054_399, w_054_401, w_054_411, w_054_413, w_054_414, w_054_432, w_054_437, w_054_440, w_054_444, w_054_469, w_054_470, w_054_477, w_054_479, w_054_482, w_054_492, w_054_499, w_054_508, w_054_509, w_054_518, w_054_532, w_054_535, w_054_537, w_054_540, w_054_544, w_054_546, w_054_549, w_054_553, w_054_570, w_054_572, w_054_577, w_054_578, w_054_579, w_054_581, w_054_592, w_054_596, w_054_599, w_054_606, w_054_618, w_054_620, w_054_628, w_054_629, w_054_630, w_054_631, w_054_632, w_054_633, w_054_634, w_054_635, w_054_636, w_054_637;
  wire w_055_001, w_055_005, w_055_007, w_055_012, w_055_021, w_055_023, w_055_036, w_055_044, w_055_053, w_055_057, w_055_061, w_055_076, w_055_087, w_055_090, w_055_094, w_055_100, w_055_104, w_055_109, w_055_111, w_055_113, w_055_123, w_055_128, w_055_148, w_055_149, w_055_154, w_055_155, w_055_157, w_055_160, w_055_162, w_055_164, w_055_167, w_055_169, w_055_170, w_055_173, w_055_181, w_055_213, w_055_214, w_055_216, w_055_220, w_055_226, w_055_232, w_055_233, w_055_242, w_055_243, w_055_245, w_055_253, w_055_254, w_055_259, w_055_260, w_055_261, w_055_284, w_055_291, w_055_292, w_055_300, w_055_306, w_055_311, w_055_324, w_055_325, w_055_327, w_055_335, w_055_339, w_055_361, w_055_363, w_055_370, w_055_373, w_055_382, w_055_385, w_055_389, w_055_420, w_055_421, w_055_422, w_055_423, w_055_435, w_055_443, w_055_466, w_055_469, w_055_473, w_055_475, w_055_494, w_055_525, w_055_526, w_055_567, w_055_576, w_055_590, w_055_594, w_055_598, w_055_602, w_055_604, w_055_610, w_055_636, w_055_647, w_055_650, w_055_660, w_055_661, w_055_671, w_055_672, w_055_693, w_055_715, w_055_716, w_055_717, w_055_735, w_055_744, w_055_750, w_055_772, w_055_775, w_055_786, w_055_821, w_055_828, w_055_835, w_055_852, w_055_856;
  wire w_056_000, w_056_018, w_056_020, w_056_023, w_056_033, w_056_085, w_056_086, w_056_112, w_056_114, w_056_124, w_056_125, w_056_161, w_056_164, w_056_165, w_056_178, w_056_182, w_056_192, w_056_193, w_056_196, w_056_203, w_056_211, w_056_217, w_056_231, w_056_233, w_056_246, w_056_251, w_056_254, w_056_273, w_056_298, w_056_315, w_056_333, w_056_382, w_056_411, w_056_441, w_056_492, w_056_503, w_056_504, w_056_512, w_056_519, w_056_589, w_056_615, w_056_625, w_056_637, w_056_650, w_056_658, w_056_659, w_056_668, w_056_679, w_056_717, w_056_727, w_056_745, w_056_751, w_056_795, w_056_800, w_056_810, w_056_821, w_056_830, w_056_833, w_056_835, w_056_876, w_056_890, w_056_894, w_056_928, w_056_929, w_056_936, w_056_972, w_056_980, w_056_1064, w_056_1109, w_056_1115, w_056_1121, w_056_1172, w_056_1176, w_056_1184, w_056_1223, w_056_1229, w_056_1269, w_056_1275, w_056_1290, w_056_1315, w_056_1342, w_056_1363, w_056_1388, w_056_1391, w_056_1409, w_056_1424, w_056_1446, w_056_1460, w_056_1465, w_056_1468, w_056_1502, w_056_1511, w_056_1534, w_056_1537, w_056_1540, w_056_1562, w_056_1615, w_056_1623, w_056_1651, w_056_1671;
  wire w_057_025, w_057_034, w_057_037, w_057_058, w_057_105, w_057_137, w_057_145, w_057_177, w_057_186, w_057_190, w_057_209, w_057_222, w_057_225, w_057_228, w_057_233, w_057_239, w_057_240, w_057_250, w_057_276, w_057_277, w_057_284, w_057_298, w_057_330, w_057_369, w_057_399, w_057_413, w_057_430, w_057_454, w_057_487, w_057_516, w_057_551, w_057_592, w_057_606, w_057_632, w_057_645, w_057_653, w_057_660, w_057_676, w_057_709, w_057_743, w_057_790, w_057_816, w_057_828, w_057_829, w_057_832, w_057_854, w_057_857, w_057_861, w_057_883, w_057_915, w_057_928, w_057_936, w_057_983, w_057_984, w_057_1003, w_057_1031, w_057_1038, w_057_1047, w_057_1060, w_057_1103, w_057_1124, w_057_1156, w_057_1158, w_057_1166, w_057_1174, w_057_1216, w_057_1249, w_057_1252, w_057_1266, w_057_1301, w_057_1307, w_057_1337, w_057_1351, w_057_1360, w_057_1410, w_057_1414, w_057_1445, w_057_1467, w_057_1517, w_057_1525, w_057_1536, w_057_1562, w_057_1591, w_057_1599, w_057_1600, w_057_1605, w_057_1615, w_057_1646, w_057_1717, w_057_1740, w_057_1768, w_057_1817, w_057_1838;
  wire w_058_011, w_058_025, w_058_034, w_058_038, w_058_041, w_058_054, w_058_058, w_058_064, w_058_074, w_058_080, w_058_097, w_058_108, w_058_125, w_058_147, w_058_174, w_058_186, w_058_190, w_058_196, w_058_199, w_058_203, w_058_212, w_058_220, w_058_240, w_058_242, w_058_266, w_058_302, w_058_315, w_058_360, w_058_367, w_058_392, w_058_403, w_058_415, w_058_431, w_058_436, w_058_459, w_058_481, w_058_498, w_058_521, w_058_531, w_058_533, w_058_553, w_058_589, w_058_608, w_058_616, w_058_625, w_058_649, w_058_701, w_058_732, w_058_743, w_058_762, w_058_768, w_058_780, w_058_794, w_058_809, w_058_814, w_058_822, w_058_828, w_058_840, w_058_843, w_058_875, w_058_885, w_058_891, w_058_919, w_058_935, w_058_938, w_058_955, w_058_961, w_058_1006, w_058_1019, w_058_1023, w_058_1027, w_058_1033, w_058_1040, w_058_1050, w_058_1064, w_058_1086, w_058_1121, w_058_1144, w_058_1145, w_058_1146, w_058_1160, w_058_1169, w_058_1187, w_058_1190, w_058_1220, w_058_1236, w_058_1255, w_058_1291, w_058_1294, w_058_1300, w_058_1346, w_058_1347, w_058_1412, w_058_1424, w_058_1469, w_058_1473, w_058_1478, w_058_1485, w_058_1500, w_058_1589, w_058_1606, w_058_1624, w_058_1629, w_058_1630, w_058_1712, w_058_1721, w_058_1743, w_058_1762, w_058_1779;
  wire w_059_008, w_059_014, w_059_017, w_059_020, w_059_023, w_059_042, w_059_052, w_059_059, w_059_065, w_059_080, w_059_082, w_059_084, w_059_093, w_059_096, w_059_113, w_059_117, w_059_125, w_059_127, w_059_139, w_059_152, w_059_158, w_059_165, w_059_172, w_059_175, w_059_179, w_059_183, w_059_184, w_059_206, w_059_207, w_059_210, w_059_214, w_059_228, w_059_229, w_059_246, w_059_272, w_059_278, w_059_284, w_059_288, w_059_289, w_059_293, w_059_296, w_059_298, w_059_303, w_059_318, w_059_333, w_059_344, w_059_346, w_059_353, w_059_360, w_059_361, w_059_381, w_059_383, w_059_395, w_059_403, w_059_429, w_059_435, w_059_445, w_059_450, w_059_457, w_059_463, w_059_478, w_059_482, w_059_485, w_059_489, w_059_492, w_059_497, w_059_503, w_059_509, w_059_518, w_059_549, w_059_561, w_059_565, w_059_572, w_059_573, w_059_577, w_059_597, w_059_599, w_059_606, w_059_608, w_059_619, w_059_622, w_059_632, w_059_651, w_059_653, w_059_692;
  wire w_060_003, w_060_005, w_060_006, w_060_007, w_060_009, w_060_010, w_060_011, w_060_012, w_060_013, w_060_016, w_060_018, w_060_019, w_060_020, w_060_022, w_060_024, w_060_025, w_060_026, w_060_028, w_060_029, w_060_030, w_060_031, w_060_032, w_060_033, w_060_034, w_060_035, w_060_037, w_060_038, w_060_039, w_060_040, w_060_041, w_060_046, w_060_047, w_060_052, w_060_053, w_060_054, w_060_055, w_060_056, w_060_057, w_060_058, w_060_059, w_060_060, w_060_062, w_060_063, w_060_065, w_060_066, w_060_067, w_060_069, w_060_070, w_060_072, w_060_074, w_060_076, w_060_077, w_060_080, w_060_081, w_060_082, w_060_084, w_060_088, w_060_091, w_060_093, w_060_094, w_060_095, w_060_096, w_060_097, w_060_098, w_060_100, w_060_101, w_060_102, w_060_103, w_060_104, w_060_106;
  wire w_061_000, w_061_009, w_061_012, w_061_049, w_061_055, w_061_071, w_061_076, w_061_084, w_061_089, w_061_106, w_061_108, w_061_114, w_061_121, w_061_151, w_061_161, w_061_182, w_061_184, w_061_201, w_061_212, w_061_213, w_061_216, w_061_217, w_061_223, w_061_232, w_061_236, w_061_240, w_061_255, w_061_260, w_061_263, w_061_274, w_061_279, w_061_280, w_061_293, w_061_297, w_061_300, w_061_303, w_061_322, w_061_337, w_061_363, w_061_367, w_061_373, w_061_374, w_061_375, w_061_392, w_061_400, w_061_404, w_061_409, w_061_411, w_061_424, w_061_426, w_061_430, w_061_435, w_061_437, w_061_450, w_061_461, w_061_468, w_061_473, w_061_479, w_061_486, w_061_497, w_061_506, w_061_513, w_061_517, w_061_535, w_061_538, w_061_540, w_061_546, w_061_548, w_061_552, w_061_560, w_061_568, w_061_582, w_061_585, w_061_607, w_061_622, w_061_633, w_061_643, w_061_644, w_061_663;
  wire w_062_015, w_062_027, w_062_032, w_062_033, w_062_063, w_062_064, w_062_071, w_062_072, w_062_077, w_062_094, w_062_097, w_062_105, w_062_106, w_062_127, w_062_137, w_062_140, w_062_186, w_062_196, w_062_211, w_062_240, w_062_243, w_062_271, w_062_286, w_062_337, w_062_341, w_062_349, w_062_362, w_062_393, w_062_408, w_062_418, w_062_433, w_062_436, w_062_447, w_062_465, w_062_497, w_062_504, w_062_527, w_062_544, w_062_556, w_062_571, w_062_587, w_062_605, w_062_608, w_062_618, w_062_689, w_062_720, w_062_732, w_062_782, w_062_783, w_062_787, w_062_805, w_062_817, w_062_876, w_062_878, w_062_887, w_062_900, w_062_962, w_062_972, w_062_973, w_062_998, w_062_1003, w_062_1016, w_062_1111, w_062_1124, w_062_1158, w_062_1177, w_062_1180, w_062_1181, w_062_1222, w_062_1289, w_062_1292, w_062_1296, w_062_1307, w_062_1332;
  wire w_063_006, w_063_016, w_063_019, w_063_027, w_063_038, w_063_041, w_063_043, w_063_049, w_063_054, w_063_055, w_063_059, w_063_060, w_063_093, w_063_095, w_063_129, w_063_137, w_063_140, w_063_145, w_063_171, w_063_175, w_063_183, w_063_184, w_063_194, w_063_255, w_063_264, w_063_270, w_063_283, w_063_287, w_063_289, w_063_292, w_063_295, w_063_312, w_063_345, w_063_358, w_063_373, w_063_375, w_063_388, w_063_392, w_063_407, w_063_422, w_063_566, w_063_572, w_063_590, w_063_597, w_063_600, w_063_613, w_063_618, w_063_619, w_063_629, w_063_695, w_063_706, w_063_722, w_063_725, w_063_749, w_063_837, w_063_909, w_063_966, w_063_975, w_063_1029, w_063_1040, w_063_1059, w_063_1088, w_063_1094, w_063_1100, w_063_1122, w_063_1140, w_063_1149, w_063_1157, w_063_1164, w_063_1171, w_063_1173, w_063_1247, w_063_1251, w_063_1265, w_063_1294, w_063_1297, w_063_1311, w_063_1336, w_063_1337, w_063_1375, w_063_1411, w_063_1422, w_063_1429, w_063_1486, w_063_1492, w_063_1500, w_063_1501, w_063_1561, w_063_1578, w_063_1583, w_063_1594, w_063_1604;
  wire w_064_036, w_064_039, w_064_085, w_064_096, w_064_102, w_064_108, w_064_115, w_064_140, w_064_141, w_064_145, w_064_147, w_064_156, w_064_159, w_064_170, w_064_179, w_064_190, w_064_193, w_064_197, w_064_210, w_064_227, w_064_234, w_064_239, w_064_252, w_064_254, w_064_264, w_064_266, w_064_293, w_064_305, w_064_330, w_064_364, w_064_380, w_064_396, w_064_405, w_064_455, w_064_474, w_064_479, w_064_492, w_064_563, w_064_586, w_064_607, w_064_609, w_064_631, w_064_636, w_064_639, w_064_666, w_064_677, w_064_728, w_064_749, w_064_772, w_064_775, w_064_790, w_064_795, w_064_805, w_064_829, w_064_861, w_064_884, w_064_889, w_064_891, w_064_904, w_064_912, w_064_926, w_064_941, w_064_954, w_064_996, w_064_999, w_064_1012, w_064_1046, w_064_1047, w_064_1058, w_064_1064, w_064_1081, w_064_1094, w_064_1135, w_064_1137, w_064_1140, w_064_1150, w_064_1154, w_064_1161, w_064_1186, w_064_1204, w_064_1225, w_064_1238, w_064_1283, w_064_1303, w_064_1323, w_064_1337, w_064_1362, w_064_1374, w_064_1377, w_064_1392, w_064_1433, w_064_1435, w_064_1438, w_064_1440, w_064_1456, w_064_1466, w_064_1474, w_064_1509, w_064_1513, w_064_1583, w_064_1594, w_064_1602, w_064_1643, w_064_1658;
  wire w_065_000, w_065_001, w_065_002, w_065_003, w_065_004, w_065_005;
  wire w_066_007, w_066_009, w_066_013, w_066_016, w_066_022, w_066_043, w_066_047, w_066_063, w_066_066, w_066_069, w_066_075, w_066_077, w_066_086, w_066_090, w_066_116, w_066_142, w_066_154, w_066_156, w_066_162, w_066_188, w_066_213, w_066_222, w_066_223, w_066_282, w_066_291, w_066_307, w_066_324, w_066_327, w_066_332, w_066_355, w_066_363, w_066_373, w_066_378, w_066_380, w_066_404, w_066_412, w_066_430, w_066_522, w_066_537, w_066_546, w_066_558, w_066_562, w_066_574, w_066_602, w_066_640, w_066_702, w_066_714, w_066_722, w_066_731, w_066_738, w_066_753, w_066_767, w_066_798, w_066_823, w_066_845, w_066_859, w_066_863, w_066_870, w_066_889, w_066_896, w_066_898, w_066_900, w_066_909, w_066_930, w_066_971, w_066_989, w_066_1009, w_066_1027, w_066_1040, w_066_1093, w_066_1151;
  wire w_067_017, w_067_019, w_067_048, w_067_080, w_067_105, w_067_160, w_067_179, w_067_183, w_067_185, w_067_200, w_067_206, w_067_209, w_067_225, w_067_237, w_067_258, w_067_267, w_067_280, w_067_287, w_067_288, w_067_292, w_067_338, w_067_360, w_067_376, w_067_403, w_067_418, w_067_434, w_067_462, w_067_477, w_067_512, w_067_531, w_067_532, w_067_541, w_067_544, w_067_558, w_067_582, w_067_589, w_067_595, w_067_603, w_067_609, w_067_620, w_067_639, w_067_651, w_067_655, w_067_665, w_067_676, w_067_682, w_067_688, w_067_690, w_067_692, w_067_696, w_067_703, w_067_727, w_067_742, w_067_746, w_067_758, w_067_763, w_067_786, w_067_799, w_067_807, w_067_871, w_067_872, w_067_896, w_067_898, w_067_905, w_067_912, w_067_943, w_067_961, w_067_962, w_067_965;
  wire w_068_000, w_068_003, w_068_011, w_068_013, w_068_017, w_068_018, w_068_019, w_068_021, w_068_022, w_068_026, w_068_027, w_068_029, w_068_030, w_068_031, w_068_036, w_068_037, w_068_038, w_068_041, w_068_048, w_068_050, w_068_055, w_068_059, w_068_062, w_068_073, w_068_075, w_068_078, w_068_083, w_068_085, w_068_086, w_068_095, w_068_097, w_068_105, w_068_106, w_068_110, w_068_114, w_068_119, w_068_126, w_068_135, w_068_140, w_068_141, w_068_142, w_068_151, w_068_157, w_068_160, w_068_163, w_068_164, w_068_165, w_068_166, w_068_169, w_068_171, w_068_176, w_068_179, w_068_184, w_068_189, w_068_190, w_068_194, w_068_197, w_068_200, w_068_203, w_068_209, w_068_210, w_068_211, w_068_216, w_068_223, w_068_224, w_068_233, w_068_234, w_068_236, w_068_239, w_068_240, w_068_243;
  wire w_069_001, w_069_019, w_069_021, w_069_038, w_069_039, w_069_049, w_069_053, w_069_068, w_069_072, w_069_182, w_069_188, w_069_283, w_069_312, w_069_331, w_069_350, w_069_368, w_069_436, w_069_474, w_069_479, w_069_510, w_069_568, w_069_620, w_069_681, w_069_723, w_069_760, w_069_805, w_069_828, w_069_866, w_069_920, w_069_921, w_069_970, w_069_976, w_069_980, w_069_1167, w_069_1270, w_069_1276, w_069_1285, w_069_1356, w_069_1365, w_069_1369, w_069_1571, w_069_1600, w_069_1618, w_069_1620, w_069_1642, w_069_1675, w_069_1681, w_069_1723, w_069_1729, w_069_1731, w_069_1744, w_069_1762, w_069_1776, w_069_1807, w_069_1818;
  wire w_070_004, w_070_005, w_070_013, w_070_014, w_070_015, w_070_022, w_070_031, w_070_032, w_070_034, w_070_035, w_070_045, w_070_050, w_070_051, w_070_056, w_070_061, w_070_062, w_070_077, w_070_079, w_070_080, w_070_093, w_070_107, w_070_110, w_070_114, w_070_120, w_070_146, w_070_149, w_070_150, w_070_160, w_070_172, w_070_175, w_070_177, w_070_180, w_070_182, w_070_183, w_070_204, w_070_212, w_070_213, w_070_231, w_070_244, w_070_250, w_070_260, w_070_270, w_070_285, w_070_314, w_070_318, w_070_369, w_070_371, w_070_374, w_070_376, w_070_379, w_070_387, w_070_391, w_070_401, w_070_405, w_070_409, w_070_423, w_070_427, w_070_430, w_070_432, w_070_446, w_070_448, w_070_450, w_070_455, w_070_459, w_070_463, w_070_471, w_070_472;
  wire w_071_007, w_071_011, w_071_012, w_071_016, w_071_018, w_071_025, w_071_028, w_071_033, w_071_040, w_071_043, w_071_044, w_071_048, w_071_052, w_071_056, w_071_061, w_071_064, w_071_066, w_071_070, w_071_071, w_071_082, w_071_086, w_071_108, w_071_125, w_071_130, w_071_151, w_071_164, w_071_167, w_071_191, w_071_193, w_071_202, w_071_224, w_071_227, w_071_235, w_071_263, w_071_274, w_071_289, w_071_293, w_071_295, w_071_303, w_071_306, w_071_312, w_071_323, w_071_339, w_071_341, w_071_355, w_071_357, w_071_358, w_071_361, w_071_380, w_071_385, w_071_406, w_071_437, w_071_442, w_071_457, w_071_465, w_071_477, w_071_481, w_071_488, w_071_519, w_071_522, w_071_523, w_071_529, w_071_531, w_071_550;
  wire w_072_001, w_072_002, w_072_003, w_072_005, w_072_006, w_072_007, w_072_008, w_072_010, w_072_013, w_072_019, w_072_022, w_072_024, w_072_032, w_072_035, w_072_038, w_072_040, w_072_042, w_072_047, w_072_048, w_072_049, w_072_051, w_072_052, w_072_053, w_072_054, w_072_055, w_072_058, w_072_059, w_072_066, w_072_067, w_072_068, w_072_069, w_072_070, w_072_073, w_072_074, w_072_075, w_072_076, w_072_077, w_072_079, w_072_081;
  wire w_073_003, w_073_004, w_073_005, w_073_006, w_073_008, w_073_009, w_073_010, w_073_011, w_073_012, w_073_016, w_073_018, w_073_019, w_073_021, w_073_022, w_073_023, w_073_029, w_073_030, w_073_031, w_073_034, w_073_036, w_073_037, w_073_042, w_073_043, w_073_053, w_073_059, w_073_061, w_073_062, w_073_063, w_073_064, w_073_065, w_073_066, w_073_067, w_073_069, w_073_071, w_073_072, w_073_073, w_073_076, w_073_079, w_073_082, w_073_083, w_073_087, w_073_090, w_073_091, w_073_093, w_073_094, w_073_096, w_073_099, w_073_100, w_073_101;
  wire w_074_026, w_074_039, w_074_054, w_074_059, w_074_080, w_074_115, w_074_128, w_074_129, w_074_136, w_074_155, w_074_167, w_074_169, w_074_212, w_074_214, w_074_215, w_074_219, w_074_231, w_074_241, w_074_246, w_074_262, w_074_273, w_074_274, w_074_278, w_074_295, w_074_298, w_074_357, w_074_422, w_074_496, w_074_501, w_074_551, w_074_557, w_074_558, w_074_582, w_074_583, w_074_584, w_074_625, w_074_658, w_074_680, w_074_690, w_074_713, w_074_811, w_074_869, w_074_954, w_074_961, w_074_1006, w_074_1023, w_074_1032, w_074_1077, w_074_1109, w_074_1217, w_074_1229, w_074_1230, w_074_1250, w_074_1265, w_074_1283, w_074_1310, w_074_1335, w_074_1365, w_074_1427, w_074_1449, w_074_1450, w_074_1467, w_074_1470, w_074_1501, w_074_1578, w_074_1647, w_074_1683, w_074_1697;
  wire w_075_000, w_075_001, w_075_003, w_075_005, w_075_014, w_075_025, w_075_037, w_075_049, w_075_051, w_075_054, w_075_055, w_075_059, w_075_061, w_075_062, w_075_065, w_075_071, w_075_074, w_075_082, w_075_087, w_075_091, w_075_096, w_075_097, w_075_098, w_075_105, w_075_109, w_075_116, w_075_117, w_075_118, w_075_127, w_075_132, w_075_144, w_075_151, w_075_152, w_075_159, w_075_167, w_075_172, w_075_173, w_075_174, w_075_179, w_075_184, w_075_187, w_075_213, w_075_214, w_075_217, w_075_221, w_075_231, w_075_234, w_075_237, w_075_238, w_075_239, w_075_241, w_075_247, w_075_249, w_075_252, w_075_254, w_075_257, w_075_261, w_075_263, w_075_264, w_075_266, w_075_282;
  wire w_076_006, w_076_010, w_076_025, w_076_034, w_076_039, w_076_045, w_076_046, w_076_048, w_076_049, w_076_057, w_076_058, w_076_066, w_076_074, w_076_076, w_076_078, w_076_085, w_076_094, w_076_103, w_076_118, w_076_119, w_076_120, w_076_128, w_076_138, w_076_140, w_076_146, w_076_149, w_076_155, w_076_169, w_076_180, w_076_200, w_076_203, w_076_208, w_076_209, w_076_210, w_076_211, w_076_215, w_076_240, w_076_242, w_076_244, w_076_262, w_076_267, w_076_285, w_076_288, w_076_290, w_076_296, w_076_311, w_076_327, w_076_330, w_076_333, w_076_335, w_076_338, w_076_344, w_076_354, w_076_355, w_076_356;
  wire w_077_009, w_077_014, w_077_023, w_077_034, w_077_055, w_077_134, w_077_151, w_077_153, w_077_170, w_077_174, w_077_197, w_077_201, w_077_209, w_077_223, w_077_232, w_077_238, w_077_252, w_077_310, w_077_314, w_077_438, w_077_439, w_077_460, w_077_490, w_077_494, w_077_526, w_077_540, w_077_568, w_077_571, w_077_589, w_077_596, w_077_602, w_077_623, w_077_632, w_077_642, w_077_658, w_077_664, w_077_701, w_077_702, w_077_709, w_077_725, w_077_769, w_077_798, w_077_873, w_077_895, w_077_903, w_077_914, w_077_927, w_077_945, w_077_997, w_077_1006, w_077_1084, w_077_1107, w_077_1114, w_077_1148;
  wire w_078_019, w_078_037, w_078_048, w_078_053, w_078_055, w_078_088, w_078_089, w_078_092, w_078_093, w_078_103, w_078_109, w_078_113, w_078_148, w_078_195, w_078_205, w_078_217, w_078_218, w_078_236, w_078_252, w_078_261, w_078_281, w_078_285, w_078_287, w_078_289, w_078_347, w_078_349, w_078_353, w_078_434, w_078_455, w_078_479, w_078_500, w_078_538, w_078_557, w_078_632, w_078_636, w_078_723, w_078_747, w_078_778, w_078_801, w_078_829, w_078_835, w_078_854, w_078_863, w_078_864, w_078_865, w_078_872, w_078_884, w_078_937, w_078_969, w_078_995, w_078_1036, w_078_1042, w_078_1120, w_078_1150, w_078_1153, w_078_1155, w_078_1184, w_078_1276, w_078_1286, w_078_1342, w_078_1347, w_078_1349, w_078_1352, w_078_1362, w_078_1469, w_078_1496, w_078_1506, w_078_1631, w_078_1664, w_078_1688;
  wire w_079_005, w_079_015, w_079_018, w_079_020, w_079_030, w_079_034, w_079_048, w_079_078, w_079_094, w_079_104, w_079_112, w_079_115, w_079_126, w_079_128, w_079_134, w_079_142, w_079_145, w_079_159, w_079_162, w_079_176, w_079_202, w_079_216, w_079_218, w_079_233, w_079_261, w_079_270, w_079_293, w_079_321, w_079_363, w_079_374, w_079_382, w_079_395, w_079_411, w_079_425, w_079_463, w_079_502, w_079_526, w_079_536, w_079_539, w_079_556, w_079_564, w_079_568, w_079_573, w_079_577, w_079_578, w_079_588, w_079_598, w_079_612, w_079_622, w_079_640, w_079_649, w_079_651, w_079_667, w_079_718, w_079_721, w_079_747, w_079_748, w_079_753, w_079_784, w_079_789, w_079_797, w_079_819, w_079_839, w_079_847, w_079_848;
  wire w_080_000, w_080_001, w_080_007, w_080_008, w_080_010, w_080_013, w_080_018, w_080_019, w_080_021, w_080_024, w_080_028, w_080_030, w_080_034, w_080_036, w_080_040, w_080_048, w_080_049, w_080_050, w_080_051, w_080_059, w_080_061, w_080_067, w_080_068, w_080_069, w_080_070, w_080_077, w_080_082, w_080_090, w_080_095, w_080_096, w_080_099, w_080_102, w_080_103, w_080_105, w_080_106, w_080_109, w_080_110, w_080_111, w_080_112, w_080_114, w_080_115, w_080_118, w_080_119;
  wire w_081_028, w_081_040, w_081_050, w_081_055, w_081_059, w_081_077, w_081_086, w_081_093, w_081_095, w_081_107, w_081_142, w_081_162, w_081_183, w_081_208, w_081_221, w_081_223, w_081_242, w_081_249, w_081_290, w_081_311, w_081_341, w_081_354, w_081_377, w_081_385, w_081_392, w_081_407, w_081_415, w_081_416, w_081_430, w_081_437, w_081_447, w_081_468, w_081_480, w_081_481, w_081_490, w_081_532, w_081_539, w_081_558, w_081_560, w_081_571, w_081_572, w_081_576, w_081_578, w_081_582, w_081_619, w_081_647, w_081_663, w_081_665, w_081_669, w_081_678;
  wire w_082_083, w_082_092, w_082_095, w_082_099, w_082_115, w_082_120, w_082_155, w_082_179, w_082_193, w_082_233, w_082_240, w_082_260, w_082_262, w_082_265, w_082_275, w_082_303, w_082_314, w_082_337, w_082_341, w_082_358, w_082_382, w_082_409, w_082_414, w_082_422, w_082_423, w_082_426, w_082_431, w_082_466, w_082_500, w_082_507, w_082_510, w_082_515, w_082_517, w_082_527, w_082_529, w_082_549, w_082_586, w_082_589, w_082_593, w_082_597, w_082_649, w_082_658, w_082_688, w_082_691, w_082_698, w_082_721, w_082_734, w_082_745, w_082_782, w_082_799, w_082_808, w_082_813;
  wire w_083_000, w_083_001, w_083_002, w_083_003, w_083_004, w_083_005, w_083_006, w_083_007, w_083_008, w_083_010, w_083_011, w_083_013, w_083_014, w_083_015, w_083_016, w_083_017, w_083_019, w_083_020, w_083_021, w_083_022, w_083_023, w_083_024, w_083_025, w_083_026, w_083_028, w_083_029, w_083_030, w_083_031;
  wire w_084_012, w_084_013, w_084_016, w_084_019, w_084_036, w_084_041, w_084_050, w_084_055, w_084_058, w_084_065, w_084_070, w_084_071, w_084_073, w_084_079, w_084_080, w_084_091, w_084_123, w_084_139, w_084_142, w_084_144, w_084_158, w_084_164, w_084_168, w_084_197, w_084_207, w_084_211, w_084_233, w_084_260, w_084_267, w_084_270, w_084_271, w_084_275, w_084_304, w_084_314, w_084_315, w_084_317, w_084_333, w_084_334, w_084_343, w_084_351, w_084_362, w_084_364, w_084_366, w_084_367, w_084_375, w_084_379, w_084_385, w_084_391, w_084_405, w_084_410, w_084_418, w_084_458, w_084_470, w_084_474, w_084_481, w_084_483;
  wire w_085_001, w_085_030, w_085_033, w_085_046, w_085_058, w_085_059, w_085_064, w_085_071, w_085_081, w_085_098, w_085_099, w_085_108, w_085_109, w_085_111, w_085_115, w_085_122, w_085_127, w_085_134, w_085_135, w_085_146, w_085_153, w_085_177, w_085_181, w_085_184, w_085_200, w_085_201, w_085_204, w_085_221, w_085_254, w_085_256, w_085_270, w_085_274, w_085_302, w_085_314, w_085_355, w_085_357, w_085_363, w_085_373, w_085_385, w_085_388, w_085_395, w_085_418, w_085_427, w_085_439, w_085_454, w_085_486, w_085_490, w_085_496, w_085_505, w_085_511, w_085_513, w_085_522, w_085_536, w_085_568, w_085_571, w_085_576, w_085_593, w_085_602, w_085_607, w_085_609, w_085_653, w_085_660, w_085_676;
  wire w_086_025, w_086_044, w_086_049, w_086_055, w_086_066, w_086_095, w_086_096, w_086_108, w_086_119, w_086_160, w_086_166, w_086_176, w_086_178, w_086_203, w_086_235, w_086_267, w_086_288, w_086_291, w_086_301, w_086_326, w_086_342, w_086_370, w_086_371, w_086_402, w_086_515, w_086_539, w_086_555, w_086_569, w_086_633, w_086_652, w_086_677, w_086_742, w_086_748, w_086_755, w_086_780, w_086_812, w_086_838, w_086_896, w_086_909, w_086_923, w_086_991, w_086_1093, w_086_1118, w_086_1168, w_086_1257, w_086_1269, w_086_1316, w_086_1430, w_086_1493, w_086_1567, w_086_1569, w_086_1575, w_086_1642;
  wire w_087_021, w_087_063, w_087_110, w_087_115, w_087_146, w_087_206, w_087_242, w_087_289, w_087_304, w_087_347, w_087_393, w_087_462, w_087_467, w_087_524, w_087_566, w_087_590, w_087_607, w_087_662, w_087_709, w_087_772, w_087_840, w_087_874, w_087_971, w_087_973, w_087_978, w_087_984, w_087_1001, w_087_1009, w_087_1021, w_087_1050, w_087_1062, w_087_1068, w_087_1097, w_087_1098, w_087_1104, w_087_1123, w_087_1173, w_087_1211, w_087_1279, w_087_1302, w_087_1307, w_087_1314, w_087_1366, w_087_1383, w_087_1426, w_087_1451, w_087_1494, w_087_1547, w_087_1581, w_087_1584, w_087_1603, w_087_1609, w_087_1682;
  wire w_088_020, w_088_030, w_088_059, w_088_067, w_088_114, w_088_118, w_088_125, w_088_139, w_088_189, w_088_210, w_088_213, w_088_239, w_088_258, w_088_279, w_088_286, w_088_291, w_088_293, w_088_326, w_088_366, w_088_421, w_088_429, w_088_437, w_088_447, w_088_455, w_088_458, w_088_467, w_088_482, w_088_507, w_088_520, w_088_528, w_088_552, w_088_594, w_088_597, w_088_629, w_088_642, w_088_651, w_088_663, w_088_698, w_088_699, w_088_729, w_088_768, w_088_815, w_088_900, w_088_931, w_088_948, w_088_1020, w_088_1028, w_088_1150, w_088_1152, w_088_1154, w_088_1192, w_088_1214, w_088_1239, w_088_1307, w_088_1340, w_088_1369;
  wire w_089_019, w_089_060, w_089_066, w_089_067, w_089_080, w_089_081, w_089_101, w_089_107, w_089_114, w_089_127, w_089_150, w_089_155, w_089_156, w_089_179, w_089_191, w_089_222, w_089_282, w_089_309, w_089_328, w_089_329, w_089_340, w_089_360, w_089_363, w_089_373, w_089_377, w_089_390, w_089_402, w_089_408, w_089_419, w_089_427, w_089_438, w_089_449, w_089_524, w_089_547, w_089_578, w_089_604, w_089_627, w_089_629, w_089_635, w_089_647, w_089_649, w_089_679, w_089_688, w_089_689, w_089_693, w_089_721, w_089_727, w_089_808, w_089_815, w_089_832, w_089_873, w_089_874, w_089_948, w_089_951, w_089_962, w_089_1077, w_089_1140, w_089_1149, w_089_1169, w_089_1204, w_089_1209, w_089_1226, w_089_1242, w_089_1252, w_089_1258, w_089_1266, w_089_1277, w_089_1290, w_089_1302;
  wire w_090_015, w_090_085, w_090_095, w_090_145, w_090_146, w_090_172, w_090_195, w_090_196, w_090_201, w_090_210, w_090_223, w_090_226, w_090_244, w_090_250, w_090_266, w_090_314, w_090_341, w_090_363, w_090_384, w_090_392, w_090_393, w_090_413, w_090_414, w_090_427, w_090_457, w_090_467, w_090_474, w_090_510, w_090_553, w_090_606, w_090_615, w_090_648, w_090_663, w_090_672, w_090_696, w_090_709, w_090_716, w_090_747, w_090_813, w_090_874, w_090_875, w_090_906, w_090_919, w_090_940, w_090_984, w_090_1067, w_090_1125, w_090_1139, w_090_1154, w_090_1208;
  wire w_091_003, w_091_004, w_091_006, w_091_008, w_091_012, w_091_021, w_091_022, w_091_024, w_091_025, w_091_030, w_091_033, w_091_039, w_091_049, w_091_052, w_091_054, w_091_056, w_091_059, w_091_065, w_091_069, w_091_077, w_091_081, w_091_088, w_091_089, w_091_090, w_091_097, w_091_099, w_091_100, w_091_101, w_091_105, w_091_106, w_091_107, w_091_112, w_091_113, w_091_119, w_091_122, w_091_124, w_091_125, w_091_128, w_091_130, w_091_132, w_091_133, w_091_140, w_091_141, w_091_145, w_091_150, w_091_159, w_091_162, w_091_163, w_091_176, w_091_177, w_091_180, w_091_182;
  wire w_092_004, w_092_026, w_092_091, w_092_104, w_092_107, w_092_126, w_092_129, w_092_136, w_092_143, w_092_151, w_092_158, w_092_163, w_092_164, w_092_200, w_092_201, w_092_204, w_092_230, w_092_240, w_092_281, w_092_293, w_092_311, w_092_335, w_092_337, w_092_367, w_092_396, w_092_426, w_092_428, w_092_517, w_092_523, w_092_526, w_092_527, w_092_540, w_092_584, w_092_591, w_092_616, w_092_639, w_092_648, w_092_651, w_092_767, w_092_850, w_092_881, w_092_886, w_092_912, w_092_926, w_092_943, w_092_970, w_092_1039, w_092_1156, w_092_1159, w_092_1194;
  wire w_093_001, w_093_004, w_093_005, w_093_009, w_093_010, w_093_011, w_093_012, w_093_015, w_093_016, w_093_017, w_093_020, w_093_022, w_093_023, w_093_025, w_093_034, w_093_040, w_093_045, w_093_048, w_093_049, w_093_052, w_093_054, w_093_055, w_093_059, w_093_062, w_093_063, w_093_065, w_093_066, w_093_068, w_093_070;
  wire w_094_002, w_094_005, w_094_006, w_094_007, w_094_008, w_094_009, w_094_011, w_094_012, w_094_013, w_094_014, w_094_016, w_094_022, w_094_024, w_094_036, w_094_044, w_094_045, w_094_046, w_094_049, w_094_050, w_094_051, w_094_053, w_094_055, w_094_056, w_094_058, w_094_061, w_094_063, w_094_068, w_094_074, w_094_076, w_094_081, w_094_083, w_094_085, w_094_087, w_094_090, w_094_091, w_094_095, w_094_096, w_094_098, w_094_100;
  wire w_095_020, w_095_042, w_095_045, w_095_054, w_095_059, w_095_067, w_095_068, w_095_099, w_095_117, w_095_130, w_095_148, w_095_157, w_095_167, w_095_180, w_095_198, w_095_233, w_095_279, w_095_329, w_095_353, w_095_373, w_095_387, w_095_445, w_095_468, w_095_476, w_095_479, w_095_486, w_095_503, w_095_506, w_095_528, w_095_576, w_095_580, w_095_581, w_095_639, w_095_660, w_095_675, w_095_718, w_095_734, w_095_736, w_095_755, w_095_834, w_095_836, w_095_841, w_095_845, w_095_859, w_095_884, w_095_898, w_095_900;
  wire w_096_002, w_096_003, w_096_007, w_096_012, w_096_027, w_096_039, w_096_042, w_096_048, w_096_054, w_096_058, w_096_073, w_096_076, w_096_085, w_096_099, w_096_108, w_096_109, w_096_110, w_096_117, w_096_118, w_096_134, w_096_142, w_096_143, w_096_144, w_096_147, w_096_161, w_096_162, w_096_173, w_096_176, w_096_183, w_096_195, w_096_196, w_096_201, w_096_208, w_096_218, w_096_224, w_096_225, w_096_227, w_096_228;
  wire w_097_020, w_097_119, w_097_143, w_097_239, w_097_257, w_097_266, w_097_278, w_097_279, w_097_310, w_097_354, w_097_370, w_097_386, w_097_390, w_097_439, w_097_446, w_097_456, w_097_469, w_097_473, w_097_489, w_097_555, w_097_556, w_097_562, w_097_573, w_097_579, w_097_685, w_097_704, w_097_712, w_097_717, w_097_718, w_097_740, w_097_743, w_097_753, w_097_761, w_097_801, w_097_810, w_097_817, w_097_882, w_097_887;
  wire w_098_001, w_098_004, w_098_010, w_098_031, w_098_146, w_098_197, w_098_254, w_098_263, w_098_274, w_098_276, w_098_307, w_098_333, w_098_368, w_098_370, w_098_387, w_098_389, w_098_426, w_098_432, w_098_460, w_098_494, w_098_498, w_098_509, w_098_513, w_098_602, w_098_607, w_098_609, w_098_613, w_098_685, w_098_698, w_098_734, w_098_740, w_098_798, w_098_801, w_098_803, w_098_804, w_098_815, w_098_836, w_098_930, w_098_977, w_098_1010, w_098_1051, w_098_1076;
  wire w_099_036, w_099_037, w_099_039, w_099_048, w_099_080, w_099_096, w_099_136, w_099_139, w_099_140, w_099_149, w_099_161, w_099_172, w_099_191, w_099_211, w_099_214, w_099_224, w_099_282, w_099_292, w_099_389, w_099_412, w_099_429, w_099_453, w_099_495, w_099_519, w_099_545, w_099_553, w_099_611, w_099_632, w_099_677, w_099_686, w_099_691, w_099_714, w_099_796, w_099_816, w_099_818, w_099_837, w_099_937, w_099_994, w_099_1076, w_099_1080, w_099_1093;
  wire w_100_000, w_100_021, w_100_082, w_100_147, w_100_155, w_100_186, w_100_214, w_100_278, w_100_298, w_100_323, w_100_347, w_100_401, w_100_467, w_100_472, w_100_494, w_100_516, w_100_538, w_100_550, w_100_576, w_100_579, w_100_597, w_100_602, w_100_610, w_100_627, w_100_667, w_100_688, w_100_712, w_100_770, w_100_777, w_100_900, w_100_1069, w_100_1090, w_100_1155, w_100_1177, w_100_1197, w_100_1259, w_100_1316, w_100_1332, w_100_1363, w_100_1408, w_100_1442, w_100_1550, w_100_1567, w_100_1601, w_100_1813;
  wire w_101_033, w_101_079, w_101_094, w_101_120, w_101_142, w_101_145, w_101_154, w_101_166, w_101_203, w_101_221, w_101_227, w_101_244, w_101_324, w_101_354, w_101_356, w_101_367, w_101_368, w_101_432, w_101_437, w_101_453, w_101_496, w_101_523, w_101_539, w_101_566, w_101_594, w_101_615, w_101_655, w_101_661, w_101_670, w_101_672, w_101_684, w_101_745;
  wire w_102_010, w_102_017, w_102_030, w_102_072, w_102_126, w_102_130, w_102_211, w_102_294, w_102_346, w_102_363, w_102_370, w_102_462, w_102_505, w_102_507, w_102_519, w_102_520, w_102_594, w_102_605, w_102_763, w_102_797, w_102_848, w_102_931, w_102_948, w_102_1039, w_102_1199, w_102_1214, w_102_1216, w_102_1259, w_102_1260, w_102_1261, w_102_1262, w_102_1263, w_102_1264, w_102_1268, w_102_1269, w_102_1270, w_102_1271, w_102_1272, w_102_1273, w_102_1274, w_102_1275, w_102_1276, w_102_1278;
  wire w_103_031, w_103_062, w_103_064, w_103_088, w_103_098, w_103_113, w_103_133, w_103_146, w_103_169, w_103_196, w_103_232, w_103_233, w_103_237, w_103_252, w_103_286, w_103_294, w_103_304, w_103_321, w_103_329, w_103_369, w_103_375, w_103_378, w_103_445, w_103_462, w_103_523, w_103_538, w_103_553, w_103_554, w_103_561, w_103_590, w_103_629, w_103_647, w_103_663, w_103_692, w_103_718, w_103_833, w_103_977, w_103_994, w_103_1055, w_103_1200, w_103_1257, w_103_1264, w_103_1299, w_103_1313, w_103_1337, w_103_1375, w_103_1398, w_103_1422;
  wire w_104_128, w_104_176, w_104_202, w_104_233, w_104_385, w_104_430, w_104_529, w_104_613, w_104_634, w_104_635, w_104_663, w_104_684, w_104_695, w_104_723, w_104_759, w_104_773, w_104_776, w_104_784, w_104_800, w_104_813, w_104_938, w_104_1006, w_104_1022, w_104_1031, w_104_1049, w_104_1173, w_104_1248, w_104_1263, w_104_1410, w_104_1424, w_104_1546, w_104_1580, w_104_1581, w_104_1647, w_104_1651, w_104_1694, w_104_1704, w_104_1763, w_104_1768;
  wire w_105_000, w_105_012, w_105_043, w_105_048, w_105_063, w_105_074, w_105_090, w_105_117, w_105_123, w_105_126, w_105_146, w_105_297, w_105_330, w_105_442, w_105_458, w_105_476, w_105_507, w_105_552, w_105_635, w_105_636, w_105_671, w_105_740, w_105_819, w_105_872, w_105_875, w_105_956, w_105_957, w_105_1029, w_105_1042, w_105_1050, w_105_1105, w_105_1136, w_105_1171, w_105_1183, w_105_1248, w_105_1249, w_105_1352, w_105_1403, w_105_1459, w_105_1472, w_105_1578, w_105_1716, w_105_1809, w_105_1812;
  wire w_106_037, w_106_043, w_106_078, w_106_089, w_106_090, w_106_096, w_106_148, w_106_158, w_106_172, w_106_185, w_106_215, w_106_231, w_106_252, w_106_276, w_106_278, w_106_334, w_106_336, w_106_347, w_106_355, w_106_356, w_106_363, w_106_370, w_106_380, w_106_424, w_106_471, w_106_479, w_106_520, w_106_524, w_106_533, w_106_585, w_106_677, w_106_716, w_106_720, w_106_722, w_106_753, w_106_764, w_106_848, w_106_854, w_106_902, w_106_1034, w_106_1069, w_106_1199, w_106_1235, w_106_1249, w_106_1269, w_106_1377;
  wire w_107_000, w_107_007, w_107_055, w_107_188, w_107_211, w_107_272, w_107_282, w_107_286, w_107_296, w_107_308, w_107_332, w_107_364, w_107_398, w_107_430, w_107_432, w_107_440, w_107_468, w_107_488, w_107_495, w_107_544, w_107_571, w_107_576, w_107_581, w_107_651, w_107_660, w_107_684, w_107_731, w_107_821, w_107_888, w_107_971, w_107_995, w_107_1115, w_107_1194, w_107_1322;
  wire w_108_007, w_108_008, w_108_009, w_108_019, w_108_022, w_108_054, w_108_055, w_108_067, w_108_076, w_108_128, w_108_134, w_108_149, w_108_207, w_108_225, w_108_245, w_108_251, w_108_261, w_108_266, w_108_277, w_108_286, w_108_309, w_108_374, w_108_381, w_108_387, w_108_398, w_108_428, w_108_467, w_108_499, w_108_500, w_108_540, w_108_549, w_108_591, w_108_652, w_108_673, w_108_693, w_108_705, w_108_717, w_108_731, w_108_734;
  wire w_109_030, w_109_032, w_109_039, w_109_046, w_109_057, w_109_073, w_109_077, w_109_097, w_109_105, w_109_143, w_109_145, w_109_162, w_109_164, w_109_167, w_109_175, w_109_177, w_109_180, w_109_182, w_109_184, w_109_189, w_109_196, w_109_206, w_109_208, w_109_222, w_109_277, w_109_280, w_109_296, w_109_313, w_109_330, w_109_335, w_109_340, w_109_373;
  wire w_110_026, w_110_095, w_110_168, w_110_201, w_110_216, w_110_237, w_110_254, w_110_289, w_110_293, w_110_297, w_110_308, w_110_329, w_110_340, w_110_430, w_110_471, w_110_529, w_110_582, w_110_610, w_110_625, w_110_803, w_110_835, w_110_857, w_110_862, w_110_905, w_110_914, w_110_975, w_110_981, w_110_1010, w_110_1241, w_110_1345, w_110_1372, w_110_1446, w_110_1479, w_110_1502, w_110_1508, w_110_1611, w_110_1612, w_110_1613, w_110_1614, w_110_1615, w_110_1616, w_110_1617, w_110_1621, w_110_1622, w_110_1623, w_110_1624, w_110_1625, w_110_1626, w_110_1627, w_110_1628, w_110_1629, w_110_1630, w_110_1631, w_110_1633;
  wire w_111_000, w_111_029, w_111_030, w_111_069, w_111_080, w_111_085, w_111_122, w_111_125, w_111_151, w_111_153, w_111_168, w_111_204, w_111_239, w_111_251, w_111_256, w_111_263, w_111_264, w_111_289, w_111_292, w_111_331, w_111_333, w_111_343, w_111_352, w_111_376, w_111_383, w_111_417, w_111_418, w_111_426, w_111_447, w_111_482, w_111_485, w_111_509, w_111_604, w_111_632, w_111_666, w_111_679, w_111_712;
  wire w_112_022, w_112_034, w_112_109, w_112_137, w_112_166, w_112_191, w_112_215, w_112_254, w_112_274, w_112_279, w_112_296, w_112_301, w_112_350, w_112_359, w_112_391, w_112_416, w_112_465, w_112_514, w_112_552, w_112_554, w_112_596, w_112_597, w_112_602, w_112_605, w_112_631, w_112_635, w_112_677, w_112_707, w_112_716, w_112_756, w_112_770, w_112_804, w_112_815, w_112_831, w_112_850, w_112_865, w_112_987;
  wire w_113_007, w_113_013, w_113_053, w_113_093, w_113_097, w_113_148, w_113_176, w_113_293, w_113_372, w_113_390, w_113_432, w_113_438, w_113_458, w_113_464, w_113_469, w_113_526, w_113_555, w_113_575, w_113_692, w_113_708, w_113_764, w_113_769, w_113_771, w_113_814, w_113_832, w_113_869, w_113_910, w_113_925, w_113_979, w_113_1021;
  wire w_114_000, w_114_007, w_114_015, w_114_020, w_114_062, w_114_116, w_114_126, w_114_129, w_114_161, w_114_207, w_114_231, w_114_252, w_114_290, w_114_294, w_114_302, w_114_355, w_114_435, w_114_479, w_114_490, w_114_511, w_114_541, w_114_572, w_114_613, w_114_627, w_114_632, w_114_658, w_114_732, w_114_785, w_114_885, w_114_1015, w_114_1047, w_114_1175, w_114_1212, w_114_1247, w_114_1318;
  wire w_115_014, w_115_017, w_115_020, w_115_066, w_115_079, w_115_111, w_115_112, w_115_129, w_115_212, w_115_286, w_115_295, w_115_296, w_115_321, w_115_333, w_115_376, w_115_388, w_115_405, w_115_410, w_115_413, w_115_416, w_115_420, w_115_429, w_115_432, w_115_434, w_115_460, w_115_501, w_115_508, w_115_509, w_115_524, w_115_540, w_115_559, w_115_569, w_115_579, w_115_598, w_115_603, w_115_627;
  wire w_116_086, w_116_103, w_116_115, w_116_188, w_116_228, w_116_359, w_116_364, w_116_386, w_116_390, w_116_395, w_116_409, w_116_421, w_116_436, w_116_454, w_116_599, w_116_670, w_116_730, w_116_805, w_116_878, w_116_901, w_116_912, w_116_959, w_116_1036, w_116_1050, w_116_1268, w_116_1342, w_116_1364, w_116_1463, w_116_1491, w_116_1531, w_116_1549, w_116_1550, w_116_1551, w_116_1552, w_116_1553, w_116_1554, w_116_1555, w_116_1556, w_116_1557, w_116_1558, w_116_1562, w_116_1563, w_116_1564, w_116_1565, w_116_1566, w_116_1567, w_116_1568, w_116_1569, w_116_1570, w_116_1571, w_116_1572, w_116_1574;
  wire w_117_012, w_117_017, w_117_028, w_117_052, w_117_099, w_117_142, w_117_148, w_117_179, w_117_353, w_117_365, w_117_394, w_117_412, w_117_428, w_117_474, w_117_492, w_117_498, w_117_499, w_117_532, w_117_539, w_117_559, w_117_570, w_117_589, w_117_633, w_117_651, w_117_762, w_117_767, w_117_827, w_117_844, w_117_872, w_117_997, w_117_1219, w_117_1471;
  wire w_118_004, w_118_125, w_118_129, w_118_143, w_118_152, w_118_222, w_118_228, w_118_232, w_118_233, w_118_264, w_118_268, w_118_342, w_118_360, w_118_465, w_118_481, w_118_540, w_118_650, w_118_651, w_118_664, w_118_692, w_118_710, w_118_721, w_118_784, w_118_795, w_118_921, w_118_923, w_118_945, w_118_1006, w_118_1036, w_118_1079, w_118_1137, w_118_1139;
  wire w_119_026, w_119_078, w_119_276, w_119_341, w_119_395, w_119_400, w_119_410, w_119_440, w_119_455, w_119_483, w_119_536, w_119_587, w_119_616, w_119_642, w_119_783, w_119_797, w_119_798, w_119_815, w_119_894, w_119_924, w_119_989, w_119_1092, w_119_1112, w_119_1202, w_119_1223, w_119_1278, w_119_1282, w_119_1318, w_119_1341, w_119_1484, w_119_1518;
  wire w_120_000, w_120_002, w_120_010, w_120_032, w_120_035, w_120_037, w_120_041, w_120_043, w_120_047, w_120_051, w_120_057, w_120_085, w_120_086, w_120_094, w_120_104, w_120_109, w_120_111, w_120_116, w_120_117, w_120_118, w_120_127, w_120_128, w_120_133, w_120_141, w_120_152, w_120_156, w_120_165, w_120_168, w_120_172;
  wire w_121_053, w_121_092, w_121_102, w_121_103, w_121_114, w_121_154, w_121_202, w_121_216, w_121_231, w_121_240, w_121_339, w_121_356, w_121_390, w_121_417, w_121_422, w_121_486, w_121_501, w_121_517, w_121_524, w_121_656, w_121_697, w_121_704, w_121_710, w_121_711, w_121_723, w_121_744, w_121_779;
  wire w_122_002, w_122_018, w_122_063, w_122_082, w_122_088, w_122_098, w_122_102, w_122_127, w_122_129, w_122_175, w_122_177, w_122_202, w_122_259, w_122_274, w_122_327, w_122_331, w_122_364, w_122_390, w_122_399, w_122_410, w_122_436, w_122_478, w_122_532, w_122_556, w_122_570, w_122_572, w_122_601, w_122_605;
  wire w_123_000, w_123_004, w_123_063, w_123_088, w_123_134, w_123_182, w_123_237, w_123_334, w_123_346, w_123_374, w_123_399, w_123_400, w_123_428, w_123_455, w_123_478, w_123_494, w_123_508, w_123_518, w_123_590, w_123_615, w_123_616, w_123_618, w_123_627, w_123_668, w_123_792, w_123_832, w_123_865, w_123_970, w_123_984, w_123_990, w_123_1084, w_123_1098, w_123_1121, w_123_1173, w_123_1252;
  wire w_124_046, w_124_048, w_124_061, w_124_064, w_124_083, w_124_111, w_124_112, w_124_135, w_124_142, w_124_152, w_124_155, w_124_165, w_124_223, w_124_260, w_124_274, w_124_280, w_124_377, w_124_381, w_124_387, w_124_393, w_124_457, w_124_466, w_124_488, w_124_489, w_124_662, w_124_740;
  wire w_125_047, w_125_095, w_125_105, w_125_175, w_125_221, w_125_252, w_125_354, w_125_362, w_125_394, w_125_397, w_125_448, w_125_526, w_125_545, w_125_560, w_125_683, w_125_733, w_125_811, w_125_840, w_125_887, w_125_956, w_125_981, w_125_1050, w_125_1055, w_125_1126, w_125_1201, w_125_1361, w_125_1449;
  wire w_126_001, w_126_004, w_126_039, w_126_083, w_126_105, w_126_106, w_126_111, w_126_122, w_126_138, w_126_139, w_126_165, w_126_173, w_126_177, w_126_181, w_126_199, w_126_220, w_126_243, w_126_256, w_126_270, w_126_284, w_126_295, w_126_305, w_126_330, w_126_344, w_126_363, w_126_389, w_126_403, w_126_420;
  wire w_127_186, w_127_251, w_127_298, w_127_307, w_127_372, w_127_399, w_127_426, w_127_476, w_127_482, w_127_516, w_127_624, w_127_697, w_127_734, w_127_783, w_127_802, w_127_807, w_127_866, w_127_889, w_127_932, w_127_1024;
  wire w_128_002, w_128_008, w_128_012, w_128_031, w_128_033, w_128_038, w_128_058, w_128_061, w_128_083, w_128_084, w_128_091, w_128_109, w_128_112, w_128_116, w_128_133, w_128_168, w_128_170, w_128_176, w_128_191, w_128_197, w_128_207, w_128_222, w_128_242, w_128_243, w_128_246, w_128_258, w_128_259, w_128_264;
  wire w_129_010, w_129_041, w_129_066, w_129_090, w_129_245, w_129_332, w_129_368, w_129_429, w_129_518, w_129_607, w_129_608, w_129_648, w_129_675, w_129_681, w_129_744, w_129_747, w_129_783, w_129_795, w_129_808, w_129_877;
  wire w_130_000, w_130_029, w_130_035, w_130_055, w_130_110, w_130_143, w_130_152, w_130_195, w_130_212, w_130_221, w_130_259, w_130_333, w_130_347, w_130_499, w_130_508, w_130_562, w_130_648, w_130_696, w_130_700, w_130_707, w_130_721, w_130_977;
  wire w_131_011, w_131_031, w_131_038, w_131_070, w_131_071, w_131_127, w_131_169, w_131_311, w_131_329, w_131_345, w_131_370, w_131_374, w_131_376, w_131_405, w_131_410, w_131_440, w_131_538, w_131_539, w_131_562, w_131_592, w_131_634, w_131_766, w_131_803, w_131_847, w_131_901, w_131_968, w_131_981, w_131_1014;
  wire w_132_001, w_132_004, w_132_007, w_132_009, w_132_011, w_132_012, w_132_013, w_132_015, w_132_017, w_132_021, w_132_025, w_132_028, w_132_029, w_132_031, w_132_032, w_132_033, w_132_034, w_132_039, w_132_042, w_132_043, w_132_046, w_132_051, w_132_055, w_132_057, w_132_063, w_132_065, w_132_068, w_132_072, w_132_079, w_132_085, w_132_087, w_132_089, w_132_096, w_132_104;
  wire w_133_036, w_133_042, w_133_081, w_133_138, w_133_147, w_133_170, w_133_214, w_133_267, w_133_293, w_133_303, w_133_320, w_133_345, w_133_374, w_133_392, w_133_411, w_133_475, w_133_543, w_133_656, w_133_657, w_133_719, w_133_737, w_133_739, w_133_761, w_133_813, w_133_853, w_133_907;
  wire w_134_006, w_134_012, w_134_019, w_134_096, w_134_097, w_134_135, w_134_150, w_134_254, w_134_295, w_134_321, w_134_352, w_134_375, w_134_414, w_134_430, w_134_468, w_134_477, w_134_487, w_134_804, w_134_828, w_134_893, w_134_944, w_134_1109, w_134_1192, w_134_1230;
  wire w_135_004, w_135_018, w_135_073, w_135_078, w_135_103, w_135_114, w_135_145, w_135_160, w_135_182, w_135_221, w_135_226, w_135_258, w_135_304, w_135_336, w_135_346, w_135_378, w_135_385, w_135_387, w_135_459, w_135_482, w_135_506, w_135_553, w_135_570, w_135_601, w_135_606;
  wire w_136_049, w_136_080, w_136_086, w_136_160, w_136_168, w_136_223, w_136_321, w_136_402, w_136_458, w_136_501, w_136_504, w_136_511, w_136_629, w_136_661, w_136_665, w_136_769, w_136_806, w_136_823, w_136_898;
  wire w_137_007, w_137_012, w_137_039, w_137_112, w_137_146, w_137_178, w_137_239, w_137_276, w_137_339, w_137_344, w_137_355, w_137_379, w_137_389, w_137_399, w_137_417, w_137_449, w_137_463, w_137_507, w_137_514, w_137_653, w_137_735, w_137_871, w_137_952;
  wire w_138_004, w_138_005, w_138_007, w_138_008, w_138_010, w_138_013, w_138_017, w_138_031, w_138_040, w_138_041, w_138_044, w_138_049, w_138_058, w_138_064, w_138_067, w_138_100, w_138_101, w_138_106, w_138_109, w_138_111, w_138_132, w_138_135, w_138_142, w_138_151, w_138_160, w_138_172;
  wire w_139_001, w_139_066, w_139_069, w_139_070, w_139_076, w_139_102, w_139_120, w_139_129, w_139_156, w_139_244, w_139_283, w_139_348, w_139_404, w_139_516, w_139_580, w_139_697, w_139_715, w_139_942, w_139_952, w_139_1104, w_139_1263, w_139_1326, w_139_1379, w_139_1455, w_139_1525, w_139_1723, w_139_1735;
  wire w_140_045, w_140_067, w_140_100, w_140_212, w_140_267, w_140_376, w_140_406, w_140_442, w_140_483, w_140_529, w_140_548, w_140_570, w_140_691, w_140_745, w_140_799, w_140_948, w_140_1319, w_140_1423, w_140_1554, w_140_1596;
  wire w_141_004, w_141_009, w_141_024, w_141_046, w_141_060, w_141_070, w_141_073, w_141_076, w_141_077, w_141_106, w_141_123, w_141_140, w_141_148, w_141_180, w_141_255, w_141_261, w_141_267, w_141_297, w_141_328, w_141_336, w_141_369, w_141_495, w_141_542, w_141_591, w_141_606, w_141_636, w_141_720;
  wire w_142_022, w_142_050, w_142_140, w_142_170, w_142_237, w_142_279, w_142_340, w_142_350, w_142_457, w_142_544, w_142_557, w_142_565, w_142_644, w_142_649, w_142_697, w_142_752, w_142_776, w_142_945, w_142_1185;
  wire w_143_056, w_143_098, w_143_103, w_143_109, w_143_110, w_143_116, w_143_323, w_143_328, w_143_347, w_143_363, w_143_370, w_143_404, w_143_466, w_143_515, w_143_753, w_143_941, w_143_988, w_143_1303, w_143_1344, w_143_1469, w_143_1478, w_143_1529;
  wire w_144_014, w_144_044, w_144_058, w_144_077, w_144_139, w_144_147, w_144_197, w_144_271, w_144_274, w_144_352, w_144_511, w_144_609, w_144_688, w_144_703, w_144_704, w_144_726, w_144_763, w_144_874, w_144_965, w_144_993, w_144_1040, w_144_1102, w_144_1115, w_144_1212, w_144_1226, w_144_1387, w_144_1570;
  wire w_145_005, w_145_006, w_145_007, w_145_009, w_145_012, w_145_013, w_145_015, w_145_016, w_145_017, w_145_020, w_145_023, w_145_024, w_145_027, w_145_032, w_145_033, w_145_034, w_145_035, w_145_036, w_145_037, w_145_038, w_145_040;
  wire w_146_007, w_146_028, w_146_055, w_146_057, w_146_071, w_146_075, w_146_115, w_146_120, w_146_134, w_146_191, w_146_199, w_146_202, w_146_220, w_146_232, w_146_234, w_146_260, w_146_297, w_146_335, w_146_366, w_146_375, w_146_395, w_146_401, w_146_403, w_146_407, w_146_418, w_146_424;
  wire w_147_008, w_147_030, w_147_036, w_147_040, w_147_041, w_147_049, w_147_053, w_147_066, w_147_074, w_147_076, w_147_080, w_147_093, w_147_105, w_147_126, w_147_153, w_147_156, w_147_159, w_147_176, w_147_189, w_147_190, w_147_198;
  wire w_148_120, w_148_274, w_148_490, w_148_530, w_148_715, w_148_806, w_148_903, w_148_932, w_148_1020, w_148_1416, w_148_1503, w_148_1730, w_148_1796, w_148_1819, w_148_1863, w_148_1903, w_148_1915, w_148_1916, w_148_1917, w_148_1918, w_148_1919, w_148_1920, w_148_1921, w_148_1922, w_148_1923, w_148_1924, w_148_1925;
  wire w_149_028, w_149_076, w_149_090, w_149_093, w_149_095, w_149_218, w_149_252, w_149_309, w_149_329, w_149_381, w_149_489, w_149_580, w_149_581, w_149_590, w_149_594, w_149_805, w_149_1027, w_149_1111, w_149_1125, w_149_1158;
  wire w_150_006, w_150_016, w_150_106, w_150_128, w_150_144, w_150_229, w_150_421, w_150_493, w_150_654, w_150_715, w_150_768, w_150_817, w_150_849, w_150_894, w_150_1118, w_150_1283, w_150_1395, w_150_1409, w_150_1570, w_150_1648, w_150_1721, w_150_1759, w_150_1761;
  wire w_151_097, w_151_103, w_151_165, w_151_179, w_151_190, w_151_350, w_151_370, w_151_380, w_151_434, w_151_454, w_151_553, w_151_587, w_151_595, w_151_694, w_151_765, w_151_834, w_151_922, w_151_1014, w_151_1043, w_151_1090, w_151_1109, w_151_1182, w_151_1310, w_151_1378;
  wire w_152_031, w_152_039, w_152_045, w_152_065, w_152_081, w_152_120, w_152_142, w_152_169, w_152_176, w_152_177, w_152_216, w_152_220, w_152_249, w_152_253, w_152_345, w_152_358, w_152_367, w_152_417, w_152_430, w_152_510, w_152_511;
  wire w_153_143, w_153_156, w_153_162, w_153_233, w_153_356, w_153_373, w_153_475, w_153_496, w_153_505, w_153_641, w_153_728, w_153_745, w_153_814, w_153_843, w_153_886, w_153_1016, w_153_1254, w_153_1324;
  wire w_154_000, w_154_008, w_154_013, w_154_015, w_154_051, w_154_066, w_154_071, w_154_073, w_154_096, w_154_098, w_154_106, w_154_112, w_154_123, w_154_124, w_154_136, w_154_142, w_154_148, w_154_171, w_154_181, w_154_182;
  wire w_155_006, w_155_073, w_155_074, w_155_174, w_155_207, w_155_284, w_155_561, w_155_762, w_155_784, w_155_805, w_155_838, w_155_982, w_155_1152, w_155_1257, w_155_1682;
  wire w_156_023, w_156_038, w_156_041, w_156_059, w_156_065, w_156_124, w_156_132, w_156_160, w_156_193, w_156_322, w_156_348, w_156_359, w_156_368, w_156_447, w_156_471, w_156_497, w_156_524, w_156_558, w_156_598;
  wire w_157_020, w_157_040, w_157_065, w_157_174, w_157_188, w_157_230, w_157_337, w_157_357, w_157_405, w_157_489, w_157_563, w_157_739, w_157_762, w_157_993, w_157_1078, w_157_1082, w_157_1161, w_157_1237;
  wire w_158_036, w_158_042, w_158_074, w_158_092, w_158_094, w_158_099, w_158_122, w_158_162, w_158_180, w_158_205, w_158_257, w_158_277, w_158_336, w_158_355, w_158_358, w_158_371, w_158_375;
  wire w_159_149, w_159_186, w_159_215, w_159_336, w_159_344, w_159_596, w_159_767, w_159_802, w_159_806, w_159_842, w_159_858, w_159_974, w_159_1151, w_159_1268, w_159_1288;
  wire w_160_009, w_160_016, w_160_041, w_160_053, w_160_082, w_160_100, w_160_145, w_160_154, w_160_196, w_160_212, w_160_220, w_160_228, w_160_237, w_160_337, w_160_339;
  wire w_161_027, w_161_029, w_161_072, w_161_116, w_161_120, w_161_121, w_161_171, w_161_175, w_161_178, w_161_200, w_161_250, w_161_272, w_161_298, w_161_328, w_161_368, w_161_455, w_161_515, w_161_520;
  wire w_162_019, w_162_027, w_162_093, w_162_105, w_162_117, w_162_130, w_162_242, w_162_278, w_162_340, w_162_591, w_162_746, w_162_795, w_162_808, w_162_813, w_162_890, w_162_894, w_162_904;
  wire w_163_015, w_163_041, w_163_147, w_163_216, w_163_272, w_163_290, w_163_331, w_163_614, w_163_779, w_163_790, w_163_792, w_163_1322, w_163_1548, w_163_1558, w_163_1572, w_163_1585, w_163_1642;
  wire w_164_034, w_164_060, w_164_070, w_164_078, w_164_093, w_164_134, w_164_146, w_164_204, w_164_269, w_164_307, w_164_337, w_164_359, w_164_369, w_164_498, w_164_565, w_164_732, w_164_761, w_164_782, w_164_795, w_164_888;
  wire w_165_030, w_165_058, w_165_106, w_165_130, w_165_136, w_165_163, w_165_170, w_165_227, w_165_253, w_165_264;
  wire w_166_048, w_166_057, w_166_104, w_166_148, w_166_162, w_166_227, w_166_233, w_166_249, w_166_333, w_166_335, w_166_509, w_166_531, w_166_597, w_166_615, w_166_628, w_166_656, w_166_699, w_166_812;
  wire w_167_004, w_167_006, w_167_010, w_167_012, w_167_026, w_167_028, w_167_033, w_167_054, w_167_055, w_167_059, w_167_071, w_167_079, w_167_088, w_167_089, w_167_102, w_167_127, w_167_132;
  wire w_168_005, w_168_035, w_168_077, w_168_225, w_168_240, w_168_259, w_168_320, w_168_341, w_168_399, w_168_402, w_168_470, w_168_529, w_168_608, w_168_649;
  wire w_169_068, w_169_241, w_169_308, w_169_372, w_169_408, w_169_480, w_169_499, w_169_507, w_169_548, w_169_577, w_169_676, w_169_742, w_169_1109, w_169_1242, w_169_1286, w_169_1320;
  wire w_170_045, w_170_095, w_170_167, w_170_196, w_170_322, w_170_364, w_170_623, w_170_642, w_170_766, w_170_819, w_170_903, w_170_947, w_170_988, w_170_991, w_170_1050, w_170_1270, w_170_1475, w_170_1654, w_170_1720, w_170_1727, w_170_1808, w_170_1844;
  wire w_171_037, w_171_053, w_171_085, w_171_095, w_171_101, w_171_109, w_171_112, w_171_152, w_171_237, w_171_267, w_171_290, w_171_471, w_171_493, w_171_505, w_171_539, w_171_593, w_171_654, w_171_704, w_171_731, w_171_750, w_171_794, w_171_858, w_171_971, w_171_1112;
  wire w_172_003, w_172_004, w_172_015, w_172_046, w_172_059, w_172_071, w_172_081, w_172_087, w_172_088, w_172_095, w_172_119, w_172_120, w_172_131, w_172_145, w_172_150;
  wire w_173_079, w_173_112, w_173_258, w_173_425, w_173_447, w_173_470, w_173_537, w_173_558, w_173_569, w_173_612, w_173_762, w_173_948, w_173_991, w_173_1074, w_173_1159;
  wire w_174_048, w_174_073, w_174_078, w_174_324, w_174_370, w_174_380, w_174_392, w_174_401, w_174_581, w_174_624, w_174_675, w_174_742, w_174_780;
  wire w_175_047, w_175_050, w_175_062, w_175_064, w_175_066, w_175_076, w_175_080, w_175_084, w_175_088, w_175_090, w_175_091, w_175_094, w_175_102, w_175_110, w_175_111;
  wire w_176_041, w_176_168, w_176_212, w_176_355, w_176_366, w_176_396, w_176_449, w_176_513, w_176_700, w_176_763, w_176_823, w_176_863, w_176_1151, w_176_1327, w_176_1462;
  wire w_177_208, w_177_222, w_177_782, w_177_900, w_177_917, w_177_1001, w_177_1126, w_177_1191, w_177_1314, w_177_1547, w_177_1601, w_177_1639, w_177_1895;
  wire w_178_031, w_178_032, w_178_123, w_178_285, w_178_361, w_178_365, w_178_455, w_178_479, w_178_552, w_178_586, w_178_635, w_178_658;
  wire w_179_029, w_179_031, w_179_116, w_179_122, w_179_222, w_179_226, w_179_260, w_179_351, w_179_361, w_179_397, w_179_717, w_179_748, w_179_807, w_179_974, w_179_1212, w_179_1221, w_179_1418, w_179_1432, w_179_1625;
  wire w_180_015, w_180_040, w_180_056, w_180_132, w_180_179, w_180_239, w_180_291, w_180_313, w_180_322, w_180_336, w_180_352, w_180_356, w_180_418, w_180_422, w_180_443, w_180_447, w_180_482, w_180_529, w_180_551, w_180_572, w_180_575;
  wire w_181_001, w_181_095, w_181_202, w_181_306, w_181_478, w_181_622, w_181_782, w_181_839, w_181_849, w_181_1114;
  wire w_182_019, w_182_066, w_182_109, w_182_157, w_182_194, w_182_234, w_182_241, w_182_243, w_182_285, w_182_309, w_182_361, w_182_398, w_182_401, w_182_439;
  wire w_183_035, w_183_051, w_183_054, w_183_130, w_183_147, w_183_273, w_183_299, w_183_362, w_183_438, w_183_455, w_183_481, w_183_686, w_183_740, w_183_998, w_183_1020, w_183_1069, w_183_1281, w_183_1551, w_183_1567, w_183_1770, w_183_1773, w_183_1795;
  wire w_184_001, w_184_002, w_184_003, w_184_004, w_184_006, w_184_007, w_184_008, w_184_009, w_184_010;
  wire w_185_077, w_185_333, w_185_506, w_185_943, w_185_1010, w_185_1161, w_185_1466, w_185_1801, w_185_1853;
  wire w_186_000, w_186_011, w_186_015, w_186_025, w_186_064, w_186_119, w_186_151, w_186_162, w_186_165, w_186_180, w_186_191, w_186_203, w_186_295, w_186_307, w_186_315, w_186_332, w_186_344, w_186_379, w_186_385;
  wire w_187_067, w_187_075, w_187_078, w_187_081, w_187_222, w_187_243, w_187_263, w_187_264, w_187_270, w_187_330, w_187_346, w_187_394, w_187_411, w_187_436;
  wire w_188_057, w_188_082, w_188_159, w_188_178, w_188_238, w_188_247, w_188_313, w_188_329, w_188_384, w_188_417, w_188_436, w_188_553;
  wire w_189_010, w_189_011, w_189_015, w_189_019, w_189_024, w_189_026, w_189_043, w_189_052;
  wire w_190_004, w_190_036, w_190_121, w_190_135, w_190_391, w_190_479, w_190_664, w_190_1082, w_190_1290, w_190_1332, w_190_1392, w_190_1437, w_190_1779, w_190_1780;
  wire w_191_076, w_191_098, w_191_138, w_191_221, w_191_270, w_191_375, w_191_445, w_191_626, w_191_793, w_191_816, w_191_841, w_191_1010, w_191_1058, w_191_1112, w_191_1190, w_191_1216, w_191_1390, w_191_1487, w_191_1753;
  wire w_192_087, w_192_089, w_192_108, w_192_118, w_192_190, w_192_318, w_192_328, w_192_338, w_192_346, w_192_359, w_192_382, w_192_428, w_192_461, w_192_473, w_192_486;
  wire w_193_008, w_193_032, w_193_095, w_193_139, w_193_173, w_193_179, w_193_189, w_193_336, w_193_422;
  wire w_194_074, w_194_103, w_194_234, w_194_257, w_194_467, w_194_552, w_194_580, w_194_643, w_194_705, w_194_797, w_194_853, w_194_862;
  wire w_195_041, w_195_079, w_195_086, w_195_194, w_195_202, w_195_311, w_195_410, w_195_498, w_195_1310, w_195_1332, w_195_1391, w_195_1485;
  wire w_196_050, w_196_160, w_196_282, w_196_289, w_196_349, w_196_432, w_196_440, w_196_463, w_196_555, w_196_697;
  wire w_197_073, w_197_082, w_197_288, w_197_296, w_197_493, w_197_707, w_197_777, w_197_860, w_197_1015, w_197_1036, w_197_1099, w_197_1182;
  wire w_198_122, w_198_198, w_198_224, w_198_290, w_198_398, w_198_481, w_198_625, w_198_923, w_198_926, w_198_1118, w_198_1152, w_198_1352, w_198_1377, w_198_1645, w_198_1667, w_198_1676, w_198_1725;
  wire w_199_005, w_199_041, w_199_095, w_199_127, w_199_480, w_199_620, w_199_771, w_199_865, w_199_989, w_199_1086, w_199_1092, w_199_1351, w_199_1604, w_199_1644;
  wire w_200_051, w_200_056, w_200_067, w_200_137, w_200_143, w_200_145, w_200_163, w_200_197, w_200_278, w_200_293, w_200_312, w_200_317, w_200_341, w_200_386, w_200_395, w_200_406, w_200_422, w_200_432;
  wire w_201_006, w_201_021, w_201_025, w_201_029, w_201_031, w_201_033, w_201_058, w_201_059, w_201_117, w_201_130, w_201_166, w_201_184, w_201_230, w_201_265, w_201_314;
  wire w_202_090, w_202_095, w_202_356, w_202_372, w_202_431, w_202_662, w_202_727, w_202_782, w_202_924, w_202_1120, w_202_1580, w_202_1780;
  wire w_203_305, w_203_384, w_203_566, w_203_599, w_203_650, w_203_766;
  wire w_204_064, w_204_196, w_204_245, w_204_353, w_204_438, w_204_674, w_204_725, w_204_1002, w_204_1159, w_204_1212;
  wire w_205_298, w_205_483, w_205_554, w_205_699, w_205_721, w_205_933, w_205_1143;
  wire w_206_165, w_206_484, w_206_621, w_206_712, w_206_741, w_206_775, w_206_918, w_206_964;
  wire w_207_160, w_207_233, w_207_479, w_207_585, w_207_587, w_207_668, w_207_727, w_207_1006, w_207_1070, w_207_1116, w_207_1312, w_207_1454, w_207_1687;
  wire w_208_175, w_208_304, w_208_305, w_208_324, w_208_518, w_208_573, w_208_663, w_208_702, w_208_813, w_208_912, w_208_1069, w_208_1436;
  wire w_209_000, w_209_084, w_209_174, w_209_313, w_209_517, w_209_638, w_209_764, w_209_1088, w_209_1547, w_209_1548, w_209_1549, w_209_1550, w_209_1551, w_209_1552, w_209_1553, w_209_1554, w_209_1555;
  wire w_210_033, w_210_113, w_210_344, w_210_367, w_210_372, w_210_375, w_210_412, w_210_428, w_210_430, w_210_614, w_210_1039, w_210_1199, w_210_1329;
  wire w_211_021, w_211_042, w_211_043, w_211_104, w_211_155, w_211_212, w_211_294, w_211_336, w_211_365;
  wire w_212_009, w_212_066, w_212_134, w_212_332, w_212_762, w_212_1185, w_212_1705;
  wire w_213_020, w_213_021, w_213_035, w_213_041, w_213_152, w_213_172, w_213_342, w_213_379, w_213_423, w_213_469, w_213_512, w_213_562, w_213_743;
  wire w_214_015, w_214_075, w_214_078, w_214_082, w_214_230, w_214_277, w_214_282, w_214_392, w_214_394, w_214_401, w_214_469, w_214_542, w_214_558, w_214_568, w_214_620, w_214_697, w_214_704, w_214_754;
  wire w_215_125, w_215_143, w_215_199, w_215_746, w_215_1078;
  wire w_216_232, w_216_236, w_216_266, w_216_299, w_216_306, w_216_318, w_216_467, w_216_540, w_216_642, w_216_644, w_216_649, w_216_667, w_216_731, w_216_743, w_216_759, w_216_873, w_216_1118, w_216_1133;
  wire w_217_005, w_217_007, w_217_023, w_217_031, w_217_072, w_217_073, w_217_076, w_217_186, w_217_197, w_217_203;
  wire w_218_058, w_218_066, w_218_302, w_218_338, w_218_385, w_218_388, w_218_404, w_218_555, w_218_637, w_218_640, w_218_721, w_218_739, w_218_783, w_218_833, w_218_1074, w_218_1258;
  wire w_219_020, w_219_036, w_219_172, w_219_184;
  wire w_220_1285;
  wire w_221_482, w_221_531, w_221_1056, w_221_1147;
  wire w_222_066, w_222_116, w_222_411, w_222_545, w_222_633, w_222_642, w_222_818, w_222_957, w_222_1038, w_222_1290;
  wire w_223_022, w_223_179, w_223_221, w_223_272, w_223_338, w_223_536, w_223_721, w_223_990, w_223_1010, w_223_1210, w_223_1368;
  wire w_224_049, w_224_145, w_224_249, w_224_413, w_224_605, w_224_834;
  wire w_225_186, w_225_276, w_225_418, w_225_547, w_225_642, w_225_802, w_225_915, w_225_962;
  wire w_226_005, w_226_239, w_226_257, w_226_276, w_226_350, w_226_439, w_226_477, w_226_631, w_226_639, w_226_655, w_226_665;
  wire w_227_002, w_227_009, w_227_085, w_227_104, w_227_172;
  wire w_228_032, w_228_090, w_228_137, w_228_153, w_228_179, w_228_186, w_228_194;
  wire w_229_071, w_229_075, w_229_192, w_229_279, w_229_1171, w_229_1253, w_229_1356, w_229_1460, w_229_1499, w_229_1590, w_229_1608;
  wire w_230_121, w_230_132, w_230_237, w_230_275, w_230_282, w_230_560, w_230_594, w_230_606, w_230_630;
  wire w_231_023, w_231_482, w_231_484, w_231_978, w_231_1101, w_231_1104, w_231_1239, w_231_1269, w_231_1286, w_231_1321, w_231_1386, w_231_1618, w_231_1772;
  wire w_232_002, w_232_153, w_232_183, w_232_385, w_232_388, w_232_480, w_232_507, w_232_608, w_232_641, w_232_667;
  wire w_233_056, w_233_083, w_233_120, w_233_152, w_233_161, w_233_219, w_233_228, w_233_242, w_233_251, w_233_279;
  wire w_234_011, w_234_048, w_234_255, w_234_284, w_234_445, w_234_462, w_234_587, w_234_664, w_234_819, w_234_1004, w_234_1075, w_234_1138;
  wire w_235_106, w_235_291, w_235_327, w_235_350, w_235_371, w_235_498, w_235_551, w_235_573, w_235_640, w_235_669, w_235_733, w_235_757, w_235_791, w_235_892, w_235_947, w_235_1042, w_235_1043, w_235_1044, w_235_1045, w_235_1046, w_235_1047, w_235_1048, w_235_1052, w_235_1053, w_235_1054, w_235_1055, w_235_1056, w_235_1057, w_235_1058, w_235_1059, w_235_1060, w_235_1062;
  wire w_236_005, w_236_099, w_236_182, w_236_391, w_236_403;
  wire w_237_042, w_237_138, w_237_475, w_237_519, w_237_569, w_237_638, w_237_705, w_237_819;
  wire w_238_062, w_238_073, w_238_085, w_238_139, w_238_143, w_238_272, w_238_332, w_238_366, w_238_425, w_238_509;
  wire w_239_061, w_239_196, w_239_367, w_239_566, w_239_601, w_239_726;
  wire w_240_270, w_240_317, w_240_427, w_240_531, w_240_576, w_240_590, w_240_888, w_240_1305;
  wire w_241_010, w_241_064, w_241_096, w_241_299, w_241_502, w_241_1084, w_241_1472;
  wire w_242_001, w_242_012, w_242_014, w_242_017, w_242_030, w_242_046, w_242_064, w_242_075, w_242_084;
  wire w_243_096, w_243_197, w_243_657, w_243_851, w_243_975, w_243_1061, w_243_1147, w_243_1362, w_243_1460;
  wire w_244_026, w_244_200, w_244_317, w_244_535, w_244_543, w_244_796, w_244_892;
  wire w_245_076, w_245_306, w_245_1128, w_245_1762;
  wire w_246_016, w_246_112, w_246_168, w_246_881, w_246_986, w_246_1367, w_246_1436, w_246_1548, w_246_1608;
  wire w_247_514, w_247_604, w_247_657, w_247_759, w_247_786, w_247_877, w_247_1352, w_247_1659;
  wire w_248_024, w_248_028, w_248_051, w_248_059, w_248_124, w_248_127, w_248_147, w_248_161, w_248_291, w_248_327, w_248_354, w_248_445, w_248_450;
  wire w_249_066, w_249_123, w_249_423, w_249_488, w_249_765, w_249_943;
  wire w_250_051, w_250_116, w_250_183, w_250_207, w_250_208, w_250_222, w_250_245;
  wire w_251_010, w_251_109, w_251_123, w_251_157, w_251_169, w_251_204, w_251_245, w_251_281, w_251_282;
  wire w_252_005, w_252_160, w_252_191, w_252_284, w_252_349, w_252_382, w_252_500, w_252_591, w_252_597, w_252_617, w_252_658;
  wire w_253_001, w_253_003, w_253_005;
  wire w_254_015, w_254_039, w_254_114, w_254_167, w_254_340;
  wire w_255_042, w_255_132, w_255_136, w_255_140, w_255_196, w_255_206, w_255_230, w_255_238;
  wire w_256_060, w_256_122, w_256_321, w_256_362, w_256_421, w_256_436, w_256_496, w_256_516, w_256_553, w_256_557, w_256_622, w_256_894, w_256_915, w_256_943, w_256_957;
  wire w_257_146, w_257_235, w_257_360, w_257_796, w_257_1198, w_257_1239, w_257_1369, w_257_1467;
  wire w_258_154, w_258_178, w_258_378, w_258_413;
  wire w_259_070, w_259_081, w_259_220, w_259_272, w_259_392;
  wire w_260_008, w_260_029, w_260_033, w_260_043, w_260_048;
  wire w_261_075, w_261_128, w_261_168, w_261_278;
  wire w_262_119, w_262_131, w_262_144, w_262_184, w_262_238, w_262_290;
  wire w_263_000, w_263_053, w_263_115, w_263_216, w_263_293, w_263_422, w_263_426, w_263_558;
  wire w_264_021, w_264_181, w_264_257, w_264_337, w_264_425, w_264_430, w_264_435, w_264_438, w_264_518, w_264_556;
  wire w_265_098, w_265_127, w_265_223, w_265_335, w_265_375, w_265_456, w_265_476, w_265_699, w_265_1117, w_265_1327, w_265_1382, w_265_1397;
  wire w_266_035, w_266_061, w_266_233, w_266_295, w_266_332, w_266_478, w_266_497, w_266_543;
  wire w_267_180, w_267_201, w_267_254, w_267_329, w_267_397, w_267_399, w_267_432, w_267_476, w_267_705, w_267_861, w_267_865;
  wire w_268_033, w_268_357, w_268_361, w_268_1259;
  wire w_269_453, w_269_1665, w_269_1751, w_269_1792, w_269_1961, w_269_1979;
  wire w_270_079, w_270_226, w_270_265, w_270_271, w_270_345, w_270_392, w_270_531, w_270_663;
  wire w_271_056, w_271_175, w_271_200, w_271_323, w_271_982;
  wire w_272_054, w_272_095, w_272_366, w_272_662, w_272_679, w_272_972, w_272_974;
  wire w_273_071, w_273_075, w_273_156, w_273_350, w_273_376, w_273_595, w_273_610, w_273_623, w_273_751, w_273_869, w_273_880;
  wire w_274_015, w_274_028, w_274_034, w_274_039, w_274_044, w_274_045, w_274_052, w_274_054, w_274_070, w_274_071, w_274_077;
  wire w_275_027, w_275_365, w_275_392, w_275_420, w_275_427, w_275_486, w_275_490;
  wire w_276_024, w_276_078, w_276_091, w_276_119, w_276_134, w_276_145, w_276_176, w_276_188;
  wire w_277_056, w_277_085, w_277_292;
  wire w_278_052, w_278_414, w_278_502, w_278_723, w_278_772, w_278_946, w_278_1207, w_278_1377;
  wire w_279_118, w_279_187, w_279_205, w_279_250, w_279_362, w_279_544, w_279_570, w_279_589;
  wire w_280_045, w_280_266, w_280_365, w_280_389;
  wire w_281_044, w_281_131, w_281_393, w_281_595, w_281_879, w_281_975;
  wire w_282_305, w_282_474, w_282_537, w_282_707, w_282_1923;
  wire w_283_034, w_283_086, w_283_135, w_283_224, w_283_357, w_283_663, w_283_992, w_283_1042, w_283_1149, w_283_1219, w_283_1343, w_283_1410, w_283_1461, w_283_1561, w_283_1724;
  wire w_284_047, w_284_140, w_284_147, w_284_819, w_284_987, w_284_1406, w_284_1530;
  wire w_285_021, w_285_142, w_285_152, w_285_264, w_285_314, w_285_457, w_285_470, w_285_507, w_285_671;
  wire w_286_076, w_286_086, w_286_163, w_286_239, w_286_530, w_286_531, w_286_538, w_286_539;
  wire w_287_020, w_287_022, w_287_027, w_287_129, w_287_148, w_287_194, w_287_271, w_287_287, w_287_352;
  wire w_288_036, w_288_172, w_288_272, w_288_321, w_288_700, w_288_709, w_288_823;
  wire w_289_199, w_289_281, w_289_377, w_289_398, w_289_817, w_289_856, w_289_921, w_289_1017, w_289_1199;
  wire w_290_007, w_290_095, w_290_110, w_290_217, w_290_254, w_290_399;
  wire w_291_126, w_291_244, w_291_638, w_291_793;
  wire w_292_019, w_292_033, w_292_145, w_292_461, w_292_557, w_292_708, w_292_732, w_292_765, w_292_804, w_292_892;
  wire w_293_147, w_293_212, w_293_441, w_293_464, w_293_484, w_293_535, w_293_608, w_293_660, w_293_759, w_293_875, w_293_989, w_293_1017, w_293_1517;
  wire w_294_087, w_294_252, w_294_314, w_294_499, w_294_564, w_294_630, w_294_813;
  wire w_295_332, w_295_369, w_295_422, w_295_546, w_295_616, w_295_718, w_295_949, w_295_1351, w_295_1365;
  wire w_296_305, w_296_333, w_296_491, w_296_801;
  wire w_297_041, w_297_083, w_297_111;
  wire w_298_387, w_298_578, w_298_675, w_298_828, w_298_1289, w_298_1342, w_298_1674;
  wire w_299_086, w_299_100, w_299_113, w_299_308, w_299_340, w_299_691, w_299_740, w_299_1020, w_299_1159, w_299_1179, w_299_1221, w_299_1489, w_299_1560, w_299_1759, w_299_1760, w_299_1761;
  wire w_300_014, w_300_714, w_300_853, w_300_1378, w_300_1448;
  wire w_301_1084, w_301_1225, w_301_1280, w_301_1829;
  wire w_302_121, w_302_122, w_302_195, w_302_321, w_302_402, w_302_624, w_302_660, w_302_1277, w_302_1591;
  wire w_303_008, w_303_045, w_303_690;
  wire w_304_846, w_304_1341, w_304_1575, w_304_1593;
  wire w_305_000, w_305_006, w_305_008, w_305_011, w_305_012, w_305_018, w_305_019, w_305_020, w_305_021, w_305_022, w_305_023, w_305_024;
  wire w_306_005, w_306_282, w_306_427, w_306_1195, w_306_1228, w_306_1282;
  wire w_307_008, w_307_013, w_307_048, w_307_119, w_307_203, w_307_230, w_307_243, w_307_271, w_307_274;
  wire w_308_235, w_308_256, w_308_281, w_308_457, w_308_778, w_308_1117, w_308_1148;
  wire w_309_001, w_309_086, w_309_136, w_309_174;
  wire w_310_019, w_310_043, w_310_065, w_310_136, w_310_189, w_310_223, w_310_274, w_310_332, w_310_477, w_310_505;
  wire w_311_135, w_311_230, w_311_245, w_311_254, w_311_386, w_311_453, w_311_514, w_311_641;
  wire w_312_054, w_312_133, w_312_146, w_312_162, w_312_218, w_312_425, w_312_514;
  wire w_313_000, w_313_001, w_313_005, w_313_017, w_313_025, w_313_028, w_313_033;
  wire w_314_151, w_314_499;
  wire w_315_093, w_315_232, w_315_234, w_315_444, w_315_445, w_315_556, w_315_720;
  wire w_316_082, w_316_101, w_316_288, w_316_510, w_316_915;
  wire w_317_092, w_317_649, w_317_1030, w_317_1544, w_317_1547, w_317_1606;
  wire w_318_012, w_318_097, w_318_192, w_318_277, w_318_336, w_318_360, w_318_507;
  wire w_319_307, w_319_1589;
  wire w_320_201, w_320_214, w_320_484, w_320_632;
  wire w_321_082, w_321_092, w_321_097, w_321_120, w_321_129, w_321_196;
  wire w_322_112, w_322_143, w_322_296, w_322_1155;
  wire w_323_111, w_323_288, w_323_305, w_323_309, w_323_312, w_323_386, w_323_403, w_323_446, w_323_461;
  wire w_324_008, w_324_092, w_324_105, w_324_145, w_324_183, w_324_469, w_324_530, w_324_742;
  wire w_325_661, w_325_1102, w_325_1215, w_325_1228, w_325_1468, w_325_1534;
  wire w_326_363, w_326_383, w_326_737, w_326_1155;
  wire w_327_290, w_327_428, w_327_516, w_327_519, w_327_1023, w_327_1107;
  wire w_328_005, w_328_006, w_328_008, w_328_010, w_328_013;
  wire w_329_059, w_329_203, w_329_228, w_329_249, w_329_262, w_329_460;
  wire w_330_248, w_330_693, w_330_731, w_330_753, w_330_814, w_330_958, w_330_1024;
  wire w_331_107, w_331_550, w_331_838, w_331_899;
  wire w_332_063, w_332_177, w_332_319, w_332_572, w_332_617, w_332_1090;
  wire w_333_070;
  wire w_334_223, w_334_261, w_334_343, w_334_566, w_334_567, w_334_597, w_334_650;
  wire w_335_006, w_335_072, w_335_362;
  wire w_336_141, w_336_181, w_336_577, w_336_663, w_336_1049, w_336_1116, w_336_1225, w_336_1630;
  wire w_337_027, w_337_038, w_337_094, w_337_158, w_337_234, w_337_266, w_337_369;
  wire w_338_073, w_338_1435, w_338_1654, w_338_1705;
  wire w_339_121, w_339_235, w_339_405, w_339_439, w_339_524;
  wire w_340_114;
  wire w_341_141, w_341_249, w_341_302;
  wire w_342_013, w_342_1028, w_342_1576, w_342_1768, w_342_1769, w_342_1770, w_342_1771, w_342_1772, w_342_1773, w_342_1774, w_342_1775, w_342_1776, w_342_1777, w_342_1781, w_342_1782, w_342_1783, w_342_1784, w_342_1785, w_342_1786, w_342_1788;
  wire w_343_016, w_343_227, w_343_894, w_343_1177;
  wire w_344_052, w_344_117, w_344_139, w_344_141, w_344_150, w_344_207;
  wire w_345_1056, w_345_1240, w_345_1481;
  wire w_346_341, w_346_528, w_346_640, w_346_679;
  wire w_347_053, w_347_705, w_347_950, w_347_1219, w_347_1311, w_347_1576, w_347_1601;
  wire w_348_167;
  wire w_349_052, w_349_104;
  wire w_350_207, w_350_314, w_350_377, w_350_444, w_350_527, w_350_529;
  wire w_351_000, w_351_021, w_351_028, w_351_035;
  wire w_352_320, w_352_406, w_352_422, w_352_672;
  wire w_353_138, w_353_181, w_353_240, w_353_380, w_353_448, w_353_531, w_353_691, w_353_720, w_353_985, w_353_1174;
  wire w_354_064, w_354_278, w_354_391, w_354_412, w_354_460, w_354_1250, w_354_1261;
  wire w_355_018, w_355_076, w_355_089, w_355_155, w_355_213, w_355_226, w_355_291, w_355_525;
  wire w_356_068, w_356_335, w_356_714;
  wire w_357_026, w_357_083, w_357_141, w_357_293, w_357_401;
  wire w_358_471, w_358_675, w_358_692, w_358_1178, w_358_1499;
  wire w_359_131, w_359_526, w_359_650, w_359_1125;
  wire w_360_496, w_360_542, w_360_762;
  wire w_361_090, w_361_238, w_361_317;
  wire w_362_105, w_362_212, w_362_293, w_362_337, w_362_481, w_362_483, w_362_1655;
  wire w_363_075, w_363_507, w_363_598, w_363_803;
  wire w_364_185, w_364_233, w_364_722, w_364_1423;
  wire w_365_064, w_365_198, w_365_216, w_365_534, w_365_536, w_365_620, w_365_832, w_365_858;
  wire w_366_011;
  wire w_367_489;
  wire w_368_156, w_368_455, w_368_653, w_368_783, w_368_986, w_368_1314, w_368_1526, w_368_1696;
  wire w_369_228, w_369_346, w_369_649, w_369_1046, w_369_1193, w_369_1531;
  wire w_370_066, w_370_067, w_370_077, w_370_616, w_370_890, w_370_1007, w_370_1459;
  wire w_371_092, w_371_098, w_371_343, w_371_387, w_371_548, w_371_710;
  wire w_372_215, w_372_317, w_372_366, w_372_404, w_372_428;
  wire w_373_465, w_373_471, w_373_1442, w_373_1800;
  wire w_374_012, w_374_145, w_374_304, w_374_798, w_374_1192, w_374_1496;
  wire w_375_1233;
  wire w_376_209, w_376_513, w_376_677, w_376_750;
  wire w_377_072, w_377_193, w_377_256;
  wire w_378_048, w_378_278, w_378_565, w_378_597;
  wire w_379_043, w_379_194, w_379_781, w_379_829;
  wire w_380_321, w_380_434;
  wire w_381_179, w_381_531, w_381_634, w_381_839;
  wire w_382_163, w_382_185, w_382_653, w_382_672, w_382_678;
  wire w_383_097, w_383_133, w_383_187, w_383_219, w_383_235, w_383_377;
  wire w_384_1443;
  wire w_385_227, w_385_326;
  wire w_386_011, w_386_236;
  wire w_387_317, w_387_619, w_387_691, w_387_720, w_387_967;
  wire w_388_219, w_388_339, w_388_630, w_388_751, w_388_936;
  wire w_389_671, w_389_787, w_389_1252, w_389_1431, w_389_1549, w_389_1637;
  wire w_390_195, w_390_434, w_390_717;
  wire w_391_015, w_391_048;
  wire w_392_480, w_392_598, w_392_982, w_392_1327, w_392_1798;
  wire w_393_523;
  wire w_394_008, w_394_013, w_394_030, w_394_037;
  wire w_395_657, w_395_966;
  wire w_396_001, w_396_254, w_396_282, w_396_560;
  wire w_397_455, w_397_673, w_397_1350, w_397_1463;
  wire w_398_086, w_398_235, w_398_258, w_398_887, w_398_1205, w_398_1585;
  wire w_399_076, w_399_191, w_399_563, w_399_1417, w_399_1788, w_399_1789, w_399_1790, w_399_1791, w_399_1792, w_399_1793, w_399_1794, w_399_1795, w_399_1796, w_399_1797, w_399_1798, w_399_1802, w_399_1803, w_399_1804, w_399_1806;
  wire w_400_067, w_400_224;
  wire w_401_063, w_401_383, w_401_517, w_401_544;
  wire w_402_176, w_402_569, w_402_632, w_402_872, w_402_998;
  wire w_403_004, w_403_097, w_403_146, w_403_215, w_403_223;
  wire w_404_052, w_404_266, w_404_800;
  wire w_405_122, w_405_171, w_405_284;
  wire w_406_175, w_406_471, w_406_554, w_406_677, w_406_835, w_406_870, w_406_964;
  wire w_407_014, w_407_182;
  wire w_408_005, w_408_011, w_408_015, w_408_017;
  wire w_409_138, w_409_623, w_409_732, w_409_773;
  wire w_410_008, w_410_069, w_410_103, w_410_111, w_410_164;
  wire w_411_668, w_411_987, w_411_1244, w_411_1382, w_411_1447;
  wire w_412_000, w_412_028, w_412_161, w_412_437;
  wire w_413_194;
  wire w_414_110;
  wire w_415_024, w_415_058, w_415_207;
  wire w_416_198, w_416_298, w_416_307, w_416_364, w_416_432, w_416_600, w_416_1113;
  wire w_417_017, w_417_456;
  wire w_418_170, w_418_475, w_418_479, w_418_673, w_418_1325, w_418_1382;
  wire w_419_069, w_419_087, w_419_178;
  wire w_420_832, w_420_1439;
  wire w_421_031, w_421_096, w_421_143, w_421_154, w_421_269, w_421_275, w_421_311;
  wire w_422_251, w_422_306, w_422_351, w_422_384, w_422_579;
  wire w_423_080, w_423_206;
  wire w_424_002, w_424_010, w_424_016, w_424_021, w_424_022, w_424_025;
  wire w_425_174, w_425_247;
  wire w_426_621;
  wire w_427_021, w_427_055, w_427_082, w_427_169, w_427_172, w_427_245, w_427_257;
  wire w_428_864;
  wire w_429_200, w_429_1594;
  wire w_430_014, w_430_067, w_430_069, w_430_088, w_430_130;
  wire w_431_218, w_431_239, w_431_1031, w_431_1266;
  wire w_432_171, w_432_726, w_432_727, w_432_728, w_432_729, w_432_730, w_432_731, w_432_735, w_432_736, w_432_737, w_432_738, w_432_739, w_432_741;
  wire w_433_070, w_433_394, w_433_430, w_433_560, w_433_592, w_433_631, w_433_824;
  wire w_434_621, w_434_633;
  wire w_435_916;
  wire w_436_667, w_436_1391, w_436_1601;
  wire w_437_1451, w_437_1574;
  wire w_438_1586;
  wire w_439_508, w_439_531;
  wire w_440_591, w_440_709, w_440_814, w_440_896;
  wire w_441_128, w_441_750, w_441_948;
  wire w_442_118, w_442_759, w_442_803, w_442_1693;
  wire w_443_305, w_443_369, w_443_718;
  wire w_444_085, w_444_113;
  wire w_445_301, w_445_361, w_445_394;
  wire w_446_046, w_446_247, w_446_536, w_446_605, w_446_698, w_446_722, w_446_752;
  wire w_447_169;
  wire w_448_252, w_448_423;
  wire w_449_347, w_449_402, w_449_1041;
  wire w_451_401, w_451_616, w_451_632;
  wire w_452_108, w_452_176, w_452_289, w_452_775;
  wire w_453_073, w_453_109, w_453_115, w_453_196;
  wire w_454_021, w_454_025, w_454_043, w_454_142, w_454_260;
  wire w_456_283, w_456_442, w_456_731, w_456_769, w_456_979;
  wire w_457_975, w_457_1221, w_457_1222, w_457_1223, w_457_1224, w_457_1225, w_457_1226;
  wire w_458_073, w_458_412, w_458_1066;
  wire w_459_383, w_459_833;
  wire w_460_906, w_460_1204;
  wire w_461_047, w_461_171, w_461_280, w_461_310, w_461_319, w_461_651, w_461_696;
  wire w_462_021, w_462_025, w_462_134;
  wire w_463_044, w_463_144, w_463_172, w_463_340, w_463_433, w_463_473;
  wire w_464_379;
  wire w_465_050, w_465_943;
  wire w_466_005, w_466_103, w_466_234, w_466_271;
  wire w_467_390, w_467_689, w_467_1137;
  wire w_468_214, w_468_249, w_468_253;
  wire w_469_046, w_469_351, w_469_529;
  wire w_470_456, w_470_1212;
  wire w_471_265, w_471_359, w_471_553;
  wire w_473_022, w_473_245, w_473_1043;
  wire w_474_300, w_474_412;
  wire w_475_095, w_475_175, w_475_219;
  wire w_476_073, w_476_096, w_476_191, w_476_312, w_476_313, w_476_379, w_476_389;
  wire w_477_023, w_477_098, w_477_104;
  wire w_478_293, w_478_367, w_478_665, w_478_815, w_478_1092, w_478_1191, w_478_1446;
  wire w_479_615, w_479_638, w_479_643, w_479_694, w_479_1024, w_479_1741;
  wire w_480_021, w_480_062;
  wire w_481_093, w_481_1485;
  wire w_482_410, w_482_839;
  wire w_483_094, w_483_314, w_483_425;
  wire w_484_010, w_484_362, w_484_492, w_484_493, w_484_494, w_484_498, w_484_499, w_484_500, w_484_501, w_484_502, w_484_503, w_484_504, w_484_505, w_484_506, w_484_507, w_484_509;
  wire w_485_176;
  wire w_487_032, w_487_525, w_487_617, w_487_790, w_487_1069, w_487_1147;
  wire w_488_278, w_488_641, w_488_908, w_488_978;
  wire w_489_036, w_489_1324, w_489_1344;
  wire w_490_288, w_490_1421;
  wire w_491_048, w_491_164;
  wire w_492_043, w_492_085, w_492_086, w_492_128;
  wire w_493_062, w_493_157, w_493_225, w_493_430, w_493_441, w_493_572, w_493_573, w_493_574, w_493_575, w_493_576, w_493_577, w_493_578, w_493_582, w_493_583, w_493_584, w_493_585, w_493_586, w_493_587, w_493_589;
  wire w_494_945, w_494_1233, w_494_1931, w_494_1932, w_494_1933, w_494_1934, w_494_1935, w_494_1936;
  wire w_495_1004, w_495_1084;
  wire w_496_101, w_496_495, w_496_628, w_496_797, w_496_959, w_496_1215;
  wire w_497_331, w_497_364, w_497_391;
  wire w_498_402, w_498_507, w_498_636;
  wire w_499_181, w_499_371, w_499_436, w_499_1419, w_499_1719;
  wire w_500_004, w_500_891, w_500_1299;
  wire w_501_352;
  wire w_502_002, w_502_250, w_502_289;
  wire w_503_023, w_503_261, w_503_299, w_503_404, w_503_694;
  wire w_504_065, w_504_152, w_504_314, w_504_564;
  wire w_505_342, w_505_916, w_505_1503, w_505_1562;
  wire w_506_135, w_506_138, w_506_472;
  wire w_507_047, w_507_110;
  wire w_508_018;
  wire w_509_068, w_509_110, w_509_148, w_509_294, w_509_322, w_509_386;
  wire w_510_051, w_510_177, w_510_180, w_510_260, w_510_261;
  wire w_512_268, w_512_374, w_512_679, w_512_823, w_512_1078;
  wire w_513_409, w_513_1030;
  wire w_514_053, w_514_848, w_514_955, w_514_1099, w_514_1390;
  wire w_515_094, w_515_186, w_515_456, w_515_657, w_515_679;
  wire w_516_317, w_516_699;
  wire w_517_039;
  wire w_518_204;
  wire w_519_189;
  wire w_520_598, w_520_667, w_520_1416;
  wire w_521_852;
  wire w_522_090;
  wire w_523_021, w_523_688;
  wire w_524_121, w_524_464, w_524_1502, w_524_1505;
  wire w_525_175, w_525_366, w_525_1141, w_525_1399;
  wire w_528_041, w_528_110, w_528_145;
  wire w_529_180;
  wire w_530_1263, w_530_1605;
  wire w_531_121, w_531_628, w_531_1378, w_531_1379, w_531_1380, w_531_1381, w_531_1382, w_531_1383, w_531_1384, w_531_1385, w_531_1386, w_531_1387, w_531_1388, w_531_1392, w_531_1393, w_531_1394, w_531_1395, w_531_1397;
  wire w_532_271, w_532_410;
  wire w_534_014, w_534_1008, w_534_1231;
  wire w_536_150;
  wire w_537_388, w_537_615;
  wire w_538_357, w_538_363, w_538_713, w_538_864;
  wire w_539_231;
  wire w_540_182, w_540_326, w_540_341;
  wire w_541_073;
  wire w_542_089, w_542_308;
  wire w_543_374, w_543_594, w_543_740;
  wire w_544_028, w_544_040, w_544_081, w_544_100;
  wire w_545_1135, w_545_1157;
  wire w_546_065, w_546_078, w_546_258, w_546_1098;
  wire w_547_082, w_547_437;
  wire w_548_325, w_548_356, w_548_509, w_548_636, w_548_843, w_548_923;
  wire w_549_164, w_549_222, w_549_244, w_549_284, w_549_352;
  wire w_550_785;
  wire w_551_082, w_551_271, w_551_365, w_551_674, w_551_929, w_551_1193;
  wire w_552_027;
  wire w_554_288, w_554_319;
  wire w_555_332, w_555_481, w_555_1052, w_555_1335, w_555_1534;
  wire w_556_147, w_556_235, w_556_258, w_556_272;
  wire w_557_485, w_557_825, w_557_1075;
  wire w_559_669, w_559_922;
  wire w_560_327, w_560_345, w_560_1113, w_560_1382;
  wire w_561_252, w_561_339;
  wire w_562_017;
  wire w_563_139, w_563_242, w_563_721, w_563_905, w_563_960, w_563_961, w_563_962, w_563_963;
  wire w_564_071;
  wire w_566_066, w_566_957;
  wire w_568_047, w_568_596, w_568_913;
  wire w_569_388;
  wire w_570_560, w_570_1461;
  wire w_571_034, w_571_1088;
  wire w_575_205, w_575_519, w_575_539;
  wire w_576_511, w_576_846, w_576_1032;
  wire w_578_287, w_578_425, w_578_634;
  wire w_579_134, w_579_721, w_579_1003, w_579_1598;
  wire w_582_1282, w_582_1357;
  wire w_583_066, w_583_224, w_583_291;
  wire w_584_730, w_584_893;
  wire w_585_214, w_585_360;
  wire w_586_135, w_586_969, w_586_1406;
  wire w_587_856, w_587_869;
  wire w_588_356;
  wire w_589_707;
  wire w_590_780, w_590_1014;
  wire w_591_300, w_591_762, w_591_1100;
  wire w_592_086, w_592_142, w_592_687;
  wire w_593_207;
  wire w_595_157, w_595_178, w_595_321;
  wire w_596_124, w_596_343;
  wire w_597_068, w_597_813;
  wire w_598_265;
  wire w_599_010, w_599_034, w_599_056;
  wire w_600_523, w_600_663;
  wire w_601_015, w_601_063, w_601_438, w_601_471;
  wire w_602_517;
  wire w_606_070;
  wire w_607_622, w_607_675;
  wire w_609_034, w_609_330;
  wire w_610_889, w_610_890, w_610_891, w_610_892, w_610_893, w_610_894, w_610_895, w_610_896, w_610_897, w_610_898, w_610_899;
  wire w_611_122, w_611_200, w_611_393;
  wire w_613_092, w_613_379, w_613_1491;
  wire w_614_162, w_614_388, w_614_500;
  wire w_615_216;
  wire w_616_164, w_616_1323;
  wire w_617_575, w_617_871;
  wire w_618_405;
  wire w_619_033, w_619_080;
  wire w_620_074, w_620_379;
  wire w_621_071, w_621_268;
  wire w_622_749;
  wire w_623_435, w_623_635;
  wire w_624_1288;
  wire w_625_1222;
  wire w_626_212, w_626_1103;
  wire w_627_1504;
  wire w_628_148, w_628_999, w_628_1376;
  wire w_629_028, w_629_318, w_629_760;
  wire w_630_083, w_630_312;
  wire w_631_069;
  wire w_632_266;
  wire w_633_068, w_633_696;
  wire w_634_237;
  wire w_635_326, w_635_649;
  wire w_636_262, w_636_299;
  wire w_637_159, w_637_508;
  wire w_638_432, w_638_1113, w_638_1129;
  wire w_639_313, w_639_1097, w_639_1572, w_639_1573;
  wire w_640_066, w_640_496, w_640_710;
  wire w_641_262, w_641_515, w_641_594, w_641_787;
  wire w_642_231, w_642_268;
  wire w_644_837, w_644_866;
  wire w_645_049, w_645_091, w_645_105;
  wire w_646_094;
  wire w_647_214, w_647_288;
  wire w_648_062, w_648_1062;
  wire w_649_568;
  wire w_650_134, w_650_173;
  wire w_651_012, w_651_352, w_651_1455, w_651_1483;
  wire w_652_003, w_652_032, w_652_064;
  wire w_654_208;
  wire w_655_134, w_655_1625;
  wire w_657_1324;
  wire w_658_866;
  wire w_659_522;
  wire w_660_005, w_660_064, w_660_207, w_660_223, w_660_298;
  wire w_662_540;
  wire w_663_732;
  wire w_664_091;
  wire w_665_324, w_665_335;
  wire w_667_474;
  wire w_668_104, w_668_967;
  wire w_669_042, w_669_044, w_669_079, w_669_137, w_669_138, w_669_139, w_669_140, w_669_141, w_669_142, w_669_143, w_669_144, w_669_145;
  wire w_670_119, w_670_353, w_670_636;
  wire w_671_330;
  wire w_673_061;
  wire w_674_038, w_674_041, w_674_050;
  wire w_675_004, w_675_012;
  wire w_676_349, w_676_1465;
  wire w_677_132;
  wire w_678_238, w_678_759, w_678_781;
  wire w_679_272, w_679_506;
  wire w_681_026, w_681_1392;
  wire w_682_001, w_682_042, w_682_097, w_682_148;
  wire w_683_161, w_683_164, w_683_238;
  wire w_685_1698;
  wire w_686_073, w_686_417;
  wire w_687_290, w_687_540, w_687_1614;
  wire w_688_909;
  wire w_690_753;
  wire w_691_286, w_691_509;
  wire w_692_115;
  wire w_694_687, w_694_874;
  wire w_696_103, w_696_418, w_696_431;
  wire w_697_644, w_697_733, w_697_939, w_697_1369;
  wire w_698_1173;
  wire w_699_079;
  wire w_700_106, w_700_818;
  wire w_701_276;
  wire w_703_042, w_703_183, w_703_312;
  wire w_704_087, w_704_803, w_704_1453;
  wire w_705_087;
  wire w_706_587, w_706_1392;
  wire w_707_418;
  wire w_708_131, w_708_987, w_708_1216;
  wire w_709_060;
  wire w_711_891;
  wire w_712_441, w_712_442, w_712_634;
  wire w_713_104, w_713_131, w_713_146, w_713_203;
  wire w_714_604;
  wire w_715_306, w_715_605, w_715_843;
  wire w_716_110, w_716_135, w_716_416, w_716_418;
  wire w_717_1135, w_717_1608;
  wire w_719_461;
  wire w_722_1277, w_722_1323, w_722_1621, w_722_1622, w_722_1623, w_722_1624, w_722_1625, w_722_1626, w_722_1627, w_722_1628;
  wire w_723_166;
  wire w_724_167, w_724_444, w_724_1149;
  wire w_726_1725;
  wire w_727_690;
  wire w_728_220, w_728_1474;
  wire w_729_404;
  wire w_730_029, w_730_695;
  wire w_731_027, w_731_059;
  wire w_733_210, w_733_461;
  wire w_737_163;
  wire w_739_100;
  wire w_740_1463;
  wire w_741_660, w_741_921;
  wire w_742_065, w_742_176;
  wire w_743_219;
  wire w_744_084, w_744_349;
  wire w_745_034, w_745_1779;
  wire w_748_059, w_748_137, w_748_352;
  wire w_749_443, w_749_660;
  wire w_751_026;
  wire w_752_789, w_752_1842;
  wire w_755_1157;
  wire w_756_029, w_756_402;
  wire w_758_301, w_758_721;
  wire w_759_359;
  wire w_761_029, w_761_408;
  wire w_762_873, w_762_973;
  wire w_763_252;
  wire w_764_117;
  wire w_766_241;
  wire w_768_099, w_768_1400, w_768_1574;
  wire w_769_203, w_769_204, w_769_205, w_769_206, w_769_207, w_769_208, w_769_209;
  wire w_770_377;
  wire w_771_455;
  wire w_773_045, w_773_106, w_773_158;
  wire w_774_273, w_774_275, w_774_358, w_774_402;
  wire w_777_1423;
  wire w_778_157;
  wire w_779_268, w_779_1214;
  wire w_781_001, w_781_1578, w_781_1927;
  wire w_782_660, w_782_860;
  wire w_783_1101;
  wire w_784_448;
  wire w_786_960, w_786_1041;
  wire w_788_162;
  wire w_789_059;
  wire w_790_373, w_790_894, w_790_1308;
  wire w_791_162;
  wire w_792_882;
  wire w_793_071, w_793_376;
  wire w_794_021, w_794_319;
  wire w_795_080;
  wire w_796_506, w_796_1386, w_796_1672;
  wire w_797_000, w_797_284;
  wire w_798_333, w_798_611;
  wire w_799_494, w_799_848, w_799_849, w_799_850, w_799_851, w_799_852, w_799_853, w_799_854, w_799_855, w_799_856, w_799_860, w_799_861, w_799_862, w_799_863, w_799_865;
  wire w_800_598;
  wire w_803_018, w_803_122, w_803_464;
  wire w_805_553;
  wire w_807_312, w_807_337;
  wire w_808_008, w_808_810, w_808_986;
  wire w_809_122, w_809_1170;
  wire w_810_657, w_810_754, w_810_824;
  wire w_811_1068, w_811_1380, w_811_1552, w_811_1656, w_811_1657, w_811_1658, w_811_1662, w_811_1663, w_811_1664, w_811_1665, w_811_1666, w_811_1667, w_811_1668, w_811_1670;
  wire w_813_1102;
  wire w_814_632;
  wire w_815_878;
  wire w_817_481, w_817_484;
  wire w_818_030, w_818_157;
  wire w_819_177, w_819_178, w_819_190;
  wire w_820_230, w_820_664;
  wire w_821_012;
  wire w_825_278;
  wire w_826_369, w_826_437, w_826_438, w_826_439, w_826_440, w_826_444, w_826_445, w_826_446, w_826_447, w_826_448, w_826_449, w_826_450, w_826_452;
  wire w_827_021, w_827_820;
  wire w_828_066, w_828_715;
  wire w_829_391;
  wire w_830_022;
  wire w_831_1052;
  wire w_832_266;
  wire w_833_562;
  wire w_834_1377;
  wire w_835_622;
  wire w_836_246;
  wire w_838_1026;
  wire w_841_642, w_841_1177, w_841_1412, w_841_1480;
  wire w_842_151;
  wire w_843_173, w_843_278;
  wire w_844_323;
  wire w_845_041;
  wire w_847_251, w_847_421;
  wire w_848_264, w_848_349, w_848_565, w_848_723;
  wire w_849_242;
  wire w_850_1264;
  wire w_851_1288, w_851_1289, w_851_1290, w_851_1291, w_851_1292, w_851_1293, w_851_1294, w_851_1295, w_851_1296, w_851_1297;
  wire w_852_269;
  wire w_855_166, w_855_946;
  wire w_856_1410;
  wire w_858_124, w_858_381;
  wire w_860_017, w_860_405, w_860_903, w_860_1045;
  wire w_862_052;
  wire w_863_096, w_863_292, w_863_389, w_863_390, w_863_391, w_863_392, w_863_393, w_863_394, w_863_398, w_863_399, w_863_400, w_863_401, w_863_402, w_863_403, w_863_404, w_863_405, w_863_406, w_863_407, w_863_408, w_863_409, w_863_411;
  wire w_864_076;
  wire w_865_178;
  wire w_866_722, w_866_1044;
  wire w_868_223;
  wire w_871_000;
  wire w_874_219;
  wire w_876_063, w_876_1135;
  wire w_877_566, w_877_632;
  wire w_880_1190;
  wire w_882_384, w_882_737;
  wire w_885_1687;
  wire w_886_088;
  wire w_888_1871;
  wire w_889_030, w_889_097;
  wire w_890_411, w_890_822;
  wire w_892_214;
  wire w_893_056;
  wire w_894_393, w_894_586, w_894_587, w_894_588, w_894_589, w_894_590, w_894_591, w_894_595, w_894_596, w_894_597, w_894_598, w_894_599, w_894_600, w_894_601, w_894_602, w_894_603, w_894_604, w_894_605, w_894_607;
  wire w_895_037;
  wire w_897_1329, w_897_1330, w_897_1331, w_897_1332, w_897_1333, w_897_1334, w_897_1335, w_897_1336, w_897_1337, w_897_1338;
  wire w_901_088, w_901_574, w_901_607;
  wire w_902_415;
  wire w_903_455;
  wire w_905_262;
  wire w_907_426;
  wire w_908_1300;
  wire w_910_116;
  wire w_911_069;
  wire w_912_120, w_912_152, w_912_239, w_912_1012;
  wire w_915_132, w_915_948;
  wire w_916_191, w_916_732;
  wire w_919_1871, w_919_1872, w_919_1873, w_919_1874, w_919_1875, w_919_1876, w_919_1877, w_919_1878;
  wire w_921_020;
  wire w_922_1398, w_922_1533;
  wire w_924_311;
  wire w_925_563, w_925_784;
  wire w_928_200;
  wire w_932_294, w_932_853;
  wire w_936_1058;
  wire w_937_329;
  wire w_939_556;
  wire w_940_013, w_940_080, w_940_140;
  wire w_941_1118, w_941_1119, w_941_1120;
  wire w_942_113;
  wire w_949_751;
  wire w_951_471;
  wire w_952_247;
  wire w_957_171;
  wire w_962_105;
  wire w_963_263;
  wire w_966_336, w_966_461, w_966_462, w_966_463, w_966_464, w_966_465, w_966_466, w_966_470, w_966_471, w_966_472, w_966_473, w_966_474, w_966_475, w_966_476, w_966_477, w_966_478, w_966_480;
  wire w_968_263, w_968_742;
  wire w_969_298;
  wire w_975_392, w_975_669, w_975_1237;
  wire w_976_215, w_976_287, w_976_288, w_976_289, w_976_290, w_976_291, w_976_292, w_976_293, w_976_294, w_976_295, w_976_299, w_976_300, w_976_301, w_976_303;
  wire w_978_267;
  wire w_979_555, w_979_812;
  wire w_980_107;
  wire w_981_087;
  wire w_987_771;
  wire w_988_096;
  wire w_991_026;
  wire w_996_217, w_996_1460, w_996_1461, w_996_1462, w_996_1463, w_996_1464, w_996_1465, w_996_1466, w_996_1467, w_996_1471, w_996_1472, w_996_1473, w_996_1474, w_996_1475, w_996_1476, w_996_1477, w_996_1478, w_996_1479, w_996_1480, w_996_1482;
  wire w_999_921;
  wire w_1002_108, w_1002_191;
  wire w_1004_487;
  wire w_1005_1726;
  wire w_1006_1160;
  wire w_1010_649;
  wire w_1011_314;
  wire w_1012_147, w_1012_353;
  wire w_1013_326;
  wire w_1017_151, w_1017_222;
  wire w_1018_190, w_1018_418, w_1018_633;
  wire w_1019_850;
  wire w_1025_1532;
  wire w_1030_528;
  wire w_1033_020;
  wire w_1034_506;
  wire w_1035_002, w_1035_074;
  wire w_1036_151, w_1036_805;
  wire w_1038_1382;
  wire w_1041_374;
  wire w_1044_059;
  wire w_1045_096;
  wire w_1047_1404;
  wire w_1049_021;
  wire w_1050_082;
  wire w_1053_806;
  wire w_1055_134, w_1055_453, w_1055_454, w_1055_455, w_1055_456, w_1055_457, w_1055_458, w_1055_459, w_1055_460, w_1055_461, w_1055_462, w_1055_463, w_1055_464;
  wire w_1056_111;
  wire w_1057_865;
  wire w_1060_189;
  wire w_1064_040;
  wire w_1065_185, w_1065_229, w_1065_406;
  wire w_1066_974;
  wire w_1069_285, w_1069_553, w_1069_579;
  wire w_1072_321;
  wire w_1075_1904, w_1075_1905, w_1075_1906, w_1075_1907, w_1075_1908, w_1075_1909, w_1075_1910, w_1075_1911, w_1075_1915, w_1075_1916, w_1075_1917, w_1075_1918, w_1075_1919, w_1075_1920, w_1075_1921, w_1075_1922, w_1075_1924;
  wire w_1076_206;
  wire w_1078_045, w_1078_081, w_1078_082, w_1078_083, w_1078_084, w_1078_085, w_1078_086, w_1078_087, w_1078_088, w_1078_089, w_1078_090, w_1078_091, w_1078_092;
  wire w_1080_723;
  wire w_1083_094;
  wire w_1087_369;
  wire w_1088_775, w_1088_842;
  wire w_1092_449;
  wire w_1093_019, w_1093_049;
  wire w_1095_044;
  wire w_1097_525, w_1097_1090;
  wire w_1099_048;
  wire w_1104_019;
  wire w_1108_010;
  wire w_1109_060;
  wire w_1111_1175;
  wire w_1112_1168, w_1112_1748, w_1112_1749, w_1112_1750, w_1112_1751, w_1112_1752, w_1112_1753, w_1112_1754, w_1112_1755, w_1112_1756;
  wire w_1114_194;
  wire w_1117_515;
  wire w_1118_533, w_1118_1455, w_1118_1456, w_1118_1457, w_1118_1458, w_1118_1459, w_1118_1460, w_1118_1461, w_1118_1462, w_1118_1463, w_1118_1464;
  wire w_1124_1428;
  wire w_1126_121;
  wire w_1128_466;
  wire w_1131_656, w_1131_664;
  wire w_1132_1117, w_1132_1118, w_1132_1119, w_1132_1120, w_1132_1121, w_1132_1122, w_1132_1123;
  wire w_1133_1692;
  wire w_1134_1163;
  wire w_1137_216;
  wire w_1139_1355;
  wire w_1142_154;
  wire w_1148_133;
  wire w_1157_360;
  wire w_1158_191;
  wire w_1161_784;
  wire w_1162_232;
  wire w_1165_045;
  wire w_1166_032;
  wire w_1168_039;
  wire w_1169_327;
  wire w_1173_1388;
  wire w_1176_1251, w_1176_1252, w_1176_1253, w_1176_1254, w_1176_1255, w_1176_1256, w_1176_1257, w_1176_1258, w_1176_1259, w_1176_1260, w_1176_1261, w_1176_1262;
  wire w_1178_104;
  wire w_1181_634, w_1181_769;
  wire w_1183_177;
  wire w_1190_258;
  wire w_1192_779;
  wire w_1194_032, w_1194_157;
  wire w_1199_581, w_1199_1954, w_1199_1955, w_1199_1956, w_1199_1960, w_1199_1961, w_1199_1962, w_1199_1963, w_1199_1964, w_1199_1965, w_1199_1966, w_1199_1967, w_1199_1968, w_1199_1969, w_1199_1970, w_1199_1971, w_1199_1973;
  wire w_1200_704;
  wire w_1203_345;
  wire w_1204_137;
  wire w_1208_1034;
  wire w_1209_041;
  wire w_1212_003, w_1212_232;
  wire w_1213_087, w_1213_239;
  wire w_1215_855;
  wire w_1224_1447;
  wire w_1226_737, w_1226_1459;
  wire w_1227_414;
  wire w_1230_965, w_1230_966, w_1230_967, w_1230_968, w_1230_969, w_1230_970;
  wire w_1231_107, w_1231_150;
  wire w_1235_950, w_1235_1006;
  wire w_1236_1603;
  wire w_1239_311, w_1239_502;
  wire w_1240_471;
  wire w_1244_049;
  wire w_1246_814;
  wire w_1252_023;
  wire w_1253_704, w_1253_710;
  wire w_1258_009, w_1258_040;
  wire w_1259_894;
  wire w_1267_451;
  wire w_1270_723;
  wire w_1274_815;
  wire w_1275_1432, w_1275_1433, w_1275_1434, w_1275_1435, w_1275_1436, w_1275_1437, w_1275_1438, w_1275_1439, w_1275_1440, w_1275_1444, w_1275_1445, w_1275_1446, w_1275_1447, w_1275_1448, w_1275_1449, w_1275_1450, w_1275_1451, w_1275_1452, w_1275_1453, w_1275_1454, w_1275_1456;
  wire w_1276_796;
  wire w_1281_436;
  wire w_1288_1602, w_1288_1603, w_1288_1604, w_1288_1605, w_1288_1606, w_1288_1607, w_1288_1611, w_1288_1612, w_1288_1613, w_1288_1614, w_1288_1615, w_1288_1616, w_1288_1617, w_1288_1618, w_1288_1619, w_1288_1620, w_1288_1622;
  wire w_1289_284, w_1289_456, w_1289_457, w_1289_458, w_1289_459, w_1289_460, w_1289_461, w_1289_462, w_1289_463;
  wire w_1293_1762;
  wire w_1297_202;
  wire w_1298_518, w_1298_519, w_1298_520, w_1298_524, w_1298_525, w_1298_526, w_1298_527, w_1298_529;
  wire w_1299_668;
  wire w_1301_098;
  wire w_1303_222;
  wire w_1304_708;
  wire w_1305_025, w_1305_036;
  wire w_1308_361, w_1308_362, w_1308_363, w_1308_364, w_1308_365, w_1308_366, w_1308_367, w_1308_368, w_1308_369, w_1308_370, w_1308_371, w_1308_372, w_1308_376, w_1308_377, w_1308_378, w_1308_379, w_1308_380, w_1308_381, w_1308_382, w_1308_384;
  wire w_1312_969, w_1312_970, w_1312_971, w_1312_972, w_1312_973, w_1312_974, w_1312_975, w_1312_976, w_1312_977, w_1312_978, w_1312_979, w_1312_980, w_1312_984, w_1312_985, w_1312_986, w_1312_988;
  wire w_1316_035;
  wire w_1320_000;
  wire w_1321_169;
  wire w_1329_047, w_1329_157, w_1329_196;
  wire w_1330_429;
  wire w_1331_343;
  wire w_1335_651;
  wire w_1339_1486;
  wire w_1354_916;
  wire w_1362_599;
  wire w_1363_168;
  wire w_1367_1256;
  wire w_1369_038;
  wire w_1375_1357;
  wire w_1376_518;
  wire w_1378_503;
  wire w_1380_542;
  wire w_1381_336;
  wire w_1391_245;
  wire w_1392_360;
  wire w_1395_110;
  wire w_1396_1004;
  wire w_1399_334;
  wire w_1400_522;
  wire w_1403_125;
  wire w_1410_066, w_1410_086;
  wire w_1422_540, w_1422_541, w_1422_542, w_1422_543, w_1422_544;
  wire w_1423_462, w_1423_463, w_1423_464, w_1423_465, w_1423_466, w_1423_467, w_1423_468, w_1423_469, w_1423_470, w_1423_471, w_1423_472;
  wire w_1427_403;
  wire w_1428_144;
  wire w_1429_723;
  wire w_1433_189;
  wire w_1440_698;
  wire w_1446_545;
  wire w_1449_388, w_1449_428, w_1449_506, w_1449_507, w_1449_508, w_1449_509;
  wire w_1454_158;
  wire w_1455_105;
  wire w_1463_378, w_1463_482;
  wire w_1468_475;
  wire w_1486_226;
  wire w_1492_357;
  wire w_1494_332;
  wire w_1496_083;
  wire w_1502_1051;
  wire w_1503_257;
  wire w_1505_029;
  wire w_1510_151;
  wire w_1511_527;
  wire w_1513_018;
  wire w_1524_069;
  wire w_1529_1173;
  wire w_1530_672;
  wire w_1534_349;
  wire w_1538_208;
  wire w_1539_021;
  wire w_1542_076;
  wire w_1549_655;
  wire w_1550_140;
  wire w_1560_137, w_1560_289;
  wire w_1561_166;
  wire w_1563_104;
  wire w_1577_015;
  wire w_1578_109;
  wire w_1579_1708, w_1579_1709, w_1579_1710, w_1579_1711, w_1579_1712, w_1579_1713, w_1579_1714, w_1579_1715;
  wire w_1580_224;
  wire w_1586_998, w_1586_1357;
  wire w_1589_1440;
  wire w_1590_840;
  wire w_1594_878;
  wire w_1596_216;
  wire w_1598_1875, w_1598_1876, w_1598_1877, w_1598_1878, w_1598_1879, w_1598_1880, w_1598_1881, w_1598_1882, w_1598_1883, w_1598_1884, w_1598_1885;
  wire w_1601_113, w_1601_114, w_1601_115, w_1601_119, w_1601_120, w_1601_121, w_1601_122, w_1601_123, w_1601_124, w_1601_125, w_1601_127;
  wire w_1603_907, w_1603_1223, w_1603_1583;
  wire w_1605_144;
  wire w_1609_218;
  wire w_1615_1009;
  wire w_1622_078;
  wire w_1629_026;
  wire w_1635_431;
  wire w_1652_404;
  wire w_1656_1927, w_1656_1928, w_1656_1929, w_1656_1930;
  wire w_1666_1997, w_1666_1998, w_1666_1999, w_1666_2000, w_1666_2001, w_1666_2002, w_1666_2003, w_1666_2004, w_1666_2005, w_1666_2006, w_1666_2007, w_1666_2008, w_1666_2012, w_1666_2013, w_1666_2014, w_1666_2016;
  wire w_1673_151;
  wire w_1687_828;
  wire w_1688_1681, w_1688_1682, w_1688_1683, w_1688_1684, w_1688_1685, w_1688_1686, w_1688_1687, w_1688_1688;
  wire w_1692_078, w_1692_766, w_1692_767, w_1692_768, w_1692_769, w_1692_770, w_1692_774, w_1692_775, w_1692_776, w_1692_777, w_1692_778, w_1692_779, w_1692_780, w_1692_782;
  wire w_1701_010;
  wire w_1716_1335;
  wire w_1721_407, w_1721_863;
  wire w_1726_437;
  wire w_1727_092;
  wire w_1732_311;
  wire w_1734_083;
  wire w_1754_1116;
  wire w_1755_243;
  wire w_1760_002, w_1760_054;
  wire w_1774_625;
  wire w_1777_499;
  wire w_1787_1409;
  wire w_1800_369;
  wire w_1801_026;
  wire w_1806_215;
  wire w_1810_274;
  wire w_1811_265;
  wire w_1816_144;
  wire w_1818_359, w_1818_360, w_1818_361, w_1818_362;
  wire w_1819_036;
  wire w_1820_561;
  wire w_1821_248, w_1821_249, w_1821_250, w_1821_251, w_1821_252, w_1821_253, w_1821_257, w_1821_258, w_1821_259, w_1821_260, w_1821_261, w_1821_262, w_1821_263, w_1821_264, w_1821_265, w_1821_266, w_1821_268;
  wire w_1824_1452, w_1824_1453, w_1824_1454;
  wire w_1833_629;
  wire w_1836_1757, w_1836_1758, w_1836_1759, w_1836_1760, w_1836_1761, w_1836_1762, w_1836_1763, w_1836_1764, w_1836_1765, w_1836_1766, w_1836_1767, w_1836_1768, w_1836_1772, w_1836_1773, w_1836_1774, w_1836_1775, w_1836_1776, w_1836_1778;
  wire w_1848_117, w_1848_118, w_1848_119, w_1848_120;
  wire w_1871_787;
  wire w_1873_820;
  wire w_1885_477;
  wire w_1890_797;
  wire w_1891_031;
  wire w_1904_1675;
  wire w_1905_377;
  wire w_1911_1096, w_1911_1097, w_1911_1098, w_1911_1099, w_1911_1100, w_1911_1101, w_1911_1102, w_1911_1103, w_1911_1104, w_1911_1105, w_1911_1106, w_1911_1107;
  wire w_1916_638;
  wire w_1927_525;
  wire w_1937_085;
  wire w_1940_595;
  wire w_1943_034;
  wire w_1964_004;
  wire w_1983_007;
  wire w_1986_071, w_1986_421;
  wire w_1990_1658;
  wire w_1994_186;
  wire w_1997_662;
  wire w_2000_000, w_2000_001, w_2000_002, w_2000_003, w_2000_004, w_2000_005, w_2000_006, w_2000_007, w_2000_008, w_2000_009, w_2000_010, w_2000_011, w_2000_012, w_2000_013, w_2000_014, w_2000_015, w_2000_016, w_2000_017, w_2000_018, w_2000_019, w_2000_020, w_2000_021, w_2000_022, w_2000_023, w_2000_024, w_2000_025, w_2000_026, w_2000_027, w_2000_028, w_2000_029, w_2000_030, w_2000_031, w_2000_032, w_2000_033, w_2000_034, w_2000_035, w_2000_036, w_2000_037, w_2000_038, w_2000_039, w_2000_040, w_2000_041, w_2000_042, w_2000_043, w_2000_044, w_2000_045, w_2000_046, w_2000_047, w_2000_048, w_2000_049, w_2000_050, w_2000_051, w_2000_052, w_2000_053, w_2000_054, w_2000_055, w_2000_056, w_2000_057, w_2000_058, w_2000_059, w_2000_060, w_2000_061, w_2000_062, w_2000_063, w_2000_064, w_2000_065, w_2000_066, w_2000_067, w_2000_068, w_2000_069, w_2000_070, w_2000_071, w_2000_072, w_2000_073, w_2000_074, w_2000_075, w_2000_076, w_2000_077, w_2000_078, w_2000_079, w_2000_080, w_2000_081, w_2000_082, w_2000_083, w_2000_084, w_2000_085, w_2000_086, w_2000_087, w_2000_088, w_2000_089, w_2000_090, w_2000_091, w_2000_092, w_2000_093, w_2000_094, w_2000_095, w_2000_096, w_2000_097, w_2000_098, w_2000_099, w_2000_100, w_2000_101, w_2000_102, w_2000_103, w_2000_104, w_2000_105, w_2000_106, w_2000_107, w_2000_108, w_2000_109, w_2000_110;
  not1 I001_000(w_001_000, w_000_000);
  nand2 I001_001(w_001_001, w_000_001, w_000_002);
  not1 I001_002(w_001_002, w_000_003);
  or2  I001_003(w_001_003, w_000_004, w_000_005);
  nand2 I001_004(w_001_004, w_000_006, w_000_007);
  nand2 I001_005(w_001_005, w_000_008, w_000_009);
  not1 I001_006(w_001_006, w_000_010);
  and2 I001_007(w_001_007, w_000_011, w_000_012);
  nand2 I001_008(w_001_008, w_000_013, w_000_014);
  not1 I001_009(w_001_009, w_000_015);
  nand2 I001_010(w_001_010, w_000_016, w_000_017);
  or2  I001_011(w_001_011, w_000_018, w_000_019);
  not1 I001_012(w_001_012, w_000_020);
  nand2 I001_013(w_001_013, w_000_021, w_000_022);
  nand2 I001_014(w_001_014, w_000_023, w_000_024);
  or2  I001_015(w_001_015, w_000_025, w_000_026);
  and2 I001_016(w_001_016, w_000_027, w_000_028);
  and2 I001_017(w_001_017, w_000_029, w_000_030);
  or2  I001_018(w_001_018, w_000_031, w_000_032);
  and2 I001_019(w_001_019, w_000_033, w_000_034);
  not1 I001_020(w_001_020, w_000_035);
  and2 I001_021(w_001_021, w_000_036, w_000_037);
  or2  I001_022(w_001_022, w_000_038, w_000_039);
  and2 I001_023(w_001_023, w_000_040, w_000_041);
  or2  I001_024(w_001_024, w_000_042, w_000_043);
  and2 I001_025(w_001_025, w_000_044, w_000_045);
  or2  I001_026(w_001_026, w_000_046, w_000_047);
  not1 I001_027(w_001_027, w_000_048);
  nand2 I001_028(w_001_028, w_000_049, w_000_050);
  and2 I001_029(w_001_029, w_000_051, w_000_052);
  and2 I001_030(w_001_030, w_000_053, w_000_054);
  nand2 I001_031(w_001_031, w_000_055, w_000_056);
  and2 I001_032(w_001_032, w_000_057, w_000_058);
  and2 I001_033(w_001_033, w_000_059, w_000_012);
  not1 I001_034(w_001_034, w_000_060);
  not1 I001_035(w_001_035, w_000_061);
  nand2 I001_036(w_001_036, w_000_062, w_000_063);
  or2  I001_038(w_001_038, w_000_065, w_000_066);
  or2  I001_039(w_001_039, w_000_067, w_000_068);
  and2 I001_040(w_001_040, w_000_069, w_000_070);
  not1 I001_041(w_001_041, w_000_071);
  or2  I001_042(w_001_042, w_000_072, w_000_073);
  nand2 I001_043(w_001_043, w_000_074, w_000_075);
  nand2 I001_044(w_001_044, w_000_076, w_000_077);
  nand2 I001_045(w_001_045, w_000_078, w_000_079);
  or2  I001_046(w_001_046, w_000_080, w_000_081);
  and2 I001_047(w_001_047, w_000_082, w_000_083);
  not1 I001_048(w_001_048, w_000_084);
  not1 I001_049(w_001_049, w_000_085);
  nand2 I001_050(w_001_050, w_000_086, w_000_087);
  nand2 I001_051(w_001_051, w_000_088, w_000_089);
  nand2 I001_052(w_001_052, w_000_019, w_000_090);
  and2 I001_053(w_001_053, w_000_091, w_000_092);
  and2 I001_054(w_001_054, w_000_093, w_000_094);
  nand2 I001_055(w_001_055, w_000_095, w_000_096);
  not1 I001_056(w_001_056, w_000_097);
  or2  I001_057(w_001_057, w_000_098, w_000_099);
  or2  I001_059(w_001_059, w_000_102, w_000_103);
  and2 I001_060(w_001_060, w_000_104, w_000_105);
  and2 I001_061(w_001_061, w_000_106, w_000_107);
  and2 I001_062(w_001_062, w_000_108, w_000_109);
  nand2 I001_063(w_001_063, w_000_110, w_000_111);
  and2 I001_064(w_001_064, w_000_112, w_000_113);
  or2  I001_065(w_001_065, w_000_114, w_000_115);
  nand2 I001_066(w_001_066, w_000_116, w_000_117);
  not1 I001_067(w_001_067, w_000_118);
  or2  I001_068(w_001_068, w_000_119, w_000_120);
  or2  I001_069(w_001_069, w_000_121, w_000_122);
  nand2 I001_070(w_001_070, w_000_123, w_000_124);
  or2  I001_071(w_001_071, w_000_125, w_000_126);
  nand2 I001_072(w_001_072, w_000_127, w_000_128);
  not1 I001_073(w_001_073, w_000_129);
  and2 I001_074(w_001_074, w_000_130, w_000_131);
  and2 I001_075(w_001_075, w_000_132, w_000_133);
  or2  I001_076(w_001_076, w_000_134, w_000_135);
  and2 I001_077(w_001_077, w_000_136, w_000_137);
  nand2 I001_078(w_001_078, w_000_138, w_000_139);
  and2 I001_079(w_001_079, w_000_140, w_000_141);
  not1 I001_080(w_001_080, w_000_142);
  nand2 I001_081(w_001_081, w_000_143, w_000_144);
  or2  I001_082(w_001_082, w_000_082, w_000_145);
  and2 I001_083(w_001_083, w_000_146, w_000_147);
  nand2 I001_084(w_001_084, w_000_148, w_000_149);
  nand2 I001_086(w_001_086, w_000_152, w_000_153);
  and2 I001_087(w_001_087, w_000_154, w_000_155);
  nand2 I001_088(w_001_088, w_000_156, w_000_157);
  not1 I001_090(w_001_090, w_000_160);
  and2 I001_091(w_001_091, w_000_161, w_000_162);
  not1 I001_092(w_001_092, w_000_163);
  or2  I001_093(w_001_093, w_000_164, w_000_165);
  not1 I001_094(w_001_094, w_000_166);
  and2 I001_095(w_001_095, w_000_167, w_000_062);
  and2 I001_096(w_001_096, w_000_168, w_000_036);
  and2 I001_097(w_001_097, w_000_169, w_000_170);
  not1 I001_098(w_001_098, w_000_171);
  nand2 I001_099(w_001_099, w_000_172, w_000_173);
  or2  I001_100(w_001_100, w_000_174, w_000_175);
  not1 I001_101(w_001_101, w_000_176);
  nand2 I001_102(w_001_102, w_000_177, w_000_178);
  nand2 I001_103(w_001_103, w_000_179, w_000_180);
  or2  I001_104(w_001_104, w_000_181, w_000_182);
  not1 I001_106(w_001_106, w_000_184);
  and2 I001_107(w_001_107, w_000_185, w_000_090);
  and2 I001_108(w_001_108, w_000_186, w_000_187);
  and2 I001_109(w_001_109, w_000_188, w_000_189);
  and2 I001_110(w_001_110, w_000_190, w_000_191);
  nand2 I001_111(w_001_111, w_000_192, w_000_193);
  and2 I001_112(w_001_112, w_000_194, w_000_009);
  and2 I001_113(w_001_113, w_000_195, w_000_196);
  nand2 I001_114(w_001_114, w_000_197, w_000_198);
  or2  I001_115(w_001_115, w_000_199, w_000_200);
  nand2 I001_116(w_001_116, w_000_201, w_000_202);
  or2  I001_117(w_001_117, w_000_203, w_000_204);
  or2  I001_119(w_001_119, w_000_207, w_000_208);
  not1 I001_120(w_001_120, w_000_209);
  not1 I001_121(w_001_121, w_000_210);
  and2 I001_122(w_001_122, w_000_211, w_000_212);
  and2 I001_123(w_001_123, w_000_081, w_000_213);
  and2 I001_124(w_001_124, w_000_214, w_000_215);
  and2 I001_125(w_001_125, w_000_216, w_000_217);
  or2  I001_126(w_001_126, w_000_218, w_000_219);
  and2 I001_127(w_001_127, w_000_042, w_000_220);
  or2  I001_128(w_001_128, w_000_221, w_000_190);
  and2 I001_129(w_001_129, w_000_222, w_000_209);
  or2  I001_130(w_001_130, w_000_223, w_000_224);
  and2 I001_131(w_001_131, w_000_225, w_000_226);
  and2 I001_132(w_001_132, w_000_227, w_000_228);
  or2  I001_133(w_001_133, w_000_229, w_000_230);
  nand2 I001_134(w_001_134, w_000_231, w_000_142);
  nand2 I001_135(w_001_135, w_000_232, w_000_233);
  and2 I001_137(w_001_137, w_000_236, w_000_237);
  not1 I001_138(w_001_138, w_000_238);
  nand2 I001_139(w_001_139, w_000_239, w_000_202);
  not1 I001_140(w_001_140, w_000_240);
  and2 I001_141(w_001_141, w_000_021, w_000_241);
  and2 I001_142(w_001_142, w_000_242, w_000_243);
  and2 I001_143(w_001_143, w_000_244, w_000_245);
  and2 I001_145(w_001_145, w_000_246, w_000_247);
  and2 I001_147(w_001_147, w_000_249, w_000_250);
  nand2 I001_148(w_001_148, w_000_251, w_000_252);
  or2  I001_149(w_001_149, w_000_253, w_000_046);
  and2 I001_150(w_001_150, w_000_254, w_000_249);
  not1 I001_151(w_001_151, w_000_255);
  or2  I001_152(w_001_152, w_000_256, w_000_257);
  or2  I001_153(w_001_153, w_000_258, w_000_259);
  or2  I001_154(w_001_154, w_000_260, w_000_261);
  nand2 I001_155(w_001_155, w_000_262, w_000_263);
  or2  I001_156(w_001_156, w_000_264, w_000_265);
  not1 I001_157(w_001_157, w_000_266);
  nand2 I001_159(w_001_159, w_000_050, w_000_268);
  and2 I001_160(w_001_160, w_000_269, w_000_270);
  or2  I001_161(w_001_161, w_000_271, w_000_272);
  nand2 I001_162(w_001_162, w_000_002, w_000_273);
  nand2 I001_163(w_001_163, w_000_274, w_000_275);
  nand2 I001_164(w_001_164, w_000_276, w_000_159);
  nand2 I001_165(w_001_165, w_000_277, w_000_134);
  nand2 I001_166(w_001_166, w_000_278, w_000_215);
  or2  I001_168(w_001_168, w_000_281, w_000_282);
  or2  I001_169(w_001_169, w_000_283, w_000_284);
  or2  I001_170(w_001_170, w_000_285, w_000_286);
  nand2 I001_172(w_001_172, w_000_289, w_000_290);
  nand2 I001_173(w_001_173, w_000_291, w_000_292);
  or2  I001_174(w_001_174, w_000_293, w_000_294);
  and2 I001_175(w_001_175, w_000_295, w_000_296);
  not1 I001_176(w_001_176, w_000_232);
  or2  I001_177(w_001_177, w_000_042, w_000_297);
  or2  I001_178(w_001_178, w_000_023, w_000_298);
  or2  I001_179(w_001_179, w_000_299, w_000_300);
  or2  I001_180(w_001_180, w_000_301, w_000_302);
  or2  I001_181(w_001_181, w_000_234, w_000_303);
  not1 I001_182(w_001_182, w_000_304);
  or2  I001_183(w_001_183, w_000_305, w_000_306);
  or2  I001_184(w_001_184, w_000_307, w_000_308);
  not1 I001_185(w_001_185, w_000_309);
  not1 I001_186(w_001_186, w_000_310);
  not1 I001_187(w_001_187, w_000_311);
  and2 I001_188(w_001_188, w_000_312, w_000_313);
  not1 I001_189(w_001_189, w_000_290);
  nand2 I001_190(w_001_190, w_000_314, w_000_315);
  and2 I001_191(w_001_191, w_000_316, w_000_317);
  or2  I001_192(w_001_192, w_000_318, w_000_319);
  not1 I001_193(w_001_193, w_000_320);
  nand2 I001_194(w_001_194, w_000_321, w_000_090);
  and2 I001_195(w_001_195, w_000_322, w_000_323);
  or2  I001_196(w_001_196, w_000_189, w_000_274);
  nand2 I001_197(w_001_197, w_000_324, w_000_325);
  or2  I001_198(w_001_198, w_000_326, w_000_327);
  not1 I001_199(w_001_199, w_000_328);
  not1 I001_200(w_001_200, w_000_329);
  and2 I001_201(w_001_201, w_000_330, w_000_331);
  and2 I001_202(w_001_202, w_000_332, w_000_237);
  or2  I001_203(w_001_203, w_000_333, w_000_334);
  not1 I001_204(w_001_204, w_000_335);
  nand2 I001_205(w_001_205, w_000_336, w_000_337);
  or2  I001_206(w_001_206, w_000_338, w_000_289);
  nand2 I001_207(w_001_207, w_000_339, w_000_340);
  or2  I001_208(w_001_208, w_000_341, w_000_342);
  or2  I001_209(w_001_209, w_000_343, w_000_344);
  not1 I001_210(w_001_210, w_000_345);
  or2  I001_212(w_001_212, w_000_157, w_000_348);
  or2  I001_213(w_001_213, w_000_349, w_000_270);
  nand2 I001_214(w_001_214, w_000_350, w_000_351);
  not1 I001_216(w_001_216, w_000_354);
  nand2 I001_217(w_001_217, w_000_355, w_000_356);
  not1 I001_218(w_001_218, w_000_357);
  and2 I001_219(w_001_219, w_000_358, w_000_359);
  not1 I001_221(w_001_221, w_000_361);
  or2  I001_223(w_001_223, w_000_364, w_000_365);
  not1 I001_224(w_001_224, w_000_030);
  not1 I001_225(w_001_225, w_000_366);
  or2  I001_226(w_001_226, w_000_367, w_000_368);
  not1 I001_227(w_001_227, w_000_231);
  nand2 I001_228(w_001_228, w_000_369, w_000_370);
  not1 I001_229(w_001_229, w_000_371);
  not1 I001_230(w_001_230, w_000_372);
  not1 I001_231(w_001_231, w_000_373);
  and2 I001_232(w_001_232, w_000_374, w_000_375);
  or2  I001_233(w_001_233, w_000_376, w_000_377);
  and2 I001_234(w_001_234, w_000_378, w_000_379);
  nand2 I001_235(w_001_235, w_000_380, w_000_381);
  nand2 I001_236(w_001_236, w_000_382, w_000_127);
  not1 I001_237(w_001_237, w_000_383);
  and2 I001_238(w_001_238, w_000_384, w_000_385);
  nand2 I001_239(w_001_239, w_000_049, w_000_386);
  nand2 I001_240(w_001_240, w_000_387, w_000_388);
  nand2 I001_241(w_001_241, w_000_389, w_000_390);
  not1 I001_242(w_001_242, w_000_391);
  and2 I001_243(w_001_243, w_000_392, w_000_393);
  or2  I001_244(w_001_244, w_000_394, w_000_395);
  not1 I001_245(w_001_245, w_000_396);
  not1 I001_246(w_001_246, w_000_397);
  not1 I001_247(w_001_247, w_000_126);
  or2  I001_248(w_001_248, w_000_398, w_000_253);
  nand2 I001_249(w_001_249, w_000_399, w_000_400);
  or2  I001_250(w_001_250, w_000_179, w_000_377);
  not1 I001_251(w_001_251, w_000_401);
  and2 I001_252(w_001_252, w_000_402, w_000_403);
  and2 I001_253(w_001_253, w_000_294, w_000_404);
  not1 I001_254(w_001_254, w_000_235);
  or2  I001_255(w_001_255, w_000_405, w_000_406);
  nand2 I001_256(w_001_256, w_000_407, w_000_328);
  or2  I001_257(w_001_257, w_000_408, w_000_409);
  not1 I001_258(w_001_258, w_000_410);
  and2 I001_259(w_001_259, w_000_411, w_000_412);
  not1 I001_260(w_001_260, w_000_413);
  not1 I001_261(w_001_261, w_000_414);
  nand2 I001_262(w_001_262, w_000_415, w_000_416);
  or2  I001_263(w_001_263, w_000_417, w_000_418);
  and2 I001_264(w_001_264, w_000_419, w_000_420);
  not1 I001_265(w_001_265, w_000_421);
  nand2 I001_266(w_001_266, w_000_422, w_000_423);
  nand2 I001_267(w_001_267, w_000_424, w_000_425);
  and2 I001_268(w_001_268, w_000_426, w_000_226);
  nand2 I001_269(w_001_269, w_000_427, w_000_428);
  or2  I001_270(w_001_270, w_000_429, w_000_430);
  and2 I001_271(w_001_271, w_000_431, w_000_432);
  not1 I001_272(w_001_272, w_000_433);
  not1 I001_273(w_001_273, w_000_434);
  and2 I001_274(w_001_274, w_000_379, w_000_435);
  not1 I001_275(w_001_275, w_000_436);
  and2 I001_276(w_001_276, w_000_427, w_000_234);
  not1 I001_278(w_001_278, w_000_438);
  nand2 I001_279(w_001_279, w_000_347, w_000_439);
  not1 I001_280(w_001_280, w_000_440);
  not1 I001_281(w_001_281, w_000_059);
  not1 I001_282(w_001_282, w_000_047);
  and2 I001_283(w_001_283, w_000_441, w_000_442);
  and2 I001_284(w_001_284, w_000_443, w_000_444);
  nand2 I001_285(w_001_285, w_000_445, w_000_446);
  and2 I001_286(w_001_286, w_000_278, w_000_447);
  not1 I001_287(w_001_287, w_000_448);
  nand2 I001_288(w_001_288, w_000_449, w_000_450);
  nand2 I001_289(w_001_289, w_000_324, w_000_272);
  not1 I001_290(w_001_290, w_000_154);
  nand2 I001_291(w_001_291, w_000_451, w_000_452);
  or2  I001_292(w_001_292, w_000_453, w_000_454);
  and2 I001_293(w_001_293, w_000_269, w_000_455);
  or2  I001_294(w_001_294, w_000_456, w_000_457);
  or2  I001_295(w_001_295, w_000_458, w_000_459);
  and2 I001_296(w_001_296, w_000_460, w_000_461);
  and2 I001_297(w_001_297, w_000_462, w_000_463);
  not1 I001_298(w_001_298, w_000_464);
  nand2 I001_299(w_001_299, w_000_376, w_000_465);
  nand2 I001_300(w_001_300, w_000_466, w_000_467);
  not1 I001_302(w_001_302, w_000_470);
  and2 I001_303(w_001_303, w_000_471, w_000_472);
  or2  I001_305(w_001_305, w_000_474, w_000_475);
  not1 I001_306(w_001_306, w_000_476);
  not1 I001_307(w_001_307, w_000_067);
  nand2 I001_308(w_001_308, w_000_477, w_000_478);
  nand2 I001_309(w_001_309, w_000_479, w_000_122);
  or2  I001_310(w_001_310, w_000_480, w_000_481);
  nand2 I001_311(w_001_311, w_000_482, w_000_254);
  not1 I001_312(w_001_312, w_000_483);
  or2  I001_313(w_001_313, w_000_484, w_000_485);
  or2  I001_316(w_001_316, w_000_488, w_000_489);
  and2 I001_317(w_001_317, w_000_490, w_000_491);
  nand2 I001_319(w_001_319, w_000_297, w_000_032);
  not1 I001_321(w_001_321, w_000_415);
  or2  I001_322(w_001_322, w_000_494, w_000_495);
  nand2 I001_323(w_001_323, w_000_496, w_000_297);
  or2  I001_325(w_001_325, w_000_498, w_000_499);
  and2 I001_326(w_001_326, w_000_500, w_000_501);
  or2  I001_329(w_001_329, w_000_505, w_000_285);
  not1 I001_330(w_001_330, w_000_506);
  nand2 I001_331(w_001_331, w_000_507, w_000_508);
  and2 I001_335(w_001_335, w_000_515, w_000_516);
  or2  I001_336(w_001_336, w_000_517, w_000_518);
  or2  I001_337(w_001_337, w_000_310, w_000_519);
  and2 I001_338(w_001_338, w_000_225, w_000_520);
  or2  I001_340(w_001_340, w_000_008, w_000_522);
  nand2 I001_341(w_001_341, w_000_350, w_000_523);
  or2  I001_342(w_001_342, w_000_524, w_000_525);
  or2  I001_343(w_001_343, w_000_071, w_000_526);
  or2  I001_344(w_001_344, w_000_527, w_000_528);
  nand2 I001_345(w_001_345, w_000_398, w_000_529);
  not1 I001_346(w_001_346, w_000_393);
  nand2 I001_348(w_001_348, w_000_532, w_000_533);
  nand2 I001_349(w_001_349, w_000_534, w_000_099);
  or2  I001_350(w_001_350, w_000_535, w_000_536);
  and2 I001_352(w_001_352, w_000_539, w_000_184);
  not1 I001_354(w_001_354, w_000_542);
  or2  I001_357(w_001_357, w_000_545, w_000_546);
  not1 I001_358(w_001_358, w_000_445);
  and2 I001_359(w_001_359, w_000_325, w_000_547);
  or2  I001_362(w_001_362, w_000_549, w_000_439);
  not1 I001_363(w_001_363, w_000_421);
  nand2 I001_364(w_001_364, w_000_550, w_000_551);
  not1 I001_365(w_001_365, w_000_552);
  not1 I001_366(w_001_366, w_000_553);
  or2  I001_367(w_001_367, w_000_554, w_000_555);
  or2  I001_370(w_001_370, w_000_557, w_000_558);
  nand2 I001_371(w_001_371, w_000_506, w_000_559);
  and2 I001_372(w_001_372, w_000_560, w_000_263);
  nand2 I001_373(w_001_373, w_000_561, w_000_037);
  or2  I001_374(w_001_374, w_000_562, w_000_563);
  not1 I001_377(w_001_377, w_000_567);
  or2  I001_378(w_001_378, w_000_568, w_000_569);
  or2  I001_379(w_001_379, w_000_570, w_000_571);
  nand2 I001_384(w_001_384, w_000_576, w_000_141);
  and2 I001_386(w_001_386, w_000_170, w_000_578);
  and2 I001_387(w_001_387, w_000_579, w_000_580);
  not1 I001_388(w_001_388, w_000_465);
  not1 I001_389(w_001_389, w_000_326);
  not1 I001_390(w_001_390, w_000_183);
  nand2 I001_391(w_001_391, w_000_581, w_000_582);
  and2 I001_392(w_001_392, w_000_583, w_000_393);
  not1 I001_393(w_001_393, w_000_584);
  or2  I001_394(w_001_394, w_000_585, w_000_586);
  and2 I001_395(w_001_395, w_000_587, w_000_548);
  or2  I001_397(w_001_397, w_000_589, w_000_590);
  nand2 I001_398(w_001_398, w_000_591, w_000_592);
  and2 I001_399(w_001_399, w_000_156, w_000_593);
  or2  I001_400(w_001_400, w_000_594, w_000_595);
  nand2 I001_401(w_001_401, w_000_596, w_000_597);
  not1 I001_404(w_001_404, w_000_100);
  not1 I001_405(w_001_405, w_000_600);
  and2 I001_406(w_001_406, w_000_042, w_000_601);
  nand2 I001_407(w_001_407, w_000_602, w_000_289);
  and2 I001_408(w_001_408, w_000_603, w_000_604);
  nand2 I001_409(w_001_409, w_000_605, w_000_606);
  and2 I001_411(w_001_411, w_000_608, w_000_609);
  nand2 I001_412(w_001_412, w_000_610, w_000_011);
  nand2 I001_413(w_001_413, w_000_611, w_000_192);
  or2  I001_414(w_001_414, w_000_612, w_000_613);
  nand2 I001_416(w_001_416, w_000_616, w_000_617);
  nand2 I001_417(w_001_417, w_000_377, w_000_618);
  and2 I001_418(w_001_418, w_000_573, w_000_619);
  not1 I001_419(w_001_419, w_000_125);
  or2  I001_420(w_001_420, w_000_620, w_000_496);
  not1 I001_421(w_001_421, w_000_621);
  or2  I001_422(w_001_422, w_000_622, w_000_623);
  and2 I001_423(w_001_423, w_000_624, w_000_625);
  and2 I001_424(w_001_424, w_000_305, w_000_030);
  or2  I001_425(w_001_425, w_000_626, w_000_627);
  and2 I001_426(w_001_426, w_000_562, w_000_424);
  nand2 I001_427(w_001_427, w_000_280, w_000_628);
  not1 I001_428(w_001_428, w_000_629);
  and2 I001_429(w_001_429, w_000_630, w_000_631);
  or2  I001_430(w_001_430, w_000_140, w_000_632);
  nand2 I001_431(w_001_431, w_000_633, w_000_557);
  or2  I001_432(w_001_432, w_000_431, w_000_634);
  not1 I001_435(w_001_435, w_000_639);
  nand2 I001_436(w_001_436, w_000_640, w_000_641);
  nand2 I001_438(w_001_438, w_000_644, w_000_645);
  or2  I001_440(w_001_440, w_000_232, w_000_646);
  not1 I001_442(w_001_442, w_000_433);
  nand2 I001_443(w_001_443, w_000_587, w_000_647);
  not1 I001_444(w_001_444, w_000_648);
  nand2 I001_445(w_001_445, w_000_351, w_000_649);
  and2 I001_446(w_001_446, w_000_650, w_000_651);
  not1 I001_447(w_001_447, w_000_652);
  or2  I001_448(w_001_448, w_000_653, w_000_186);
  or2  I001_449(w_001_449, w_000_654, w_000_655);
  nand2 I001_451(w_001_451, w_000_657, w_000_658);
  nand2 I001_452(w_001_452, w_000_659, w_000_660);
  and2 I001_453(w_001_453, w_000_661, w_000_139);
  nand2 I001_454(w_001_454, w_000_063, w_000_662);
  or2  I001_455(w_001_455, w_000_663, w_000_664);
  nand2 I001_457(w_001_457, w_000_667, w_000_668);
  nand2 I001_458(w_001_458, w_000_435, w_000_669);
  or2  I001_459(w_001_459, w_000_669, w_000_450);
  nand2 I001_460(w_001_460, w_000_670, w_000_671);
  not1 I001_461(w_001_461, w_000_089);
  not1 I001_466(w_001_466, w_000_679);
  nand2 I001_467(w_001_467, w_000_579, w_000_680);
  nand2 I001_470(w_001_470, w_000_683, w_000_684);
  or2  I001_471(w_001_471, w_000_685, w_000_353);
  not1 I001_472(w_001_472, w_000_686);
  not1 I001_473(w_001_473, w_000_687);
  not1 I001_474(w_001_474, w_000_688);
  and2 I001_475(w_001_475, w_000_689, w_000_690);
  or2  I001_476(w_001_476, w_000_691, w_000_480);
  not1 I001_478(w_001_478, w_000_123);
  or2  I001_479(w_001_479, w_000_693, w_000_694);
  or2  I001_480(w_001_480, w_000_312, w_000_695);
  or2  I001_481(w_001_481, w_000_696, w_000_697);
  and2 I001_482(w_001_482, w_000_698, w_000_699);
  nand2 I001_484(w_001_484, w_000_295, w_000_569);
  nand2 I001_485(w_001_485, w_000_702, w_000_703);
  and2 I001_486(w_001_486, w_000_571, w_000_704);
  or2  I001_487(w_001_487, w_000_705, w_000_172);
  nand2 I001_488(w_001_488, w_000_089, w_000_527);
  not1 I001_489(w_001_489, w_000_706);
  and2 I001_491(w_001_491, w_000_709, w_000_213);
  not1 I001_492(w_001_492, w_000_499);
  not1 I001_493(w_001_493, w_000_710);
  and2 I001_494(w_001_494, w_000_711, w_000_141);
  not1 I001_495(w_001_495, w_000_639);
  or2  I001_496(w_001_496, w_000_263, w_000_712);
  not1 I001_498(w_001_498, w_000_513);
  nand2 I001_499(w_001_499, w_000_714, w_000_257);
  nand2 I001_501(w_001_501, w_000_138, w_000_715);
  nand2 I001_502(w_001_502, w_000_716, w_000_421);
  and2 I001_503(w_001_503, w_000_717, w_000_634);
  not1 I001_504(w_001_504, w_000_718);
  and2 I001_505(w_001_505, w_000_719, w_000_720);
  and2 I001_506(w_001_506, w_000_721, w_000_722);
  nand2 I001_507(w_001_507, w_000_723, w_000_724);
  and2 I001_509(w_001_509, w_000_339, w_000_727);
  and2 I001_510(w_001_510, w_000_596, w_000_728);
  nand2 I001_511(w_001_511, w_000_729, w_000_013);
  or2  I001_512(w_001_512, w_000_519, w_000_730);
  not1 I001_513(w_001_513, w_000_731);
  and2 I001_514(w_001_514, w_000_732, w_000_279);
  nand2 I001_517(w_001_517, w_000_736, w_000_737);
  not1 I001_518(w_001_518, w_000_738);
  and2 I001_519(w_001_519, w_000_584, w_000_739);
  nand2 I001_520(w_001_520, w_000_740, w_000_741);
  or2  I001_521(w_001_521, w_000_496, w_000_440);
  nand2 I001_522(w_001_522, w_000_742, w_000_743);
  and2 I001_524(w_001_524, w_000_523, w_000_251);
  or2  I001_525(w_001_525, w_000_745, w_000_530);
  nand2 I001_526(w_001_526, w_000_704, w_000_746);
  not1 I001_527(w_001_527, w_000_302);
  or2  I001_528(w_001_528, w_000_747, w_000_748);
  nand2 I001_529(w_001_529, w_000_407, w_000_484);
  nand2 I001_530(w_001_530, w_000_749, w_000_750);
  nand2 I001_531(w_001_531, w_000_751, w_000_528);
  nand2 I001_532(w_001_532, w_000_752, w_000_753);
  nand2 I001_533(w_001_533, w_000_754, w_000_755);
  nand2 I001_535(w_001_535, w_000_438, w_000_757);
  and2 I001_537(w_001_537, w_000_098, w_000_486);
  not1 I001_538(w_001_538, w_000_752);
  nand2 I001_539(w_001_539, w_000_098, w_000_695);
  not1 I001_542(w_001_542, w_000_425);
  and2 I001_543(w_001_543, w_000_759, w_000_760);
  not1 I001_544(w_001_544, w_000_761);
  and2 I001_545(w_001_545, w_000_547, w_000_272);
  and2 I001_546(w_001_546, w_000_762, w_000_763);
  or2  I001_548(w_001_548, w_000_766, w_000_767);
  nand2 I001_549(w_001_549, w_000_035, w_000_768);
  nand2 I001_550(w_001_550, w_000_498, w_000_049);
  nand2 I001_553(w_001_553, w_000_770, w_000_771);
  and2 I001_554(w_001_554, w_000_772, w_000_773);
  or2  I001_555(w_001_555, w_000_115, w_000_560);
  or2  I001_556(w_001_556, w_000_774, w_000_775);
  and2 I001_558(w_001_558, w_000_329, w_000_777);
  or2  I001_559(w_001_559, w_000_778, w_000_634);
  and2 I001_560(w_001_560, w_000_779, w_000_585);
  nand2 I001_561(w_001_561, w_000_765, w_000_780);
  not1 I001_562(w_001_562, w_000_626);
  or2  I001_564(w_001_564, w_000_781, w_000_782);
  not1 I001_565(w_001_565, w_000_783);
  nand2 I001_566(w_001_566, w_000_784, w_000_428);
  and2 I001_567(w_001_567, w_000_785, w_000_786);
  not1 I001_568(w_001_568, w_000_300);
  not1 I001_569(w_001_569, w_000_787);
  or2  I001_570(w_001_570, w_000_763, w_000_788);
  and2 I001_571(w_001_571, w_000_789, w_000_790);
  nand2 I001_572(w_001_572, w_000_791, w_000_544);
  and2 I001_573(w_001_573, w_000_792, w_000_793);
  not1 I001_574(w_001_574, w_000_794);
  not1 I001_575(w_001_575, w_000_795);
  not1 I001_576(w_001_576, w_000_796);
  and2 I001_577(w_001_577, w_000_797, w_000_798);
  not1 I001_580(w_001_580, w_000_801);
  not1 I001_583(w_001_583, w_000_465);
  nand2 I001_584(w_001_584, w_000_804, w_000_805);
  nand2 I001_585(w_001_585, w_000_806, w_000_187);
  or2  I001_586(w_001_586, w_000_602, w_000_807);
  and2 I001_587(w_001_587, w_000_088, w_000_808);
  and2 I001_589(w_001_589, w_000_628, w_000_811);
  and2 I001_590(w_001_590, w_000_812, w_000_813);
  nand2 I001_592(w_001_592, w_000_815, w_000_816);
  and2 I001_593(w_001_593, w_000_515, w_000_487);
  not1 I001_594(w_001_594, w_000_817);
  not1 I001_595(w_001_595, w_000_818);
  or2  I001_596(w_001_596, w_000_819, w_000_820);
  and2 I001_597(w_001_597, w_000_821, w_000_293);
  nand2 I001_601(w_001_601, w_000_824, w_000_811);
  or2  I001_602(w_001_602, w_000_825, w_000_681);
  or2  I001_603(w_001_603, w_000_826, w_000_499);
  or2  I001_604(w_001_604, w_000_535, w_000_827);
  and2 I001_605(w_001_605, w_000_769, w_000_346);
  nand2 I001_606(w_001_606, w_000_828, w_000_829);
  or2  I001_609(w_001_609, w_000_832, w_000_833);
  and2 I001_610(w_001_610, w_000_114, w_000_371);
  not1 I001_612(w_001_612, w_000_835);
  and2 I001_613(w_001_613, w_000_836, w_000_697);
  and2 I001_614(w_001_614, w_000_067, w_000_837);
  nand2 I001_615(w_001_615, w_000_838, w_000_839);
  or2  I001_617(w_001_617, w_000_841, w_000_842);
  and2 I001_618(w_001_618, w_000_147, w_000_843);
  or2  I001_619(w_001_619, w_000_335, w_000_422);
  and2 I001_620(w_001_620, w_000_844, w_000_845);
  nand2 I001_621(w_001_621, w_000_339, w_000_766);
  or2  I001_622(w_001_622, w_000_846, w_000_847);
  and2 I001_623(w_001_623, w_000_848, w_000_849);
  or2  I001_624(w_001_624, w_000_850, w_000_851);
  nand2 I001_625(w_001_625, w_000_852, w_000_721);
  not1 I001_626(w_001_626, w_000_853);
  or2  I001_627(w_001_627, w_000_854, w_000_855);
  and2 I001_628(w_001_628, w_000_856, w_000_857);
  nand2 I001_629(w_001_629, w_000_798, w_000_858);
  nand2 I001_630(w_001_630, w_000_859, w_000_860);
  nand2 I001_631(w_001_631, w_000_616, w_000_267);
  nand2 I001_632(w_001_632, w_000_861, w_000_292);
  and2 I001_635(w_001_635, w_000_864, w_000_865);
  and2 I001_636(w_001_636, w_000_866, w_000_376);
  or2  I001_637(w_001_637, w_000_173, w_000_867);
  nand2 I001_638(w_001_638, w_000_868, w_000_673);
  or2  I001_639(w_001_639, w_000_481, w_000_869);
  or2  I001_640(w_001_640, w_000_396, w_000_870);
  not1 I001_641(w_001_641, w_000_280);
  nand2 I001_643(w_001_643, w_000_854, w_000_366);
  not1 I001_644(w_001_644, w_000_871);
  or2  I001_646(w_001_646, w_000_874, w_000_875);
  nand2 I001_649(w_001_649, w_000_879, w_000_880);
  and2 I001_650(w_001_650, w_000_071, w_000_881);
  nand2 I001_651(w_001_651, w_000_000, w_000_320);
  and2 I001_652(w_001_652, w_000_882, w_000_883);
  and2 I001_653(w_001_653, w_000_504, w_000_884);
  not1 I001_655(w_001_655, w_000_886);
  not1 I001_656(w_001_656, w_000_636);
  not1 I001_657(w_001_657, w_000_887);
  not1 I001_658(w_001_658, w_000_614);
  or2  I001_659(w_001_659, w_000_888, w_000_865);
  and2 I001_660(w_001_660, w_000_889, w_000_620);
  or2  I001_661(w_001_661, w_000_863, w_000_890);
  and2 I001_662(w_001_662, w_000_786, w_000_004);
  or2  I001_663(w_001_663, w_000_891, w_000_356);
  nand2 I001_665(w_001_665, w_000_569, w_000_128);
  or2  I001_666(w_001_666, w_000_892, w_000_893);
  not1 I001_667(w_001_667, w_000_894);
  not1 I001_668(w_001_668, w_000_895);
  or2  I001_669(w_001_669, w_000_896, w_000_897);
  and2 I001_671(w_001_671, w_000_238, w_000_699);
  or2  I001_672(w_001_672, w_000_000, w_000_899);
  or2  I001_673(w_001_673, w_000_900, w_000_348);
  or2  I001_674(w_001_674, w_000_017, w_000_901);
  nand2 I001_677(w_001_677, w_000_903, w_000_904);
  or2  I001_678(w_001_678, w_000_392, w_000_905);
  and2 I001_681(w_001_681, w_000_550, w_000_908);
  not1 I001_683(w_001_683, w_000_910);
  or2  I001_685(w_001_685, w_000_911, w_000_461);
  not1 I001_686(w_001_686, w_000_142);
  not1 I001_687(w_001_687, w_000_191);
  nand2 I001_688(w_001_688, w_000_912, w_000_913);
  not1 I001_689(w_001_689, w_000_538);
  not1 I001_691(w_001_691, w_000_422);
  not1 I001_692(w_001_692, w_000_915);
  nand2 I001_696(w_001_696, w_000_918, w_000_157);
  nand2 I001_697(w_001_697, w_000_602, w_000_492);
  and2 I001_698(w_001_698, w_000_296, w_000_919);
  not1 I001_699(w_001_699, w_000_840);
  or2  I001_700(w_001_700, w_000_920, w_000_512);
  and2 I001_701(w_001_701, w_000_921, w_000_922);
  and2 I001_702(w_001_702, w_000_872, w_000_428);
  and2 I001_704(w_001_704, w_000_576, w_000_337);
  not1 I001_707(w_001_707, w_000_782);
  not1 I001_708(w_001_708, w_000_523);
  or2  I001_709(w_001_709, w_000_926, w_000_927);
  or2  I001_710(w_001_710, w_000_928, w_000_353);
  nand2 I001_711(w_001_711, w_000_724, w_000_754);
  not1 I001_712(w_001_712, w_000_929);
  not1 I001_714(w_001_714, w_000_158);
  and2 I001_715(w_001_715, w_000_023, w_000_641);
  or2  I001_716(w_001_716, w_000_111, w_000_930);
  not1 I001_717(w_001_717, w_000_260);
  not1 I001_718(w_001_718, w_000_931);
  or2  I001_720(w_001_720, w_000_781, w_000_439);
  not1 I001_721(w_001_721, w_000_017);
  not1 I001_722(w_001_722, w_000_933);
  or2  I001_723(w_001_723, w_000_511, w_000_674);
  or2  I001_725(w_001_725, w_000_566, w_000_935);
  or2  I001_726(w_001_726, w_000_161, w_000_936);
  not1 I001_728(w_001_728, w_000_937);
  or2  I001_729(w_001_729, w_000_938, w_000_939);
  not1 I001_731(w_001_731, w_000_942);
  and2 I001_732(w_001_732, w_000_943, w_000_277);
  not1 I001_733(w_001_733, w_000_136);
  nand2 I001_734(w_001_734, w_000_693, w_000_037);
  not1 I001_735(w_001_735, w_000_944);
  nand2 I001_736(w_001_736, w_000_212, w_000_945);
  not1 I001_737(w_001_737, w_000_946);
  or2  I001_738(w_001_738, w_000_095, w_000_674);
  not1 I001_741(w_001_741, w_000_851);
  or2  I001_742(w_001_742, w_000_948, w_000_949);
  not1 I001_744(w_001_744, w_000_169);
  nand2 I001_745(w_001_745, w_000_563, w_000_951);
  nand2 I001_746(w_001_746, w_000_952, w_000_180);
  and2 I001_747(w_001_747, w_000_297, w_000_953);
  not1 I001_750(w_001_750, w_000_955);
  and2 I001_751(w_001_751, w_000_416, w_000_052);
  not1 I001_752(w_001_752, w_000_956);
  not1 I001_754(w_001_754, w_000_958);
  nand2 I001_755(w_001_755, w_000_949, w_000_790);
  nand2 I001_756(w_001_756, w_000_959, w_000_960);
  not1 I001_757(w_001_757, w_000_961);
  nand2 I001_758(w_001_758, w_000_229, w_000_962);
  and2 I001_759(w_001_759, w_000_963, w_000_964);
  and2 I001_761(w_001_761, w_000_966, w_000_967);
  not1 I001_762(w_001_762, w_000_968);
  not1 I001_763(w_001_763, w_000_759);
  and2 I001_764(w_001_764, w_000_969, w_000_384);
  nand2 I001_765(w_001_765, w_000_970, w_000_971);
  not1 I001_767(w_001_767, w_000_835);
  nand2 I001_768(w_001_768, w_000_450, w_000_972);
  not1 I001_769(w_001_769, w_000_973);
  not1 I001_770(w_001_770, w_000_974);
  not1 I001_771(w_001_771, w_000_264);
  nand2 I001_772(w_001_772, w_000_758, w_000_853);
  not1 I001_776(w_001_776, w_000_472);
  or2  I001_778(w_001_778, w_000_632, w_000_249);
  nand2 I001_779(w_001_779, w_000_980, w_000_376);
  not1 I001_780(w_001_780, w_000_981);
  not1 I001_781(w_001_781, w_000_982);
  nand2 I001_783(w_001_783, w_000_014, w_000_984);
  or2  I001_784(w_001_784, w_000_958, w_000_430);
  not1 I001_785(w_001_785, w_000_985);
  nand2 I001_786(w_001_786, w_000_659, w_000_986);
  nand2 I001_787(w_001_787, w_000_987, w_000_313);
  nand2 I001_790(w_001_790, w_000_988, w_000_712);
  nand2 I001_791(w_001_791, w_000_989, w_000_313);
  not1 I001_792(w_001_792, w_000_513);
  and2 I001_793(w_001_793, w_000_096, w_000_990);
  and2 I001_794(w_001_794, w_000_110, w_000_991);
  nand2 I001_796(w_001_796, w_000_993, w_000_994);
  not1 I001_797(w_001_797, w_000_995);
  and2 I001_798(w_001_798, w_000_008, w_000_996);
  and2 I001_799(w_001_799, w_000_726, w_000_295);
  or2  I001_800(w_001_800, w_000_997, w_000_998);
  and2 I001_801(w_001_801, w_000_857, w_000_251);
  or2  I001_804(w_001_804, w_000_999, w_000_626);
  or2  I001_805(w_001_805, w_000_1000, w_000_325);
  not1 I001_806(w_001_806, w_000_1001);
  not1 I001_807(w_001_807, w_000_589);
  and2 I001_808(w_001_808, w_000_1002, w_000_795);
  not1 I001_809(w_001_809, w_000_784);
  nand2 I001_810(w_001_810, w_000_1003, w_000_840);
  not1 I001_811(w_001_811, w_000_155);
  or2  I001_812(w_001_812, w_000_1004, w_000_1005);
  not1 I001_813(w_001_813, w_000_505);
  not1 I001_814(w_001_814, w_000_1006);
  nand2 I001_815(w_001_815, w_000_863, w_000_1007);
  not1 I001_816(w_001_816, w_000_408);
  not1 I001_817(w_001_817, w_000_768);
  or2  I001_818(w_001_818, w_000_1008, w_000_1009);
  and2 I001_820(w_001_820, w_000_1010, w_000_1011);
  nand2 I001_821(w_001_821, w_000_1012, w_000_435);
  nand2 I001_822(w_001_822, w_000_1013, w_000_1014);
  or2  I001_824(w_001_824, w_000_1016, w_000_1017);
  not1 I001_825(w_001_825, w_000_1018);
  and2 I001_827(w_001_827, w_000_1020, w_000_1021);
  nand2 I001_828(w_001_828, w_000_1022, w_000_733);
  not1 I001_829(w_001_829, w_000_1023);
  and2 I001_831(w_001_831, w_000_258, w_000_1025);
  and2 I001_832(w_001_832, w_000_1026, w_000_297);
  nand2 I001_833(w_001_833, w_000_1027, w_000_1028);
  or2  I001_835(w_001_835, w_000_1030, w_000_319);
  nand2 I001_836(w_001_836, w_000_1031, w_000_1032);
  and2 I001_837(w_001_837, w_000_719, w_000_896);
  not1 I001_840(w_001_840, w_000_1035);
  or2  I001_842(w_001_842, w_000_858, w_000_1037);
  and2 I001_843(w_001_843, w_000_286, w_000_1038);
  or2  I001_844(w_001_844, w_000_1039, w_000_1040);
  not1 I001_845(w_001_845, w_000_421);
  and2 I001_847(w_001_847, w_000_878, w_000_729);
  nand2 I001_848(w_001_848, w_000_758, w_000_053);
  nand2 I001_849(w_001_849, w_000_007, w_000_772);
  nand2 I001_850(w_001_850, w_000_1041, w_000_1042);
  and2 I001_851(w_001_851, w_000_308, w_000_1043);
  not1 I001_852(w_001_852, w_000_1044);
  not1 I001_853(w_001_853, w_000_485);
  not1 I001_854(w_001_854, w_000_946);
  nand2 I001_855(w_001_855, w_000_1045, w_000_751);
  or2  I001_856(w_001_856, w_000_1046, w_000_833);
  not1 I001_857(w_001_857, w_000_448);
  nand2 I001_859(w_001_859, w_000_1047, w_000_1048);
  or2  I001_860(w_001_860, w_000_1049, w_000_287);
  and2 I001_861(w_001_861, w_000_328, w_000_462);
  nand2 I001_862(w_001_862, w_000_1050, w_000_718);
  not1 I001_864(w_001_864, w_000_861);
  not1 I001_865(w_001_865, w_000_1052);
  nand2 I001_866(w_001_866, w_000_657, w_000_129);
  nand2 I001_867(w_001_867, w_000_1053, w_000_1054);
  and2 I001_868(w_001_868, w_000_1055, w_000_078);
  or2  I001_869(w_001_869, w_000_1056, w_000_1057);
  and2 I001_870(w_001_870, w_000_628, w_000_186);
  not1 I001_872(w_001_872, w_000_865);
  nand2 I001_873(w_001_873, w_000_1058, w_000_848);
  nand2 I001_875(w_001_875, w_000_1055, w_000_1060);
  or2  I001_876(w_001_876, w_000_589, w_000_1061);
  and2 I001_877(w_001_877, w_000_1062, w_000_1063);
  nand2 I001_878(w_001_878, w_000_893, w_000_1042);
  and2 I001_879(w_001_879, w_000_1064, w_000_1065);
  or2  I001_880(w_001_880, w_000_1066, w_000_550);
  or2  I001_881(w_001_881, w_000_056, w_000_737);
  not1 I001_882(w_001_882, w_000_241);
  not1 I001_883(w_001_883, w_000_1067);
  not1 I001_884(w_001_884, w_000_1068);
  or2  I001_885(w_001_885, w_000_658, w_000_264);
  nand2 I001_887(w_001_887, w_000_1070, w_000_1071);
  and2 I001_888(w_001_888, w_000_499, w_000_763);
  not1 I001_889(w_001_889, w_000_263);
  not1 I001_890(w_001_890, w_000_399);
  or2  I001_892(w_001_892, w_000_111, w_000_129);
  and2 I001_893(w_001_893, w_000_012, w_000_186);
  or2  I001_894(w_001_894, w_000_1055, w_000_779);
  nand2 I001_895(w_001_895, w_000_979, w_000_589);
  or2  I001_897(w_001_897, w_000_995, w_000_880);
  and2 I001_898(w_001_898, w_000_211, w_000_1075);
  and2 I001_899(w_001_899, w_000_711, w_000_1076);
  nand2 I001_900(w_001_900, w_000_1077, w_000_784);
  not1 I001_901(w_001_901, w_000_632);
  nand2 I001_902(w_001_902, w_000_096, w_000_1078);
  not1 I001_903(w_001_903, w_000_225);
  or2  I001_904(w_001_904, w_000_1079, w_000_763);
  not1 I001_905(w_001_905, w_000_286);
  not1 I001_906(w_001_906, w_000_894);
  or2  I001_907(w_001_907, w_000_835, w_000_1080);
  not1 I001_908(w_001_908, w_000_082);
  or2  I001_909(w_001_909, w_000_053, w_000_1081);
  or2  I001_910(w_001_910, w_000_617, w_000_1082);
  not1 I001_911(w_001_911, w_000_1083);
  nand2 I001_914(w_001_914, w_000_131, w_000_1085);
  not1 I001_915(w_001_915, w_000_709);
  or2  I001_916(w_001_916, w_000_1086, w_000_1087);
  not1 I001_919(w_001_919, w_000_485);
  and2 I001_921(w_001_921, w_000_656, w_000_388);
  or2  I001_922(w_001_922, w_000_1089, w_000_738);
  not1 I001_926(w_001_926, w_000_942);
  and2 I001_929(w_001_929, w_000_1094, w_000_1095);
  nand2 I001_931(w_001_931, w_000_1096, w_000_1097);
  and2 I001_932(w_001_932, w_000_110, w_000_702);
  or2  I001_936(w_001_936, w_000_946, w_000_1102);
  and2 I001_937(w_001_937, w_000_1103, w_000_850);
  and2 I001_939(w_001_939, w_000_1105, w_000_1106);
  not1 I001_940(w_001_940, w_000_676);
  or2  I001_941(w_001_941, w_000_253, w_000_1107);
  or2  I001_943(w_001_943, w_000_1108, w_000_1109);
  or2  I001_944(w_001_944, w_000_709, w_000_1110);
  and2 I001_946(w_001_946, w_000_1111, w_000_1112);
  not1 I001_947(w_001_947, w_000_1113);
  and2 I001_948(w_001_948, w_000_029, w_000_264);
  and2 I001_949(w_001_949, w_000_424, w_000_250);
  and2 I001_950(w_001_950, w_000_1114, w_000_1115);
  not1 I001_951(w_001_951, w_000_772);
  nand2 I001_953(w_001_953, w_000_1116, w_000_1117);
  or2  I001_954(w_001_954, w_000_709, w_000_1118);
  not1 I001_955(w_001_955, w_000_1119);
  and2 I001_956(w_001_956, w_000_850, w_000_355);
  nand2 I001_958(w_001_958, w_000_1120, w_000_1121);
  and2 I001_960(w_001_960, w_000_1124, w_000_508);
  or2  I001_961(w_001_961, w_000_1125, w_000_303);
  nand2 I001_963(w_001_963, w_000_1126, w_000_1127);
  nand2 I001_964(w_001_964, w_000_1128, w_000_1129);
  and2 I001_965(w_001_965, w_000_1130, w_000_1131);
  not1 I001_966(w_001_966, w_000_816);
  and2 I001_967(w_001_967, w_000_1132, w_000_1027);
  nand2 I001_969(w_001_969, w_000_226, w_000_1133);
  nand2 I001_970(w_001_970, w_000_1134, w_000_023);
  and2 I001_973(w_001_973, w_000_230, w_000_1138);
  nand2 I001_974(w_001_974, w_000_051, w_000_1139);
  and2 I001_976(w_001_976, w_000_1141, w_000_780);
  not1 I001_977(w_001_977, w_000_493);
  or2  I001_978(w_001_978, w_000_898, w_000_386);
  nand2 I001_980(w_001_980, w_000_202, w_000_626);
  not1 I001_981(w_001_981, w_000_1143);
  or2  I001_982(w_001_982, w_000_1144, w_000_1145);
  or2  I001_983(w_001_983, w_000_146, w_000_1146);
  and2 I001_984(w_001_984, w_000_174, w_000_1147);
  not1 I001_985(w_001_985, w_000_414);
  not1 I001_986(w_001_986, w_000_1148);
  and2 I001_987(w_001_987, w_000_1149, w_000_735);
  nand2 I001_988(w_001_988, w_000_334, w_000_1150);
  and2 I001_989(w_001_989, w_000_635, w_000_507);
  not1 I001_990(w_001_990, w_000_1151);
  nand2 I001_991(w_001_991, w_000_055, w_000_703);
  and2 I001_993(w_001_993, w_000_1153, w_000_1154);
  and2 I001_994(w_001_994, w_000_1155, w_000_1156);
  or2  I001_997(w_001_997, w_000_042, w_000_1043);
  nand2 I001_998(w_001_998, w_000_777, w_000_1159);
  not1 I001_999(w_001_999, w_000_386);
  not1 I001_1000(w_001_1000, w_000_097);
  or2  I001_1001(w_001_1001, w_000_417, w_000_061);
  and2 I001_1002(w_001_1002, w_000_824, w_000_1117);
  not1 I001_1003(w_001_1003, w_000_1160);
  nand2 I001_1005(w_001_1005, w_000_186, w_000_1109);
  not1 I001_1007(w_001_1007, w_000_495);
  not1 I001_1008(w_001_1008, w_000_417);
  not1 I001_1011(w_001_1011, w_000_1165);
  not1 I001_1012(w_001_1012, w_000_403);
  not1 I001_1013(w_001_1013, w_000_1163);
  or2  I001_1014(w_001_1014, w_000_234, w_000_339);
  not1 I001_1015(w_001_1015, w_000_1166);
  and2 I001_1019(w_001_1019, w_000_1171, w_000_1172);
  nand2 I001_1020(w_001_1020, w_000_1004, w_000_361);
  and2 I001_1022(w_001_1022, w_000_327, w_000_050);
  not1 I001_1023(w_001_1023, w_000_1173);
  nand2 I001_1025(w_001_1025, w_000_626, w_000_680);
  not1 I001_1026(w_001_1026, w_000_912);
  and2 I001_1027(w_001_1027, w_000_1175, w_000_157);
  nand2 I001_1028(w_001_1028, w_000_346, w_000_1176);
  and2 I001_1030(w_001_1030, w_000_1178, w_000_1179);
  and2 I001_1031(w_001_1031, w_000_557, w_000_584);
  and2 I001_1033(w_001_1033, w_000_337, w_000_1180);
  not1 I001_1034(w_001_1034, w_000_277);
  or2  I001_1035(w_001_1035, w_000_1181, w_000_1074);
  and2 I001_1036(w_001_1036, w_000_342, w_000_1182);
  not1 I001_1037(w_001_1037, w_000_1183);
  not1 I001_1039(w_001_1039, w_000_225);
  or2  I001_1040(w_001_1040, w_000_902, w_000_827);
  nand2 I001_1042(w_001_1042, w_000_1186, w_000_1187);
  nand2 I001_1044(w_001_1044, w_000_1142, w_000_1189);
  and2 I001_1045(w_001_1045, w_000_696, w_000_619);
  or2  I001_1046(w_001_1046, w_000_412, w_000_1190);
  or2  I001_1047(w_001_1047, w_000_754, w_000_1191);
  not1 I001_1049(w_001_1049, w_000_124);
  or2  I001_1050(w_001_1050, w_000_959, w_000_1193);
  nand2 I001_1051(w_001_1051, w_000_1194, w_000_1195);
  and2 I001_1053(w_001_1053, w_000_1197, w_000_046);
  not1 I001_1054(w_001_1054, w_000_1109);
  or2  I001_1056(w_001_1056, w_000_173, w_000_070);
  not1 I001_1057(w_001_1057, w_000_585);
  and2 I001_1058(w_001_1058, w_000_1199, w_000_1200);
  and2 I001_1059(w_001_1059, w_000_1201, w_000_052);
  nand2 I001_1060(w_001_1060, w_000_368, w_000_176);
  and2 I001_1061(w_001_1061, w_000_1202, w_000_430);
  nand2 I001_1062(w_001_1062, w_000_1203, w_000_037);
  and2 I001_1063(w_001_1063, w_000_1204, w_000_1205);
  and2 I001_1064(w_001_1064, w_000_1206, w_000_1207);
  nand2 I001_1065(w_001_1065, w_000_1208, w_000_1209);
  and2 I001_1066(w_001_1066, w_000_707, w_000_1147);
  or2  I001_1067(w_001_1067, w_000_777, w_000_1157);
  nand2 I001_1068(w_001_1068, w_000_893, w_000_992);
  not1 I001_1070(w_001_1070, w_000_1210);
  and2 I001_1071(w_001_1071, w_000_1211, w_000_431);
  and2 I001_1072(w_001_1072, w_000_1026, w_000_861);
  and2 I001_1074(w_001_1074, w_000_477, w_000_821);
  nand2 I001_1076(w_001_1076, w_000_1212, w_000_780);
  nand2 I001_1077(w_001_1077, w_000_586, w_000_279);
  or2  I001_1078(w_001_1078, w_000_1213, w_000_1214);
  and2 I001_1079(w_001_1079, w_000_609, w_000_428);
  nand2 I001_1081(w_001_1081, w_000_1215, w_000_1027);
  not1 I001_1082(w_001_1082, w_000_1216);
  nand2 I001_1083(w_001_1083, w_000_484, w_000_873);
  nand2 I001_1084(w_001_1084, w_000_1217, w_000_124);
  nand2 I001_1085(w_001_1085, w_000_158, w_000_945);
  not1 I001_1088(w_001_1088, w_000_1218);
  and2 I001_1089(w_001_1089, w_000_155, w_000_962);
  and2 I001_1090(w_001_1090, w_000_1219, w_000_1220);
  and2 I001_1092(w_001_1092, w_000_187, w_000_017);
  not1 I001_1093(w_001_1093, w_000_199);
  and2 I001_1094(w_001_1094, w_000_1221, w_000_1072);
  not1 I001_1096(w_001_1096, w_000_1223);
  not1 I001_1097(w_001_1097, w_000_1098);
  and2 I001_1098(w_001_1098, w_000_582, w_000_1224);
  or2  I001_1099(w_001_1099, w_000_1225, w_000_1226);
  and2 I001_1100(w_001_1100, w_000_1227, w_000_355);
  not1 I001_1101(w_001_1101, w_000_591);
  not1 I001_1102(w_001_1102, w_000_1228);
  and2 I001_1104(w_001_1104, w_000_1229, w_000_545);
  not1 I001_1105(w_001_1105, w_000_034);
  or2  I001_1106(w_001_1106, w_000_1230, w_000_1107);
  or2  I001_1107(w_001_1107, w_000_996, w_000_655);
  nand2 I001_1108(w_001_1108, w_000_606, w_000_1149);
  or2  I001_1109(w_001_1109, w_000_1231, w_000_083);
  not1 I001_1111(w_001_1111, w_000_850);
  nand2 I001_1112(w_001_1112, w_000_1232, w_000_1205);
  or2  I001_1113(w_001_1113, w_000_835, w_000_1191);
  nand2 I001_1115(w_001_1115, w_000_1234, w_000_323);
  not1 I001_1117(w_001_1117, w_000_1236);
  or2  I001_1118(w_001_1118, w_000_091, w_000_650);
  and2 I001_1119(w_001_1119, w_000_1237, w_000_1238);
  not1 I001_1120(w_001_1120, w_000_388);
  not1 I001_1121(w_001_1121, w_000_057);
  not1 I001_1122(w_001_1122, w_000_1239);
  nand2 I001_1123(w_001_1123, w_000_240, w_000_768);
  and2 I001_1124(w_001_1124, w_000_1240, w_000_141);
  nand2 I001_1125(w_001_1125, w_000_1241, w_000_1053);
  nand2 I001_1126(w_001_1126, w_000_1242, w_000_844);
  not1 I001_1127(w_001_1127, w_000_152);
  or2  I001_1128(w_001_1128, w_000_1243, w_000_510);
  nand2 I001_1129(w_001_1129, w_000_970, w_000_327);
  not1 I001_1130(w_001_1130, w_000_1244);
  and2 I001_1131(w_001_1131, w_000_040, w_000_1245);
  not1 I001_1132(w_001_1132, w_000_780);
  not1 I001_1133(w_001_1133, w_000_831);
  nand2 I001_1134(w_001_1134, w_000_1246, w_000_1247);
  nand2 I001_1135(w_001_1135, w_000_1019, w_000_019);
  or2  I001_1138(w_001_1138, w_000_083, w_000_1250);
  and2 I001_1140(w_001_1140, w_000_1252, w_000_1253);
  not1 I001_1141(w_001_1141, w_000_129);
  and2 I001_1142(w_001_1142, w_000_1138, w_000_929);
  and2 I001_1143(w_001_1143, w_000_718, w_000_055);
  or2  I001_1144(w_001_1144, w_000_1254, w_000_887);
  and2 I001_1145(w_001_1145, w_000_1255, w_000_718);
  nand2 I001_1146(w_001_1146, w_000_878, w_000_737);
  and2 I001_1147(w_001_1147, w_000_390, w_000_835);
  not1 I001_1148(w_001_1148, w_000_1256);
  or2  I001_1149(w_001_1149, w_000_317, w_000_1257);
  or2  I001_1151(w_001_1151, w_000_707, w_000_623);
  nand2 I001_1152(w_001_1152, w_000_836, w_000_879);
  or2  I001_1153(w_001_1153, w_000_118, w_000_1258);
  nand2 I001_1155(w_001_1155, w_000_1259, w_000_908);
  not1 I001_1156(w_001_1156, w_000_130);
  and2 I001_1158(w_001_1158, w_000_046, w_000_055);
  nand2 I001_1159(w_001_1159, w_000_1261, w_000_212);
  and2 I001_1160(w_001_1160, w_000_1128, w_000_897);
  or2  I001_1161(w_001_1161, w_000_197, w_000_130);
  or2  I001_1163(w_001_1163, w_000_403, w_000_418);
  nand2 I001_1164(w_001_1164, w_000_283, w_000_1262);
  nand2 I001_1167(w_001_1167, w_000_828, w_000_026);
  nand2 I001_1170(w_001_1170, w_000_1094, w_000_1265);
  nand2 I001_1171(w_001_1171, w_000_1266, w_000_1249);
  or2  I001_1172(w_001_1172, w_000_473, w_000_074);
  nand2 I001_1176(w_001_1176, w_000_1271, w_000_943);
  nand2 I001_1177(w_001_1177, w_000_167, w_000_1272);
  and2 I001_1179(w_001_1179, w_000_617, w_000_1204);
  nand2 I001_1181(w_001_1181, w_000_008, w_000_289);
  nand2 I001_1183(w_001_1183, w_000_1150, w_000_116);
  not1 I001_1184(w_001_1184, w_000_887);
  and2 I001_1185(w_001_1185, w_000_1274, w_000_1259);
  or2  I001_1186(w_001_1186, w_000_446, w_000_1223);
  not1 I001_1187(w_001_1187, w_000_1275);
  not1 I001_1188(w_001_1188, w_000_1276);
  or2  I001_1189(w_001_1189, w_000_1277, w_000_250);
  nand2 I001_1191(w_001_1191, w_000_921, w_000_1278);
  or2  I001_1192(w_001_1192, w_000_865, w_000_1279);
  not1 I001_1193(w_001_1193, w_000_058);
  nand2 I001_1195(w_001_1195, w_000_1282, w_000_679);
  nand2 I001_1196(w_001_1196, w_000_228, w_000_251);
  not1 I001_1197(w_001_1197, w_000_1283);
  or2  I001_1198(w_001_1198, w_000_313, w_000_1284);
  nand2 I001_1199(w_001_1199, w_000_352, w_000_1285);
  and2 I001_1200(w_001_1200, w_000_386, w_000_166);
  nand2 I001_1201(w_001_1201, w_000_1200, w_000_1286);
  not1 I001_1202(w_001_1202, w_000_473);
  or2  I001_1203(w_001_1203, w_000_579, w_000_1287);
  or2  I001_1204(w_001_1204, w_000_1288, w_000_1289);
  not1 I001_1205(w_001_1205, w_000_857);
  or2  I001_1206(w_001_1206, w_000_1290, w_000_845);
  and2 I001_1207(w_001_1207, w_000_1193, w_000_1291);
  or2  I001_1209(w_001_1209, w_000_949, w_000_1293);
  or2  I001_1211(w_001_1211, w_000_039, w_000_276);
  nand2 I001_1212(w_001_1212, w_000_1296, w_000_1091);
  and2 I001_1213(w_001_1213, w_000_1130, w_000_022);
  nand2 I001_1215(w_001_1215, w_000_526, w_000_569);
  or2  I001_1216(w_001_1216, w_000_240, w_000_1298);
  or2  I001_1217(w_001_1217, w_000_1299, w_000_1192);
  and2 I001_1220(w_001_1220, w_000_1301, w_000_1023);
  not1 I001_1221(w_001_1221, w_000_975);
  not1 I001_1222(w_001_1222, w_000_1161);
  or2  I001_1225(w_001_1225, w_000_1176, w_000_177);
  or2  I001_1226(w_001_1226, w_000_680, w_000_1055);
  nand2 I001_1227(w_001_1227, w_000_1257, w_000_1296);
  not1 I001_1228(w_001_1228, w_000_1303);
  or2  I001_1229(w_001_1229, w_000_1304, w_000_1305);
  not1 I001_1230(w_001_1230, w_000_1249);
  or2  I001_1231(w_001_1231, w_000_1224, w_000_146);
  and2 I001_1232(w_001_1232, w_000_247, w_000_916);
  nand2 I001_1233(w_001_1233, w_000_1306, w_000_077);
  not1 I001_1235(w_001_1235, w_000_440);
  or2  I001_1236(w_001_1236, w_000_1307, w_000_1308);
  not1 I001_1237(w_001_1237, w_000_349);
  and2 I001_1238(w_001_1238, w_000_1021, w_000_1309);
  or2  I001_1239(w_001_1239, w_000_669, w_000_466);
  and2 I001_1240(w_001_1240, w_000_1310, w_000_777);
  nand2 I001_1241(w_001_1241, w_000_1311, w_000_026);
  or2  I001_1242(w_001_1242, w_000_830, w_000_172);
  or2  I001_1243(w_001_1243, w_000_1312, w_000_1088);
  not1 I001_1246(w_001_1246, w_000_901);
  nand2 I001_1247(w_001_1247, w_000_1315, w_000_870);
  or2  I001_1248(w_001_1248, w_000_696, w_000_1316);
  not1 I001_1249(w_001_1249, w_000_396);
  and2 I001_1250(w_001_1250, w_000_332, w_000_863);
  and2 I001_1251(w_001_1251, w_000_435, w_000_1317);
  and2 I001_1253(w_001_1253, w_000_1222, w_000_543);
  not1 I001_1255(w_001_1255, w_000_447);
  or2  I001_1256(w_001_1256, w_000_878, w_000_908);
  and2 I001_1259(w_001_1259, w_000_1320, w_000_347);
  not1 I001_1260(w_001_1260, w_000_1321);
  nand2 I001_1261(w_001_1261, w_000_326, w_000_050);
  not1 I001_1262(w_001_1262, w_000_298);
  or2  I001_1263(w_001_1263, w_000_1322, w_000_498);
  or2  I001_1264(w_001_1264, w_000_1323, w_000_1324);
  and2 I001_1265(w_001_1265, w_000_512, w_000_576);
  and2 I001_1266(w_001_1266, w_000_847, w_000_1325);
  nand2 I001_1267(w_001_1267, w_000_349, w_000_1108);
  nand2 I001_1268(w_001_1268, w_000_736, w_000_764);
  or2  I001_1269(w_001_1269, w_000_151, w_000_415);
  or2  I001_1270(w_001_1270, w_000_1326, w_000_1114);
  and2 I001_1271(w_001_1271, w_000_1220, w_000_210);
  not1 I001_1272(w_001_1272, w_000_1270);
  and2 I001_1273(w_001_1273, w_000_941, w_000_107);
  nand2 I001_1274(w_001_1274, w_000_1327, w_000_1328);
  and2 I001_1275(w_001_1275, w_000_1189, w_000_493);
  and2 I001_1276(w_001_1276, w_000_117, w_000_653);
  and2 I001_1278(w_001_1278, w_000_1329, w_000_423);
  or2  I001_1279(w_001_1279, w_000_572, w_000_101);
  and2 I001_1280(w_001_1280, w_000_1330, w_000_1162);
  not1 I001_1281(w_001_1281, w_000_454);
  not1 I001_1282(w_001_1282, w_000_1331);
  and2 I001_1284(w_001_1284, w_000_710, w_000_1249);
  nand2 I001_1288(w_001_1288, w_000_1211, w_000_1334);
  nand2 I001_1289(w_001_1289, w_000_1019, w_000_471);
  and2 I001_1290(w_001_1290, w_000_1335, w_000_924);
  not1 I001_1293(w_001_1293, w_000_752);
  and2 I001_1296(w_001_1296, w_000_897, w_000_1338);
  nand2 I001_1298(w_001_1298, w_000_156, w_000_617);
  not1 I001_1299(w_001_1299, w_000_1340);
  or2  I001_1300(w_001_1300, w_000_322, w_000_386);
  or2  I001_1301(w_001_1301, w_000_074, w_000_1341);
  or2  I001_1302(w_001_1302, w_000_271, w_000_908);
  and2 I001_1303(w_001_1303, w_000_766, w_000_996);
  not1 I001_1304(w_001_1304, w_000_780);
  or2  I001_1305(w_001_1305, w_000_1342, w_000_1343);
  not1 I001_1306(w_001_1306, w_000_1344);
  and2 I001_1307(w_001_1307, w_000_334, w_000_1046);
  not1 I001_1308(w_001_1308, w_000_1345);
  not1 I001_1309(w_001_1309, w_000_216);
  not1 I001_1310(w_001_1310, w_000_846);
  nand2 I001_1312(w_001_1312, w_000_1347, w_000_952);
  or2  I001_1314(w_001_1314, w_000_864, w_000_190);
  not1 I001_1316(w_001_1316, w_000_672);
  not1 I001_1317(w_001_1317, w_000_1287);
  or2  I001_1319(w_001_1319, w_000_1349, w_000_1350);
  and2 I001_1320(w_001_1320, w_000_1351, w_000_1352);
  not1 I001_1321(w_001_1321, w_000_1353);
  and2 I001_1322(w_001_1322, w_000_1354, w_000_1355);
  or2  I001_1323(w_001_1323, w_000_075, w_000_1356);
  nand2 I001_1324(w_001_1324, w_000_1027, w_000_720);
  and2 I001_1325(w_001_1325, w_000_309, w_000_474);
  not1 I001_1327(w_001_1327, w_000_038);
  nand2 I001_1331(w_001_1331, w_000_370, w_000_147);
  or2  I001_1332(w_001_1332, w_000_1032, w_000_491);
  not1 I001_1333(w_001_1333, w_000_541);
  or2  I001_1335(w_001_1335, w_000_1359, w_000_1360);
  or2  I001_1337(w_001_1337, w_000_1361, w_000_1362);
  nand2 I001_1339(w_001_1339, w_000_836, w_000_1258);
  nand2 I001_1341(w_001_1341, w_000_1363, w_000_964);
  not1 I001_1342(w_001_1342, w_000_132);
  nand2 I001_1343(w_001_1343, w_000_1348, w_000_1165);
  and2 I001_1345(w_001_1345, w_000_437, w_000_1027);
  or2  I001_1346(w_001_1346, w_000_375, w_000_1023);
  nand2 I001_1349(w_001_1349, w_000_472, w_000_032);
  nand2 I001_1350(w_001_1350, w_000_082, w_000_905);
  and2 I001_1351(w_001_1351, w_000_675, w_000_428);
  nand2 I001_1353(w_001_1353, w_000_443, w_000_1365);
  nand2 I001_1354(w_001_1354, w_000_1366, w_000_1367);
  or2  I001_1355(w_001_1355, w_000_370, w_000_441);
  not1 I001_1356(w_001_1356, w_000_1368);
  not1 I001_1358(w_001_1358, w_000_1369);
  or2  I001_1359(w_001_1359, w_000_1370, w_000_902);
  not1 I001_1361(w_001_1361, w_000_1323);
  or2  I001_1362(w_001_1362, w_000_1372, w_000_228);
  not1 I001_1365(w_001_1365, w_000_1373);
  not1 I001_1366(w_001_1366, w_000_190);
  not1 I001_1367(w_001_1367, w_000_947);
  not1 I001_1369(w_001_1369, w_000_1007);
  nand2 I001_1371(w_001_1371, w_000_1375, w_000_1243);
  nand2 I001_1373(w_001_1373, w_000_149, w_000_1376);
  nand2 I001_1374(w_001_1374, w_000_377, w_000_1377);
  or2  I001_1376(w_001_1376, w_000_417, w_000_1379);
  and2 I001_1379(w_001_1379, w_000_1382, w_000_753);
  nand2 I001_1380(w_001_1380, w_000_956, w_000_856);
  not1 I001_1381(w_001_1381, w_000_801);
  nand2 I001_1382(w_001_1382, w_000_150, w_000_397);
  and2 I001_1383(w_001_1383, w_000_976, w_000_1383);
  nand2 I001_1384(w_001_1384, w_000_1126, w_000_008);
  nand2 I001_1386(w_001_1386, w_000_1277, w_000_1385);
  or2  I001_1387(w_001_1387, w_000_1386, w_000_011);
  not1 I001_1388(w_001_1388, w_000_1387);
  not1 I001_1390(w_001_1390, w_000_1174);
  nand2 I001_1392(w_001_1392, w_000_1389, w_000_967);
  or2  I001_1393(w_001_1393, w_000_218, w_000_1390);
  not1 I001_1394(w_001_1394, w_000_1391);
  or2  I001_1396(w_001_1396, w_000_1393, w_000_1394);
  and2 I001_1397(w_001_1397, w_000_1395, w_000_1396);
  or2  I001_1398(w_001_1398, w_000_1397, w_000_664);
  and2 I001_1399(w_001_1399, w_000_1398, w_000_1015);
  not1 I001_1400(w_001_1400, w_000_215);
  nand2 I001_1402(w_001_1402, w_000_352, w_000_757);
  or2  I001_1403(w_001_1403, w_000_1027, w_000_260);
  not1 I001_1405(w_001_1405, w_000_1082);
  or2  I001_1406(w_001_1406, w_000_788, w_000_1046);
  nand2 I001_1408(w_001_1408, w_000_491, w_000_1399);
  and2 I001_1409(w_001_1409, w_000_216, w_000_466);
  nand2 I001_1412(w_001_1412, w_000_981, w_000_001);
  nand2 I001_1413(w_001_1413, w_000_090, w_000_1202);
  not1 I001_1416(w_001_1416, w_000_411);
  or2  I001_1417(w_001_1417, w_000_1402, w_000_946);
  or2  I001_1418(w_001_1418, w_000_1191, w_000_1403);
  or2  I001_1422(w_001_1422, w_000_797, w_000_1406);
  not1 I001_1423(w_001_1423, w_000_799);
  and2 I001_1424(w_001_1424, w_000_280, w_000_353);
  nand2 I001_1425(w_001_1425, w_000_1334, w_000_428);
  nand2 I001_1426(w_001_1426, w_000_1220, w_000_845);
  or2  I001_1427(w_001_1427, w_000_1407, w_000_050);
  or2  I001_1428(w_001_1428, w_000_929, w_000_319);
  and2 I001_1429(w_001_1429, w_000_1270, w_000_1080);
  or2  I001_1430(w_001_1430, w_000_1143, w_000_409);
  nand2 I001_1431(w_001_1431, w_000_866, w_000_394);
  nand2 I001_1432(w_001_1432, w_000_003, w_000_1408);
  or2  I001_1435(w_001_1435, w_000_952, w_000_112);
  or2  I001_1436(w_001_1436, w_000_1063, w_000_1332);
  nand2 I001_1437(w_001_1437, w_000_1244, w_000_1315);
  or2  I001_1438(w_001_1438, w_000_1246, w_000_244);
  or2  I001_1439(w_001_1439, w_000_790, w_000_1411);
  or2  I001_1440(w_001_1440, w_000_1327, w_000_1009);
  not1 I001_1441(w_001_1441, w_000_1412);
  nand2 I001_1444(w_001_1444, w_000_625, w_000_042);
  or2  I001_1446(w_001_1446, w_000_1414, w_000_1056);
  and2 I001_1447(w_001_1447, w_000_847, w_000_975);
  nand2 I001_1449(w_001_1449, w_000_758, w_000_1415);
  and2 I001_1452(w_001_1452, w_000_1418, w_000_1017);
  not1 I001_1453(w_001_1453, w_000_092);
  or2  I001_1454(w_001_1454, w_000_1419, w_000_215);
  not1 I001_1456(w_001_1456, w_000_157);
  or2  I001_1457(w_001_1457, w_000_1421, w_000_1422);
  or2  I001_1458(w_001_1458, w_000_592, w_000_541);
  not1 I001_1459(w_001_1459, w_000_1423);
  not1 I001_1460(w_001_1460, w_000_585);
  and2 I001_1461(w_001_1461, w_000_1424, w_000_539);
  and2 I001_1462(w_001_1462, w_000_1083, w_000_172);
  or2  I001_1463(w_001_1463, w_000_872, w_000_1425);
  not1 I001_1464(w_001_1464, w_000_242);
  not1 I001_1465(w_001_1465, w_000_1426);
  not1 I001_1467(w_001_1467, w_000_409);
  not1 I001_1469(w_001_1469, w_000_1427);
  or2  I001_1470(w_001_1470, w_000_484, w_000_908);
  nand2 I001_1474(w_001_1474, w_000_076, w_000_1430);
  or2  I001_1475(w_001_1475, w_000_1301, w_000_1431);
  nand2 I001_1476(w_001_1476, w_000_1432, w_000_969);
  not1 I001_1477(w_001_1477, w_000_1433);
  or2  I001_1479(w_001_1479, w_000_1434, w_000_757);
  nand2 I001_1480(w_001_1480, w_000_1241, w_000_003);
  not1 I001_1482(w_001_1482, w_000_480);
  and2 I001_1483(w_001_1483, w_000_1018, w_000_1397);
  nand2 I001_1484(w_001_1484, w_000_011, w_000_1204);
  nand2 I001_1485(w_001_1485, w_000_440, w_000_1184);
  and2 I001_1486(w_001_1486, w_000_093, w_000_1347);
  nand2 I001_1487(w_001_1487, w_000_1435, w_000_317);
  or2  I001_1488(w_001_1488, w_000_1436, w_000_1437);
  or2  I001_1489(w_001_1489, w_000_1438, w_000_190);
  and2 I001_1491(w_001_1491, w_000_696, w_000_201);
  and2 I001_1495(w_001_1495, w_000_1385, w_000_1440);
  nand2 I001_1496(w_001_1496, w_000_177, w_000_1300);
  nand2 I001_1497(w_001_1497, w_000_270, w_000_647);
  not1 I001_1498(w_001_1498, w_000_258);
  and2 I001_1499(w_001_1499, w_000_1441, w_000_585);
  or2  I001_1500(w_001_1500, w_000_773, w_000_168);
  or2  I001_1502(w_001_1502, w_000_1189, w_000_1442);
  not1 I001_1503(w_001_1503, w_000_1443);
  not1 I001_1505(w_001_1505, w_000_1444);
  and2 I001_1506(w_001_1506, w_000_1241, w_000_1366);
  or2  I001_1507(w_001_1507, w_000_1357, w_000_669);
  nand2 I001_1508(w_001_1508, w_000_657, w_000_724);
  or2  I001_1509(w_001_1509, w_000_1305, w_000_1445);
  or2  I001_1511(w_001_1511, w_000_1447, w_000_304);
  nand2 I001_1513(w_001_1513, w_000_1051, w_000_1207);
  and2 I001_1514(w_001_1514, w_000_762, w_000_1078);
  not1 I001_1515(w_001_1515, w_000_828);
  and2 I001_1516(w_001_1516, w_000_085, w_000_268);
  not1 I001_1517(w_001_1517, w_000_1449);
  not1 I001_1520(w_001_1520, w_000_1026);
  and2 I001_1521(w_001_1521, w_000_662, w_000_1295);
  nand2 I001_1522(w_001_1522, w_000_1131, w_000_1106);
  and2 I001_1523(w_001_1523, w_000_120, w_000_649);
  or2  I001_1524(w_001_1524, w_000_323, w_000_1450);
  nand2 I001_1526(w_001_1526, w_000_290, w_000_1452);
  nand2 I001_1527(w_001_1527, w_000_375, w_000_262);
  or2  I001_1529(w_001_1529, w_000_300, w_000_860);
  not1 I001_1531(w_001_1531, w_000_824);
  not1 I001_1532(w_001_1532, w_000_300);
  nand2 I001_1533(w_001_1533, w_000_789, w_000_1431);
  not1 I001_1534(w_001_1534, w_000_1454);
  nand2 I001_1536(w_001_1536, w_000_279, w_000_707);
  not1 I001_1538(w_001_1538, w_000_1088);
  nand2 I001_1540(w_001_1540, w_000_1279, w_000_1455);
  nand2 I001_1541(w_001_1541, w_000_1356, w_000_160);
  and2 I001_1544(w_001_1544, w_000_914, w_000_450);
  not1 I001_1547(w_001_1547, w_000_1457);
  not1 I001_1548(w_001_1548, w_000_1037);
  nand2 I001_1550(w_001_1550, w_000_1459, w_000_1460);
  and2 I001_1551(w_001_1551, w_000_1461, w_000_837);
  nand2 I001_1555(w_001_1555, w_000_799, w_000_129);
  or2  I001_1556(w_001_1556, w_000_1466, w_000_509);
  and2 I001_1557(w_001_1557, w_000_803, w_000_1467);
  not1 I001_1559(w_001_1559, w_000_1183);
  or2  I001_1560(w_001_1560, w_000_095, w_000_827);
  and2 I001_1561(w_001_1561, w_000_220, w_000_737);
  not1 I001_1563(w_001_1563, w_000_1469);
  or2  I001_1564(w_001_1564, w_000_303, w_000_909);
  or2  I001_1565(w_001_1565, w_000_463, w_000_442);
  and2 I001_1566(w_001_1566, w_000_1470, w_000_1471);
  or2  I001_1567(w_001_1567, w_000_319, w_000_1442);
  not1 I001_1568(w_001_1568, w_000_487);
  or2  I001_1570(w_001_1570, w_000_777, w_000_169);
  nand2 I001_1571(w_001_1571, w_000_872, w_000_1348);
  and2 I001_1573(w_001_1573, w_000_1140, w_000_365);
  not1 I001_1575(w_001_1575, w_000_1070);
  and2 I001_1576(w_001_1576, w_000_1472, w_000_1473);
  nand2 I001_1578(w_001_1578, w_000_779, w_000_957);
  nand2 I001_1579(w_001_1579, w_000_221, w_000_504);
  not1 I001_1580(w_001_1580, w_000_818);
  not1 I001_1581(w_001_1581, w_000_1474);
  and2 I001_1582(w_001_1582, w_000_999, w_000_089);
  nand2 I001_1583(w_001_1583, w_000_1475, w_000_1476);
  nand2 I001_1585(w_001_1585, w_000_983, w_000_455);
  and2 I001_1586(w_001_1586, w_000_1477, w_000_1478);
  not1 I001_1587(w_001_1587, w_000_819);
  nand2 I001_1588(w_001_1588, w_000_202, w_000_704);
  or2  I001_1589(w_001_1589, w_000_474, w_000_128);
  or2  I001_1592(w_001_1592, w_000_393, w_000_862);
  or2  I001_1593(w_001_1593, w_000_145, w_000_213);
  or2  I001_1595(w_001_1595, w_000_956, w_000_1480);
  and2 I001_1597(w_001_1597, w_000_480, w_000_467);
  not1 I001_1599(w_001_1599, w_000_1481);
  and2 I001_1600(w_001_1600, w_000_1482, w_000_1403);
  and2 I001_1602(w_001_1602, w_000_1483, w_000_1046);
  not1 I001_1603(w_001_1603, w_000_417);
  nand2 I001_1604(w_001_1604, w_000_371, w_000_1279);
  or2  I001_1605(w_001_1605, w_000_868, w_000_1484);
  nand2 I001_1606(w_001_1606, w_000_584, w_000_282);
  nand2 I001_1607(w_001_1607, w_000_319, w_000_034);
  nand2 I001_1608(w_001_1608, w_000_1388, w_000_594);
  nand2 I001_1609(w_001_1609, w_000_207, w_000_1485);
  or2  I001_1612(w_001_1612, w_000_604, w_000_660);
  or2  I001_1613(w_001_1613, w_000_382, w_000_058);
  and2 I001_1616(w_001_1616, w_000_276, w_000_1046);
  and2 I001_1617(w_001_1617, w_000_558, w_000_1153);
  not1 I001_1622(w_001_1622, w_000_456);
  not1 I001_1625(w_001_1625, w_000_758);
  or2  I001_1627(w_001_1627, w_000_228, w_000_073);
  not1 I001_1628(w_001_1628, w_000_1490);
  not1 I001_1629(w_001_1629, w_000_728);
  and2 I001_1630(w_001_1630, w_000_737, w_000_1491);
  and2 I001_1631(w_001_1631, w_000_1145, w_000_1492);
  and2 I001_1632(w_001_1632, w_000_1409, w_000_1253);
  or2  I001_1633(w_001_1633, w_000_1493, w_000_624);
  and2 I001_1634(w_001_1634, w_000_169, w_000_1433);
  or2  I001_1636(w_001_1636, w_000_496, w_000_1495);
  nand2 I001_1637(w_001_1637, w_000_478, w_000_510);
  or2  I001_1638(w_001_1638, w_000_1058, w_000_936);
  nand2 I001_1639(w_001_1639, w_000_685, w_000_1358);
  nand2 I001_1640(w_001_1640, w_000_1465, w_000_447);
  or2  I001_1641(w_001_1641, w_000_1041, w_000_1496);
  not1 I001_1642(w_001_1642, w_000_1497);
  not1 I001_1643(w_001_1643, w_000_699);
  not1 I001_1644(w_001_1644, w_000_1224);
  and2 I001_1645(w_001_1645, w_000_1498, w_000_1499);
  or2  I001_1646(w_001_1646, w_000_218, w_000_1225);
  and2 I001_1647(w_001_1647, w_000_523, w_000_1500);
  nand2 I001_1649(w_001_1649, w_000_896, w_000_1502);
  or2  I001_1651(w_001_1651, w_000_1503, w_000_111);
  not1 I001_1653(w_001_1653, w_000_853);
  not1 I001_1654(w_001_1654, w_000_296);
  or2  I001_1655(w_001_1655, w_000_1505, w_000_1506);
  or2  I001_1656(w_001_1656, w_000_1307, w_000_1507);
  not1 I001_1657(w_001_1657, w_000_1508);
  and2 I001_1659(w_001_1659, w_000_1509, w_000_692);
  nand2 I001_1660(w_001_1660, w_000_1510, w_000_1511);
  and2 I001_1661(w_001_1661, w_000_1074, w_000_315);
  nand2 I001_1662(w_001_1662, w_000_1512, w_000_545);
  or2  I001_1664(w_001_1664, w_000_1339, w_000_1513);
  not1 I001_1665(w_001_1665, w_000_734);
  not1 I001_1666(w_001_1666, w_000_1415);
  nand2 I001_1667(w_001_1667, w_000_435, w_000_1514);
  not1 I001_1669(w_001_1669, w_000_060);
  and2 I001_1670(w_001_1670, w_000_032, w_000_813);
  and2 I001_1671(w_001_1671, w_000_011, w_000_1515);
  nand2 I001_1672(w_001_1672, w_000_1516, w_000_149);
  nand2 I001_1673(w_001_1673, w_000_1320, w_000_816);
  not1 I001_1674(w_001_1674, w_000_1295);
  or2  I001_1675(w_001_1675, w_000_1321, w_000_620);
  not1 I001_1676(w_001_1676, w_000_1012);
  not1 I001_1677(w_001_1677, w_000_1177);
  or2  I001_1680(w_001_1680, w_000_1156, w_000_1518);
  nand2 I001_1681(w_001_1681, w_000_1216, w_000_1185);
  and2 I001_1682(w_001_1682, w_000_381, w_000_1349);
  nand2 I001_1683(w_001_1683, w_000_590, w_000_980);
  or2  I001_1684(w_001_1684, w_000_1091, w_000_391);
  or2  I001_1685(w_001_1685, w_000_1519, w_000_1520);
  or2  I001_1687(w_001_1687, w_000_1287, w_000_211);
  nand2 I001_1688(w_001_1688, w_000_464, w_000_310);
  and2 I001_1689(w_001_1689, w_000_1521, w_000_931);
  or2  I002_000(w_002_000, w_001_1533, w_001_1655);
  not1 I002_001(w_002_001, w_001_388);
  nand2 I002_002(w_002_002, w_000_978, w_001_546);
  or2  I002_003(w_002_003, w_001_951, w_000_1522);
  and2 I002_004(w_002_004, w_001_868, w_001_884);
  nand2 I002_005(w_002_005, w_001_010, w_001_949);
  and2 I002_006(w_002_006, w_001_194, w_000_1112);
  nand2 I002_007(w_002_007, w_001_1120, w_000_1096);
  and2 I002_008(w_002_008, w_001_1260, w_001_617);
  not1 I002_009(w_002_009, w_000_408);
  not1 I002_010(w_002_010, w_001_429);
  not1 I002_011(w_002_011, w_000_1297);
  and2 I002_012(w_002_012, w_000_728, w_001_474);
  not1 I002_013(w_002_013, w_000_286);
  nand2 I002_014(w_002_014, w_000_856, w_001_604);
  nand2 I002_015(w_002_015, w_001_1402, w_001_1236);
  nand2 I002_016(w_002_016, w_000_427, w_000_1494);
  nand2 I002_017(w_002_017, w_000_604, w_000_073);
  nand2 I002_018(w_002_018, w_000_1523, w_001_250);
  nand2 I002_019(w_002_019, w_000_766, w_001_1278);
  or2  I002_020(w_002_020, w_000_155, w_001_671);
  nand2 I002_021(w_002_021, w_001_399, w_001_1316);
  nand2 I002_022(w_002_022, w_000_1004, w_000_721);
  nand2 I002_023(w_002_023, w_001_365, w_001_040);
  or2  I002_025(w_002_025, w_000_337, w_001_589);
  and2 I002_026(w_002_026, w_000_1005, w_001_1622);
  or2  I002_027(w_002_027, w_000_1215, w_000_451);
  nand2 I002_028(w_002_028, w_001_1583, w_000_829);
  and2 I002_029(w_002_029, w_001_1282, w_000_194);
  and2 I002_030(w_002_030, w_001_721, w_001_1382);
  not1 I002_031(w_002_031, w_000_1051);
  and2 I002_032(w_002_032, w_001_1640, w_000_062);
  not1 I002_033(w_002_033, w_001_036);
  nand2 I002_034(w_002_034, w_001_1603, w_001_1280);
  not1 I002_035(w_002_035, w_000_1215);
  not1 I002_036(w_002_036, w_001_182);
  or2  I002_037(w_002_037, w_001_1246, w_000_994);
  nand2 I002_038(w_002_038, w_001_1255, w_001_843);
  or2  I002_039(w_002_039, w_000_1524, w_000_189);
  nand2 I002_040(w_002_040, w_000_835, w_000_1525);
  not1 I002_041(w_002_041, w_001_1459);
  or2  I002_042(w_002_042, w_001_256, w_001_1683);
  and2 I002_043(w_002_043, w_000_1526, w_000_1515);
  or2  I002_044(w_002_044, w_000_509, w_000_883);
  and2 I002_045(w_002_045, w_001_078, w_001_610);
  not1 I002_046(w_002_046, w_000_799);
  or2  I002_047(w_002_047, w_000_1527, w_000_1201);
  and2 I002_048(w_002_048, w_001_660, w_001_1555);
  not1 I002_049(w_002_049, w_000_1528);
  nand2 I002_050(w_002_050, w_000_1497, w_001_697);
  not1 I002_051(w_002_051, w_001_1559);
  not1 I002_052(w_002_052, w_000_1529);
  nand2 I002_053(w_002_053, w_000_145, w_001_010);
  or2  I002_054(w_002_054, w_000_1200, w_001_036);
  and2 I002_055(w_002_055, w_000_1530, w_001_1227);
  nand2 I002_056(w_002_056, w_000_537, w_001_1332);
  and2 I002_057(w_002_057, w_001_829, w_001_1563);
  nand2 I002_058(w_002_058, w_000_1122, w_001_770);
  or2  I002_059(w_002_059, w_001_707, w_000_1022);
  or2  I002_060(w_002_060, w_001_1115, w_001_681);
  or2  I002_061(w_002_061, w_001_1247, w_000_1205);
  not1 I002_062(w_002_062, w_001_947);
  and2 I002_063(w_002_063, w_001_632, w_000_056);
  or2  I002_064(w_002_064, w_000_1531, w_001_142);
  or2  I002_065(w_002_065, w_000_1265, w_001_137);
  and2 I002_066(w_002_066, w_001_1202, w_001_1205);
  or2  I002_067(w_002_067, w_001_196, w_000_328);
  or2  I002_068(w_002_068, w_000_1532, w_000_1533);
  or2  I002_069(w_002_069, w_000_977, w_001_264);
  or2  I002_070(w_002_070, w_000_1142, w_001_1275);
  or2  I002_071(w_002_071, w_000_1022, w_000_101);
  or2  I002_072(w_002_072, w_000_1534, w_001_267);
  and2 I002_073(w_002_073, w_000_1226, w_000_583);
  nand2 I002_074(w_002_074, w_001_1213, w_000_287);
  nand2 I002_075(w_002_075, w_001_667, w_000_1146);
  and2 I002_076(w_002_076, w_000_777, w_000_127);
  and2 I002_077(w_002_077, w_001_1281, w_000_1317);
  nand2 I002_078(w_002_078, w_000_543, w_000_1031);
  nand2 I002_079(w_002_079, w_000_104, w_001_1412);
  nand2 I002_080(w_002_080, w_000_1035, w_000_441);
  nand2 I002_081(w_002_081, w_000_1535, w_000_284);
  or2  I002_082(w_002_082, w_000_702, w_000_053);
  or2  I002_083(w_002_083, w_000_116, w_001_229);
  not1 I002_084(w_002_084, w_000_857);
  or2  I002_085(w_002_085, w_000_1536, w_000_254);
  and2 I002_086(w_002_086, w_000_018, w_001_178);
  or2  I002_087(w_002_087, w_000_619, w_000_1240);
  not1 I002_088(w_002_088, w_001_186);
  nand2 I002_089(w_002_089, w_001_931, w_001_1102);
  and2 I002_090(w_002_090, w_001_1571, w_001_1088);
  or2  I002_091(w_002_091, w_001_255, w_000_1401);
  not1 I002_092(w_002_092, w_001_1655);
  not1 I002_093(w_002_093, w_001_1673);
  not1 I002_094(w_002_094, w_001_1079);
  not1 I002_095(w_002_095, w_001_159);
  not1 I002_096(w_002_096, w_001_1582);
  not1 I002_097(w_002_097, w_000_984);
  or2  I002_098(w_002_098, w_001_086, w_000_584);
  or2  I002_099(w_002_099, w_001_1673, w_000_1411);
  not1 I002_100(w_002_100, w_001_812);
  and2 I002_101(w_002_101, w_000_468, w_001_701);
  or2  I002_102(w_002_102, w_001_644, w_000_151);
  nand2 I002_103(w_002_103, w_000_1293, w_000_018);
  nand2 I002_104(w_002_104, w_000_1002, w_001_257);
  or2  I002_105(w_002_105, w_001_842, w_000_256);
  nand2 I002_106(w_002_106, w_001_1667, w_001_1630);
  and2 I002_107(w_002_107, w_000_918, w_000_385);
  nand2 I002_108(w_002_108, w_001_000, w_001_070);
  or2  I002_109(w_002_109, w_001_506, w_000_1537);
  and2 I002_110(w_002_110, w_001_276, w_001_016);
  or2  I002_111(w_002_111, w_000_1538, w_001_1474);
  not1 I002_112(w_002_112, w_000_1347);
  or2  I002_113(w_002_113, w_000_977, w_001_1130);
  nand2 I002_114(w_002_114, w_001_1515, w_000_1287);
  or2  I002_115(w_002_115, w_000_1539, w_000_417);
  nand2 I002_116(w_002_116, w_000_512, w_001_681);
  and2 I002_117(w_002_117, w_000_740, w_000_1346);
  or2  I002_118(w_002_118, w_001_821, w_001_700);
  and2 I002_119(w_002_119, w_001_484, w_000_498);
  not1 I002_120(w_002_120, w_001_1288);
  or2  I002_121(w_002_121, w_000_927, w_000_206);
  and2 I002_122(w_002_122, w_000_975, w_001_024);
  nand2 I002_123(w_002_123, w_000_1057, w_000_1540);
  or2  I002_124(w_002_124, w_000_1541, w_001_1111);
  and2 I002_125(w_002_125, w_000_1542, w_001_983);
  nand2 I002_126(w_002_126, w_001_1482, w_001_604);
  not1 I002_127(w_002_127, w_000_920);
  or2  I002_128(w_002_128, w_000_1478, w_001_272);
  or2  I002_129(w_002_129, w_000_296, w_001_1238);
  not1 I002_130(w_002_130, w_001_1559);
  nand2 I002_131(w_002_131, w_001_1227, w_000_1038);
  nand2 I002_132(w_002_132, w_001_1202, w_000_1028);
  or2  I002_133(w_002_133, w_001_510, w_001_892);
  and2 I002_134(w_002_134, w_001_164, w_001_746);
  nand2 I002_135(w_002_135, w_000_1018, w_000_366);
  nand2 I002_136(w_002_136, w_001_267, w_001_1662);
  and2 I002_137(w_002_137, w_000_1543, w_001_595);
  and2 I002_138(w_002_138, w_001_640, w_000_943);
  and2 I002_139(w_002_139, w_001_1231, w_001_1198);
  nand2 I002_140(w_002_140, w_001_460, w_001_1253);
  not1 I002_141(w_002_141, w_000_1027);
  and2 I002_142(w_002_142, w_001_056, w_001_134);
  nand2 I002_143(w_002_143, w_000_1487, w_001_099);
  and2 I002_144(w_002_144, w_001_736, w_000_886);
  and2 I002_145(w_002_145, w_000_181, w_000_1544);
  and2 I002_146(w_002_146, w_001_876, w_001_1147);
  and2 I002_147(w_002_147, w_001_752, w_000_1161);
  nand2 I002_148(w_002_148, w_001_244, w_001_1362);
  or2  I002_149(w_002_149, w_000_627, w_000_1545);
  and2 I002_150(w_002_150, w_000_1227, w_000_449);
  or2  I002_151(w_002_151, w_000_1546, w_000_980);
  or2  I002_152(w_002_152, w_001_1260, w_000_650);
  nand2 I002_153(w_002_153, w_000_1529, w_001_1233);
  nand2 I002_154(w_002_154, w_000_704, w_001_224);
  not1 I002_155(w_002_155, w_000_156);
  or2  I002_156(w_002_156, w_000_364, w_001_009);
  nand2 I002_157(w_002_157, w_001_458, w_000_901);
  or2  I002_158(w_002_158, w_001_234, w_001_522);
  not1 I002_159(w_002_159, w_001_1524);
  or2  I002_160(w_002_160, w_001_1054, w_000_1547);
  or2  I002_161(w_002_161, w_000_660, w_000_686);
  nand2 I002_162(w_002_162, w_001_1195, w_000_469);
  nand2 I002_163(w_002_163, w_000_830, w_001_663);
  and2 I002_164(w_002_164, w_001_227, w_000_1078);
  nand2 I002_165(w_002_165, w_001_1600, w_001_202);
  or2  I002_166(w_002_166, w_000_573, w_001_1422);
  not1 I002_167(w_002_167, w_000_236);
  not1 I002_168(w_002_168, w_000_923);
  or2  I002_169(w_002_169, w_001_470, w_000_743);
  or2  I002_170(w_002_170, w_000_1548, w_000_403);
  not1 I002_171(w_002_171, w_000_320);
  and2 I002_172(w_002_172, w_000_823, w_001_939);
  and2 I002_173(w_002_173, w_001_416, w_000_112);
  nand2 I002_174(w_002_174, w_000_290, w_001_095);
  or2  I002_175(w_002_175, w_001_1060, w_000_1549);
  not1 I002_176(w_002_176, w_000_1068);
  nand2 I002_177(w_002_177, w_000_993, w_000_992);
  nand2 I002_178(w_002_178, w_000_1550, w_001_168);
  and2 I002_179(w_002_179, w_000_1149, w_000_1551);
  or2  I002_180(w_002_180, w_001_364, w_000_983);
  not1 I002_181(w_002_181, w_001_768);
  nand2 I002_182(w_002_182, w_001_138, w_000_816);
  not1 I002_183(w_002_183, w_000_236);
  not1 I002_184(w_002_184, w_001_1581);
  not1 I002_185(w_002_185, w_001_493);
  not1 I002_186(w_002_186, w_001_1516);
  and2 I002_187(w_002_187, w_001_187, w_000_128);
  and2 I002_188(w_002_188, w_001_1563, w_000_1552);
  not1 I002_189(w_002_189, w_001_631);
  nand2 I002_190(w_002_190, w_000_1474, w_001_224);
  not1 I002_191(w_002_191, w_000_959);
  not1 I002_192(w_002_192, w_000_634);
  and2 I002_193(w_002_193, w_000_949, w_001_872);
  and2 I002_194(w_002_194, w_001_1484, w_000_1402);
  not1 I002_195(w_002_195, w_000_1531);
  not1 I002_196(w_002_196, w_001_023);
  not1 I002_197(w_002_197, w_001_1522);
  or2  I002_198(w_002_198, w_000_1157, w_000_908);
  or2  I002_199(w_002_199, w_000_466, w_000_1449);
  not1 I002_200(w_002_200, w_000_613);
  and2 I002_201(w_002_201, w_001_270, w_000_260);
  nand2 I002_202(w_002_202, w_000_360, w_000_1127);
  and2 I002_203(w_002_203, w_001_053, w_001_1104);
  nand2 I002_204(w_002_204, w_000_627, w_000_593);
  and2 I002_205(w_002_205, w_000_1553, w_001_363);
  nand2 I002_206(w_002_206, w_000_164, w_001_592);
  or2  I002_207(w_002_207, w_001_1220, w_001_941);
  and2 I002_208(w_002_208, w_000_821, w_000_1448);
  and2 I002_209(w_002_209, w_000_529, w_001_1271);
  not1 I002_210(w_002_210, w_000_803);
  or2  I002_211(w_002_211, w_001_1396, w_001_195);
  or2  I002_212(w_002_212, w_000_600, w_000_588);
  and2 I002_213(w_002_213, w_001_1181, w_001_542);
  or2  I002_214(w_002_214, w_000_1483, w_001_205);
  or2  I002_215(w_002_215, w_001_1343, w_001_261);
  or2  I002_216(w_002_216, w_001_194, w_001_131);
  nand2 I002_217(w_002_217, w_000_224, w_000_1333);
  not1 I002_218(w_002_218, w_001_1007);
  not1 I002_219(w_002_219, w_000_1554);
  nand2 I002_220(w_002_220, w_001_1129, w_000_1202);
  not1 I002_221(w_002_221, w_001_1037);
  nand2 I002_222(w_002_222, w_000_1555, w_000_1307);
  and2 I002_223(w_002_223, w_001_1532, w_001_445);
  nand2 I002_224(w_002_224, w_000_1484, w_001_319);
  and2 I002_225(w_002_225, w_000_429, w_000_668);
  nand2 I002_226(w_002_226, w_000_264, w_000_927);
  or2  I002_227(w_002_227, w_001_129, w_001_122);
  nand2 I002_228(w_002_228, w_000_1556, w_001_1098);
  nand2 I002_229(w_002_229, w_001_1659, w_000_1476);
  and2 I002_230(w_002_230, w_001_233, w_000_1557);
  not1 I002_231(w_002_231, w_001_1403);
  nand2 I002_232(w_002_232, w_001_071, w_000_439);
  nand2 I002_233(w_002_233, w_001_028, w_000_1558);
  and2 I002_234(w_002_234, w_001_050, w_001_223);
  and2 I002_235(w_002_235, w_000_1363, w_001_446);
  not1 I002_236(w_002_236, w_001_274);
  not1 I002_237(w_002_237, w_001_197);
  nand2 I002_238(w_002_238, w_000_439, w_000_1537);
  not1 I002_239(w_002_239, w_001_1609);
  or2  I002_240(w_002_240, w_000_296, w_000_312);
  or2  I002_241(w_002_241, w_000_512, w_000_1559);
  nand2 I002_242(w_002_242, w_000_1458, w_000_1560);
  or2  I002_243(w_002_243, w_000_848, w_001_194);
  not1 I002_244(w_002_244, w_000_082);
  or2  I002_245(w_002_245, w_000_873, w_001_1447);
  and2 I002_246(w_002_246, w_000_1056, w_001_478);
  or2  I002_247(w_002_247, w_001_791, w_000_1141);
  nand2 I002_248(w_002_248, w_000_731, w_001_1444);
  or2  I002_249(w_002_249, w_001_1270, w_000_1561);
  not1 I002_250(w_002_250, w_001_193);
  and2 I002_251(w_002_251, w_001_275, w_000_1429);
  or2  I002_252(w_002_252, w_001_877, w_001_226);
  or2  I002_253(w_002_253, w_000_394, w_000_257);
  or2  I002_255(w_002_255, w_000_1203, w_000_723);
  or2  I002_256(w_002_256, w_000_1032, w_001_1124);
  or2  I002_257(w_002_257, w_000_643, w_001_394);
  or2  I002_258(w_002_258, w_000_425, w_000_599);
  or2  I002_259(w_002_259, w_001_1565, w_000_1563);
  not1 I002_260(w_002_260, w_001_1058);
  and2 I002_261(w_002_261, w_000_1169, w_001_1138);
  or2  I002_262(w_002_262, w_001_213, w_000_567);
  or2  I002_263(w_002_263, w_000_043, w_001_1290);
  nand2 I002_264(w_002_264, w_000_1564, w_000_734);
  or2  I002_265(w_002_265, w_000_1565, w_001_1057);
  not1 I002_266(w_002_266, w_001_1339);
  and2 I002_267(w_002_267, w_000_398, w_000_223);
  nand2 I002_268(w_002_268, w_001_1361, w_000_348);
  nand2 I002_269(w_002_269, w_001_915, w_000_689);
  nand2 I002_270(w_002_270, w_001_289, w_000_1375);
  nand2 I002_271(w_002_271, w_000_461, w_000_932);
  not1 I002_272(w_002_272, w_001_299);
  and2 I002_273(w_002_273, w_000_1566, w_000_1567);
  nand2 I002_274(w_002_274, w_000_150, w_000_1568);
  nand2 I002_275(w_002_275, w_001_141, w_000_1190);
  or2  I002_276(w_002_276, w_001_189, w_000_1569);
  not1 I002_277(w_002_277, w_000_1390);
  or2  I002_278(w_002_278, w_000_1570, w_001_1112);
  not1 I002_280(w_002_280, w_001_1486);
  nand2 I002_281(w_002_281, w_000_1571, w_001_876);
  and2 I002_282(w_002_282, w_001_1092, w_001_894);
  not1 I002_283(w_002_283, w_001_303);
  or2  I002_284(w_002_284, w_000_1023, w_000_1572);
  or2  I002_285(w_002_285, w_000_175, w_001_115);
  and2 I002_286(w_002_286, w_001_113, w_001_1191);
  not1 I002_287(w_002_287, w_001_677);
  or2  I002_288(w_002_288, w_001_947, w_000_1260);
  nand2 I002_289(w_002_289, w_001_352, w_000_1540);
  not1 I002_290(w_002_290, w_001_153);
  and2 I002_291(w_002_291, w_001_867, w_000_1325);
  and2 I002_292(w_002_292, w_000_1573, w_000_459);
  and2 I002_293(w_002_293, w_001_615, w_000_514);
  or2  I002_294(w_002_294, w_001_1544, w_000_682);
  nand2 I002_295(w_002_295, w_000_1574, w_000_340);
  or2  I002_297(w_002_297, w_001_075, w_001_714);
  not1 I002_298(w_002_298, w_001_391);
  nand2 I002_299(w_002_299, w_001_243, w_001_1238);
  nand2 I002_300(w_002_300, w_000_1576, w_001_1327);
  not1 I002_301(w_002_301, w_000_871);
  and2 I002_302(w_002_302, w_001_1362, w_001_1241);
  and2 I002_303(w_002_303, w_001_240, w_000_1577);
  or2  I002_304(w_002_304, w_001_232, w_000_1578);
  or2  I002_305(w_002_305, w_001_160, w_000_802);
  nand2 I002_306(w_002_306, w_001_040, w_000_125);
  not1 I002_307(w_002_307, w_000_1452);
  and2 I002_308(w_002_308, w_000_323, w_001_1607);
  or2  I002_309(w_002_309, w_000_1201, w_001_847);
  or2  I002_310(w_002_310, w_001_1046, w_000_1284);
  and2 I002_311(w_002_311, w_000_1053, w_001_539);
  or2  I002_312(w_002_312, w_001_1341, w_000_026);
  or2  I002_313(w_002_313, w_001_504, w_001_1147);
  and2 I002_314(w_002_314, w_000_1579, w_000_1257);
  nand2 I002_315(w_002_315, w_001_489, w_000_831);
  and2 I002_316(w_002_316, w_001_1060, w_000_1027);
  or2  I002_317(w_002_317, w_000_1543, w_000_944);
  not1 I002_318(w_002_318, w_000_1580);
  nand2 I002_319(w_002_319, w_000_036, w_000_1091);
  and2 I002_320(w_002_320, w_000_238, w_000_1140);
  not1 I002_321(w_002_321, w_000_397);
  or2  I002_322(w_002_322, w_000_1238, w_001_981);
  not1 I002_323(w_002_323, w_000_393);
  and2 I002_324(w_002_324, w_001_1090, w_000_464);
  or2  I002_325(w_002_325, w_000_898, w_001_1020);
  or2  I002_326(w_002_326, w_001_1408, w_001_293);
  and2 I002_327(w_002_327, w_001_531, w_000_457);
  or2  I002_328(w_002_328, w_001_1206, w_000_427);
  and2 I002_329(w_002_329, w_001_070, w_000_825);
  or2  I002_330(w_002_330, w_000_098, w_000_1449);
  not1 I002_331(w_002_331, w_001_811);
  and2 I002_332(w_002_332, w_000_1581, w_001_1203);
  nand2 I002_333(w_002_333, w_001_1496, w_001_1632);
  and2 I002_334(w_002_334, w_000_442, w_001_613);
  and2 I002_335(w_002_335, w_000_1392, w_001_391);
  and2 I002_336(w_002_336, w_001_1217, w_001_1198);
  not1 I002_338(w_002_338, w_000_1583);
  not1 I002_339(w_002_339, w_000_896);
  or2  I002_340(w_002_340, w_001_744, w_001_235);
  and2 I002_341(w_002_341, w_001_677, w_000_074);
  not1 I002_342(w_002_342, w_000_1466);
  nand2 I002_343(w_002_343, w_001_618, w_000_558);
  nand2 I002_344(w_002_344, w_000_226, w_001_783);
  and2 I002_345(w_002_345, w_001_594, w_000_912);
  and2 I002_346(w_002_346, w_000_1584, w_001_445);
  and2 I002_347(w_002_347, w_000_681, w_001_013);
  not1 I002_348(w_002_348, w_001_087);
  and2 I002_349(w_002_349, w_001_1595, w_001_754);
  or2  I002_350(w_002_350, w_000_1313, w_001_192);
  nand2 I002_351(w_002_351, w_000_1018, w_001_885);
  and2 I002_352(w_002_352, w_001_149, w_000_1504);
  or2  I002_353(w_002_353, w_001_259, w_000_264);
  not1 I002_354(w_002_354, w_001_319);
  or2  I002_355(w_002_355, w_000_449, w_001_175);
  and2 I002_356(w_002_356, w_001_929, w_000_1585);
  not1 I002_357(w_002_357, w_001_179);
  or2  I002_358(w_002_358, w_001_887, w_000_354);
  nand2 I002_359(w_002_359, w_000_504, w_001_350);
  or2  I002_360(w_002_360, w_001_651, w_001_1337);
  not1 I002_361(w_002_361, w_000_1586);
  not1 I002_363(w_002_363, w_001_785);
  or2  I002_365(w_002_365, w_000_985, w_001_386);
  or2  I002_366(w_002_366, w_001_890, w_000_245);
  and2 I002_367(w_002_367, w_001_897, w_001_002);
  nand2 I002_368(w_002_368, w_000_1587, w_000_682);
  and2 I002_369(w_002_369, w_000_538, w_000_1588);
  nand2 I002_370(w_002_370, w_000_032, w_000_293);
  not1 I002_371(w_002_371, w_001_325);
  and2 I002_372(w_002_372, w_001_1064, w_001_1160);
  not1 I002_373(w_002_373, w_001_1406);
  not1 I002_374(w_002_374, w_001_655);
  not1 I002_375(w_002_375, w_001_1538);
  and2 I002_376(w_002_376, w_000_396, w_000_045);
  not1 I002_377(w_002_377, w_000_1015);
  not1 I002_378(w_002_378, w_001_1098);
  nand2 I002_379(w_002_379, w_000_1589, w_001_1261);
  or2  I002_380(w_002_380, w_001_878, w_001_810);
  nand2 I002_381(w_002_381, w_001_412, w_001_154);
  nand2 I002_382(w_002_382, w_000_600, w_000_342);
  and2 I002_383(w_002_383, w_001_1090, w_000_570);
  and2 I002_384(w_002_384, w_001_1585, w_001_950);
  nand2 I002_385(w_002_385, w_000_1590, w_001_051);
  not1 I002_386(w_002_386, w_000_1205);
  and2 I002_387(w_002_387, w_001_367, w_001_476);
  nand2 I002_388(w_002_388, w_000_982, w_000_1128);
  not1 I002_389(w_002_389, w_001_132);
  not1 I002_390(w_002_390, w_000_912);
  or2  I002_391(w_002_391, w_000_313, w_000_735);
  and2 I002_392(w_002_392, w_000_1591, w_000_1475);
  not1 I002_393(w_002_393, w_001_1437);
  not1 I002_394(w_002_394, w_000_277);
  nand2 I002_395(w_002_395, w_000_1157, w_001_005);
  or2  I002_396(w_002_396, w_000_1592, w_000_532);
  nand2 I002_397(w_002_397, w_000_1219, w_001_049);
  and2 I002_398(w_002_398, w_001_362, w_000_1593);
  not1 I002_399(w_002_399, w_000_1594);
  and2 I002_400(w_002_400, w_001_657, w_001_762);
  nand2 I002_401(w_002_401, w_000_1392, w_000_1530);
  or2  I002_402(w_002_402, w_000_1595, w_000_1596);
  nand2 I002_403(w_002_403, w_000_644, w_000_1537);
  nand2 I002_404(w_002_404, w_001_248, w_001_922);
  and2 I002_405(w_002_405, w_001_1259, w_000_1226);
  not1 I002_406(w_002_406, w_000_551);
  and2 I002_407(w_002_407, w_001_1666, w_001_143);
  not1 I002_408(w_002_408, w_000_1597);
  nand2 I002_409(w_002_409, w_000_1598, w_001_1604);
  and2 I002_410(w_002_410, w_000_248, w_001_631);
  and2 I002_411(w_002_411, w_000_569, w_001_491);
  or2  I002_412(w_002_412, w_001_060, w_001_181);
  and2 I002_413(w_002_413, w_001_1084, w_000_1000);
  not1 I002_414(w_002_414, w_000_1496);
  not1 I002_416(w_002_416, w_001_012);
  nand2 I002_417(w_002_417, w_001_302, w_000_1242);
  not1 I002_418(w_002_418, w_000_163);
  not1 I002_419(w_002_419, w_001_046);
  or2  I002_420(w_002_420, w_001_1207, w_000_1520);
  and2 I002_421(w_002_421, w_000_1012, w_000_965);
  and2 I002_422(w_002_422, w_000_1125, w_000_1442);
  or2  I002_423(w_002_423, w_000_876, w_000_1599);
  nand2 I002_424(w_002_424, w_001_307, w_001_967);
  nand2 I002_425(w_002_425, w_000_1130, w_001_041);
  not1 I002_426(w_002_426, w_000_445);
  or2  I002_427(w_002_427, w_000_317, w_001_1403);
  or2  I002_428(w_002_428, w_001_720, w_000_1490);
  or2  I002_429(w_002_429, w_000_932, w_000_1600);
  and2 I002_430(w_002_430, w_000_1495, w_000_633);
  and2 I002_431(w_002_431, w_001_1600, w_000_1405);
  not1 I002_432(w_002_432, w_001_1447);
  and2 I002_433(w_002_433, w_000_244, w_001_1076);
  or2  I002_434(w_002_434, w_000_831, w_000_144);
  nand2 I002_435(w_002_435, w_000_1601, w_001_669);
  not1 I002_436(w_002_436, w_001_470);
  not1 I002_437(w_002_437, w_000_1602);
  not1 I002_438(w_002_438, w_001_120);
  and2 I002_439(w_002_439, w_000_1122, w_001_190);
  nand2 I002_440(w_002_440, w_000_181, w_001_1688);
  not1 I002_441(w_002_441, w_000_249);
  or2  I002_442(w_002_442, w_001_492, w_001_1003);
  and2 I002_443(w_002_443, w_001_1456, w_001_247);
  nand2 I002_444(w_002_444, w_001_1015, w_001_457);
  not1 I002_445(w_002_445, w_001_267);
  not1 I002_446(w_002_446, w_001_051);
  nand2 I002_447(w_002_447, w_001_692, w_000_1603);
  and2 I002_448(w_002_448, w_000_1604, w_000_858);
  and2 I002_449(w_002_449, w_001_012, w_001_1198);
  not1 I002_450(w_002_450, w_000_654);
  and2 I002_451(w_002_451, w_001_1062, w_001_772);
  or2  I002_452(w_002_452, w_000_362, w_000_995);
  and2 I002_453(w_002_453, w_001_1088, w_000_1605);
  or2  I002_454(w_002_454, w_000_1606, w_001_492);
  and2 I002_456(w_002_456, w_001_113, w_001_1145);
  or2  I002_457(w_002_457, w_001_902, w_001_1454);
  nand2 I002_458(w_002_458, w_001_183, w_001_1643);
  not1 I002_459(w_002_459, w_000_1607);
  nand2 I002_460(w_002_460, w_000_1438, w_000_134);
  nand2 I002_461(w_002_461, w_001_978, w_000_1608);
  or2  I002_462(w_002_462, w_000_374, w_001_1106);
  or2  I002_463(w_002_463, w_000_603, w_001_1135);
  not1 I002_464(w_002_464, w_000_590);
  or2  I002_465(w_002_465, w_001_1125, w_000_759);
  nand2 I002_466(w_002_466, w_000_404, w_000_1609);
  not1 I002_467(w_002_467, w_000_296);
  or2  I002_468(w_002_468, w_001_1627, w_001_453);
  and2 I002_469(w_002_469, w_000_828, w_001_596);
  or2  I002_470(w_002_470, w_000_1199, w_000_1129);
  or2  I002_471(w_002_471, w_001_071, w_000_078);
  and2 I002_472(w_002_472, w_001_1189, w_000_1610);
  or2  I002_473(w_002_473, w_000_1611, w_001_097);
  and2 I002_474(w_002_474, w_001_780, w_001_894);
  not1 I002_475(w_002_475, w_001_032);
  not1 I002_476(w_002_476, w_001_628);
  nand2 I002_477(w_002_477, w_001_180, w_000_1504);
  or2  I002_478(w_002_478, w_001_1576, w_000_917);
  and2 I002_479(w_002_479, w_001_107, w_000_1342);
  and2 I002_480(w_002_480, w_001_000, w_000_200);
  nand2 I002_481(w_002_481, w_001_980, w_000_271);
  not1 I002_482(w_002_482, w_000_656);
  and2 I002_483(w_002_483, w_001_1636, w_000_1590);
  and2 I002_484(w_002_484, w_000_1094, w_000_1612);
  not1 I002_485(w_002_485, w_000_1088);
  nand2 I002_486(w_002_486, w_001_1195, w_001_197);
  and2 I002_487(w_002_487, w_000_1613, w_000_130);
  nand2 I002_488(w_002_488, w_001_1463, w_001_102);
  or2  I002_489(w_002_489, w_001_800, w_000_286);
  or2  I002_490(w_002_490, w_000_228, w_001_108);
  nand2 I002_491(w_002_491, w_001_1617, w_001_061);
  or2  I002_492(w_002_492, w_000_564, w_001_672);
  not1 I002_493(w_002_493, w_001_602);
  not1 I002_494(w_002_494, w_001_1085);
  or2  I002_495(w_002_495, w_000_548, w_000_1614);
  or2  I002_496(w_002_496, w_000_463, w_001_116);
  and2 I002_497(w_002_497, w_001_345, w_001_555);
  and2 I002_498(w_002_498, w_001_524, w_001_000);
  not1 I002_499(w_002_499, w_000_255);
  nand2 I002_500(w_002_500, w_000_1017, w_000_1615);
  nand2 I002_501(w_002_501, w_001_977, w_000_259);
  or2  I002_502(w_002_502, w_000_273, w_001_142);
  and2 I002_503(w_002_503, w_000_1616, w_000_1504);
  not1 I002_504(w_002_504, w_000_059);
  not1 I002_505(w_002_505, w_001_936);
  nand2 I002_506(w_002_506, w_001_870, w_001_828);
  or2  I002_507(w_002_507, w_001_197, w_001_480);
  and2 I002_508(w_002_508, w_000_1457, w_000_1153);
  nand2 I002_509(w_002_509, w_001_1426, w_000_351);
  nand2 I002_510(w_002_510, w_000_652, w_001_040);
  not1 I002_511(w_002_511, w_001_452);
  and2 I002_512(w_002_512, w_000_1388, w_000_1617);
  not1 I002_513(w_002_513, w_001_746);
  nand2 I002_514(w_002_514, w_001_1296, w_000_065);
  and2 I002_515(w_002_515, w_000_1522, w_001_219);
  or2  I002_516(w_002_516, w_000_1618, w_001_1251);
  and2 I002_517(w_002_517, w_000_1619, w_000_1620);
  nand2 I002_519(w_002_519, w_000_472, w_001_148);
  or2  I002_521(w_002_521, w_001_542, w_001_810);
  nand2 I002_522(w_002_522, w_001_685, w_000_910);
  not1 I002_523(w_002_523, w_000_1260);
  not1 I002_524(w_002_524, w_001_124);
  not1 I002_525(w_002_525, w_001_548);
  not1 I002_526(w_002_526, w_000_1434);
  nand2 I002_527(w_002_527, w_001_016, w_001_038);
  and2 I002_528(w_002_528, w_000_888, w_000_1507);
  not1 I002_529(w_002_529, w_001_1133);
  and2 I002_530(w_002_530, w_000_1472, w_001_1500);
  nand2 I002_531(w_002_531, w_000_1188, w_001_974);
  nand2 I002_532(w_002_532, w_001_460, w_001_1020);
  not1 I002_533(w_002_533, w_001_806);
  or2  I002_534(w_002_534, w_000_822, w_001_1366);
  not1 I002_535(w_002_535, w_001_606);
  and2 I002_536(w_002_536, w_000_592, w_001_1447);
  or2  I002_537(w_002_537, w_001_1272, w_000_321);
  nand2 I002_538(w_002_538, w_000_1509, w_000_1220);
  or2  I002_539(w_002_539, w_001_032, w_000_197);
  nand2 I002_540(w_002_540, w_001_1355, w_000_1375);
  or2  I002_541(w_002_541, w_001_1093, w_001_150);
  nand2 I002_542(w_002_542, w_000_155, w_000_725);
  not1 I002_543(w_002_543, w_001_1547);
  not1 I002_544(w_002_544, w_001_178);
  or2  I002_545(w_002_545, w_000_1621, w_001_1074);
  nand2 I002_546(w_002_546, w_001_1107, w_001_1314);
  not1 I002_547(w_002_547, w_000_1022);
  not1 I002_548(w_002_548, w_001_1551);
  and2 I002_549(w_002_549, w_000_1622, w_000_1623);
  nand2 I002_550(w_002_550, w_001_635, w_000_038);
  and2 I002_551(w_002_551, w_001_1264, w_000_1624);
  not1 I002_552(w_002_552, w_000_1625);
  or2  I002_553(w_002_553, w_000_1626, w_000_1607);
  and2 I002_554(w_002_554, w_001_1325, w_000_947);
  and2 I002_555(w_002_555, w_001_850, w_000_435);
  or2  I002_556(w_002_556, w_000_778, w_000_832);
  not1 I002_557(w_002_557, w_001_1222);
  not1 I002_558(w_002_558, w_000_838);
  not1 I002_559(w_002_559, w_000_040);
  and2 I002_560(w_002_560, w_000_1182, w_001_1639);
  and2 I002_561(w_002_561, w_000_1111, w_001_1570);
  nand2 I002_562(w_002_562, w_000_1598, w_000_1627);
  not1 I002_563(w_002_563, w_001_840);
  not1 I002_564(w_002_564, w_000_553);
  not1 I002_565(w_002_565, w_000_786);
  and2 I002_566(w_002_566, w_000_1086, w_001_1027);
  nand2 I002_567(w_002_567, w_001_1163, w_001_1633);
  and2 I002_568(w_002_568, w_001_1426, w_001_286);
  nand2 I002_569(w_002_569, w_001_384, w_000_1213);
  not1 I002_570(w_002_570, w_001_1279);
  and2 I002_571(w_002_571, w_001_445, w_000_476);
  and2 I002_572(w_002_572, w_000_1614, w_000_1050);
  or2  I002_573(w_002_573, w_001_429, w_000_527);
  or2  I002_574(w_002_574, w_001_512, w_001_818);
  not1 I002_575(w_002_575, w_000_1147);
  not1 I002_576(w_002_576, w_001_193);
  not1 I002_577(w_002_577, w_000_1521);
  or2  I002_578(w_002_578, w_001_849, w_000_343);
  or2  I002_579(w_002_579, w_001_787, w_001_451);
  nand2 I002_580(w_002_580, w_000_1504, w_001_1211);
  and2 I002_581(w_002_581, w_000_804, w_000_270);
  not1 I002_582(w_002_582, w_000_561);
  and2 I002_583(w_002_583, w_001_699, w_000_386);
  or2  I002_584(w_002_584, w_000_1628, w_000_854);
  or2  I002_585(w_002_585, w_000_1197, w_001_279);
  and2 I002_586(w_002_586, w_000_1083, w_001_226);
  nand2 I002_587(w_002_587, w_000_1128, w_000_1629);
  and2 I002_588(w_002_588, w_000_047, w_000_714);
  and2 I002_589(w_002_589, w_001_1570, w_001_175);
  and2 I002_590(w_002_590, w_000_821, w_000_202);
  nand2 I002_591(w_002_591, w_000_1630, w_000_1631);
  and2 I002_592(w_002_592, w_000_1271, w_001_700);
  and2 I002_593(w_002_593, w_000_1070, w_000_174);
  and2 I003_000(w_003_000, w_002_058, w_000_951);
  not1 I003_001(w_003_001, w_001_521);
  or2  I003_002(w_003_002, w_000_829, w_001_704);
  not1 I003_003(w_003_003, w_002_138);
  and2 I003_004(w_003_004, w_002_308, w_001_121);
  or2  I003_005(w_003_005, w_000_1632, w_000_1633);
  or2  I003_006(w_003_006, w_000_692, w_002_354);
  or2  I003_007(w_003_007, w_002_194, w_000_591);
  not1 I003_008(w_003_008, w_001_1112);
  nand2 I003_009(w_003_009, w_002_159, w_002_499);
  nand2 I003_010(w_003_010, w_002_177, w_002_325);
  not1 I003_011(w_003_011, w_001_1082);
  nand2 I003_012(w_003_012, w_002_363, w_002_487);
  not1 I003_013(w_003_013, w_002_126);
  or2  I003_014(w_003_014, w_001_475, w_001_020);
  nand2 I003_015(w_003_015, w_002_463, w_002_338);
  and2 I003_016(w_003_016, w_001_1226, w_001_007);
  or2  I003_017(w_003_017, w_000_185, w_000_879);
  nand2 I003_018(w_003_018, w_002_314, w_000_370);
  nand2 I003_019(w_003_019, w_002_022, w_002_145);
  not1 I003_020(w_003_020, w_001_1067);
  or2  I003_021(w_003_021, w_001_778, w_002_448);
  nand2 I003_022(w_003_022, w_001_1381, w_001_1159);
  nand2 I003_023(w_003_023, w_000_1166, w_001_1345);
  nand2 I003_024(w_003_024, w_001_224, w_000_171);
  not1 I003_025(w_003_025, w_000_893);
  or2  I003_026(w_003_026, w_000_1049, w_002_072);
  nand2 I003_027(w_003_027, w_002_303, w_002_349);
  or2  I003_028(w_003_028, w_001_797, w_002_405);
  not1 I003_029(w_003_029, w_001_1564);
  or2  I003_030(w_003_030, w_001_731, w_002_103);
  not1 I003_031(w_003_031, w_001_1274);
  or2  I003_032(w_003_032, w_000_164, w_002_102);
  not1 I003_033(w_003_033, w_000_1634);
  and2 I003_034(w_003_034, w_002_131, w_001_1107);
  or2  I003_035(w_003_035, w_002_541, w_002_220);
  or2  I003_036(w_003_036, w_002_508, w_001_1296);
  and2 I003_037(w_003_037, w_001_027, w_001_1259);
  or2  I003_038(w_003_038, w_000_885, w_000_688);
  not1 I003_039(w_003_039, w_001_1384);
  and2 I003_040(w_003_040, w_001_1129, w_000_400);
  not1 I003_041(w_003_041, w_000_1507);
  and2 I003_042(w_003_042, w_002_048, w_001_148);
  not1 I003_043(w_003_043, w_001_1251);
  nand2 I003_044(w_003_044, w_002_195, w_001_1400);
  or2  I003_045(w_003_045, w_001_214, w_002_042);
  and2 I003_046(w_003_046, w_001_1444, w_001_518);
  and2 I003_047(w_003_047, w_000_000, w_001_260);
  not1 I003_048(w_003_048, w_001_078);
  not1 I003_049(w_003_049, w_001_1356);
  and2 I003_050(w_003_050, w_000_1130, w_000_791);
  not1 I003_051(w_003_051, w_002_150);
  nand2 I003_052(w_003_052, w_002_061, w_000_046);
  or2  I003_053(w_003_053, w_000_1635, w_000_303);
  nand2 I003_054(w_003_054, w_002_180, w_002_050);
  or2  I003_055(w_003_055, w_002_015, w_002_122);
  nand2 I003_056(w_003_056, w_001_1260, w_002_343);
  nand2 I003_057(w_003_057, w_000_674, w_000_789);
  and2 I003_058(w_003_058, w_001_269, w_001_1685);
  nand2 I003_059(w_003_059, w_000_544, w_002_513);
  nand2 I003_060(w_003_060, w_001_103, w_002_438);
  not1 I003_061(w_003_061, w_000_1168);
  nand2 I003_062(w_003_062, w_000_1072, w_000_516);
  or2  I003_063(w_003_063, w_000_047, w_002_042);
  not1 I003_064(w_003_064, w_002_238);
  not1 I003_065(w_003_065, w_001_005);
  not1 I003_066(w_003_066, w_001_363);
  nand2 I003_067(w_003_067, w_002_319, w_002_340);
  not1 I003_068(w_003_068, w_000_1017);
  not1 I003_069(w_003_069, w_000_238);
  nand2 I003_070(w_003_070, w_000_762, w_002_459);
  not1 I003_071(w_003_071, w_000_385);
  not1 I003_072(w_003_072, w_002_428);
  and2 I003_073(w_003_073, w_002_448, w_000_1247);
  nand2 I003_074(w_003_074, w_002_085, w_000_1636);
  and2 I003_075(w_003_075, w_001_129, w_002_303);
  nand2 I003_076(w_003_076, w_002_220, w_002_119);
  nand2 I003_077(w_003_077, w_000_1476, w_000_1637);
  not1 I003_078(w_003_078, w_001_413);
  and2 I003_079(w_003_079, w_001_1435, w_000_1638);
  nand2 I003_080(w_003_080, w_002_292, w_001_155);
  or2  I003_081(w_003_081, w_002_023, w_002_065);
  not1 I003_082(w_003_082, w_002_368);
  or2  I003_083(w_003_083, w_002_128, w_002_032);
  or2  I003_084(w_003_084, w_000_1639, w_000_939);
  nand2 I003_085(w_003_085, w_002_164, w_000_358);
  and2 I003_086(w_003_086, w_001_239, w_001_1367);
  nand2 I003_087(w_003_087, w_002_334, w_000_048);
  or2  I003_088(w_003_088, w_000_465, w_001_922);
  nand2 I003_089(w_003_089, w_002_593, w_001_911);
  or2  I003_090(w_003_090, w_000_174, w_001_311);
  or2  I003_091(w_003_091, w_000_1234, w_001_612);
  or2  I003_092(w_003_092, w_002_010, w_000_1640);
  nand2 I003_093(w_003_093, w_000_144, w_002_111);
  and2 I003_094(w_003_094, w_002_189, w_002_539);
  or2  I003_095(w_003_095, w_001_1053, w_002_102);
  and2 I003_096(w_003_096, w_001_264, w_001_1654);
  or2  I003_097(w_003_097, w_002_163, w_000_774);
  nand2 I003_098(w_003_098, w_002_490, w_002_441);
  not1 I003_099(w_003_099, w_000_1641);
  not1 I003_100(w_003_100, w_002_130);
  not1 I003_101(w_003_101, w_000_454);
  nand2 I003_102(w_003_102, w_001_009, w_000_1237);
  not1 I003_103(w_003_103, w_000_1554);
  not1 I003_104(w_003_104, w_002_045);
  and2 I003_105(w_003_105, w_001_001, w_001_025);
  and2 I003_106(w_003_106, w_000_1470, w_001_1382);
  and2 I003_107(w_003_107, w_000_1086, w_001_1304);
  nand2 I003_108(w_003_108, w_002_278, w_002_140);
  or2  I003_109(w_003_109, w_002_191, w_000_054);
  nand2 I003_110(w_003_110, w_001_1608, w_000_1163);
  or2  I003_111(w_003_111, w_001_1688, w_002_508);
  not1 I003_112(w_003_112, w_000_863);
  and2 I003_113(w_003_113, w_001_245, w_002_090);
  nand2 I003_114(w_003_114, w_001_056, w_000_1642);
  or2  I003_115(w_003_115, w_002_068, w_002_580);
  or2  I003_116(w_003_116, w_002_041, w_001_1462);
  nand2 I003_117(w_003_117, w_002_383, w_002_218);
  not1 I003_118(w_003_118, w_001_1320);
  and2 I003_119(w_003_119, w_001_183, w_002_500);
  or2  I003_120(w_003_120, w_000_1184, w_002_285);
  nand2 I003_121(w_003_121, w_002_431, w_001_791);
  or2  I003_122(w_003_122, w_000_559, w_000_1258);
  not1 I003_123(w_003_123, w_001_1072);
  not1 I003_124(w_003_124, w_001_050);
  nand2 I003_125(w_003_125, w_000_1068, w_001_068);
  and2 I003_126(w_003_126, w_000_294, w_001_944);
  nand2 I003_127(w_003_127, w_002_481, w_001_162);
  and2 I003_128(w_003_128, w_001_1229, w_002_522);
  not1 I003_129(w_003_129, w_002_487);
  or2  I003_130(w_003_130, w_001_126, w_002_345);
  not1 I003_131(w_003_131, w_001_747);
  or2  I003_132(w_003_132, w_002_033, w_000_431);
  nand2 I003_133(w_003_133, w_001_1077, w_001_1298);
  and2 I003_134(w_003_134, w_001_131, w_001_861);
  nand2 I003_135(w_003_135, w_000_091, w_000_1643);
  or2  I003_136(w_003_136, w_000_1138, w_000_146);
  not1 I003_137(w_003_137, w_001_843);
  and2 I003_138(w_003_138, w_000_1590, w_001_160);
  or2  I003_139(w_003_139, w_002_039, w_002_303);
  not1 I003_140(w_003_140, w_002_547);
  not1 I003_141(w_003_141, w_001_1625);
  or2  I003_142(w_003_142, w_001_182, w_000_073);
  and2 I003_143(w_003_143, w_002_003, w_001_000);
  or2  I003_144(w_003_144, w_000_996, w_002_002);
  and2 I003_145(w_003_145, w_001_186, w_001_1144);
  nand2 I003_147(w_003_147, w_000_1644, w_002_063);
  and2 I003_148(w_003_148, w_001_138, w_000_918);
  or2  I003_149(w_003_149, w_000_1471, w_001_240);
  or2  I003_150(w_003_150, w_001_1683, w_000_734);
  nand2 I003_151(w_003_151, w_000_028, w_002_416);
  and2 I003_152(w_003_152, w_000_1174, w_001_1134);
  and2 I003_153(w_003_153, w_000_562, w_001_249);
  and2 I003_154(w_003_154, w_002_078, w_000_1183);
  not1 I003_155(w_003_155, w_001_1508);
  or2  I003_156(w_003_156, w_001_1438, w_000_904);
  or2  I003_157(w_003_157, w_001_1638, w_001_583);
  nand2 I003_158(w_003_158, w_002_163, w_002_145);
  not1 I003_159(w_003_159, w_001_183);
  not1 I003_160(w_003_160, w_002_436);
  or2  I003_161(w_003_161, w_001_1196, w_001_273);
  and2 I003_162(w_003_162, w_000_257, w_001_807);
  nand2 I003_163(w_003_163, w_002_004, w_001_125);
  nand2 I003_164(w_003_164, w_000_1645, w_001_1322);
  or2  I003_165(w_003_165, w_001_1026, w_000_893);
  and2 I003_166(w_003_166, w_001_767, w_001_903);
  nand2 I003_167(w_003_167, w_000_194, w_002_253);
  or2  I003_168(w_003_168, w_002_498, w_001_216);
  not1 I003_169(w_003_169, w_002_292);
  and2 I003_170(w_003_170, w_001_1647, w_000_1182);
  or2  I003_171(w_003_171, w_001_857, w_001_1361);
  nand2 I003_172(w_003_172, w_002_255, w_002_508);
  not1 I003_173(w_003_173, w_000_1411);
  or2  I003_174(w_003_174, w_001_1605, w_000_275);
  not1 I003_175(w_003_175, w_000_773);
  or2  I003_176(w_003_176, w_000_431, w_002_131);
  nand2 I003_177(w_003_177, w_002_373, w_002_352);
  and2 I003_178(w_003_178, w_000_1209, w_001_288);
  and2 I003_179(w_003_179, w_001_895, w_002_018);
  or2  I003_180(w_003_180, w_000_618, w_001_652);
  nand2 I003_181(w_003_181, w_002_333, w_002_501);
  or2  I003_182(w_003_182, w_002_340, w_000_1353);
  and2 I003_183(w_003_183, w_002_523, w_002_539);
  and2 I003_184(w_003_184, w_001_1465, w_001_154);
  or2  I003_185(w_003_185, w_000_852, w_001_761);
  nand2 I003_186(w_003_186, w_001_338, w_002_467);
  not1 I003_187(w_003_187, w_001_049);
  not1 I003_188(w_003_188, w_001_550);
  nand2 I003_189(w_003_189, w_000_891, w_001_1683);
  nand2 I003_190(w_003_190, w_001_206, w_002_276);
  not1 I003_191(w_003_191, w_000_688);
  and2 I003_192(w_003_192, w_001_793, w_000_992);
  not1 I003_193(w_003_193, w_000_1051);
  nand2 I003_194(w_003_194, w_002_432, w_001_154);
  or2  I003_195(w_003_195, w_001_072, w_001_1187);
  or2  I003_196(w_003_196, w_000_430, w_001_062);
  or2  I003_197(w_003_197, w_000_310, w_002_094);
  or2  I003_198(w_003_198, w_000_782, w_000_1340);
  and2 I003_199(w_003_199, w_000_333, w_002_346);
  and2 I003_200(w_003_200, w_000_388, w_001_428);
  and2 I003_201(w_003_201, w_002_471, w_002_407);
  and2 I003_202(w_003_202, w_001_1070, w_002_487);
  not1 I003_203(w_003_203, w_000_547);
  or2  I003_204(w_003_204, w_002_400, w_001_1486);
  and2 I003_205(w_003_205, w_001_827, w_002_218);
  and2 I003_206(w_003_206, w_002_104, w_001_282);
  and2 I003_207(w_003_207, w_002_158, w_001_1031);
  or2  I003_208(w_003_208, w_000_033, w_000_205);
  nand2 I003_209(w_003_209, w_000_1646, w_001_526);
  and2 I003_210(w_003_210, w_002_218, w_001_049);
  nand2 I003_211(w_003_211, w_001_1600, w_002_419);
  not1 I003_212(w_003_212, w_001_048);
  not1 I003_213(w_003_213, w_002_062);
  nand2 I003_214(w_003_214, w_000_814, w_002_095);
  and2 I003_215(w_003_215, w_000_480, w_000_1647);
  and2 I003_216(w_003_216, w_001_014, w_001_443);
  or2  I003_217(w_003_217, w_000_1256, w_001_096);
  nand2 I003_218(w_003_218, w_000_1386, w_002_122);
  and2 I003_219(w_003_219, w_000_212, w_002_021);
  not1 I003_220(w_003_220, w_001_1437);
  and2 I003_221(w_003_221, w_001_195, w_002_411);
  or2  I003_222(w_003_222, w_000_586, w_002_099);
  nand2 I003_223(w_003_223, w_000_542, w_001_1308);
  not1 I003_224(w_003_224, w_002_258);
  or2  I003_225(w_003_225, w_000_1184, w_000_728);
  and2 I003_226(w_003_226, w_000_940, w_000_1247);
  not1 I003_227(w_003_227, w_002_442);
  not1 I003_228(w_003_228, w_000_921);
  nand2 I003_229(w_003_229, w_000_1639, w_000_367);
  and2 I003_230(w_003_230, w_002_416, w_002_012);
  not1 I003_231(w_003_231, w_001_757);
  or2  I003_232(w_003_232, w_000_1166, w_002_265);
  or2  I003_233(w_003_233, w_000_1648, w_001_855);
  nand2 I003_234(w_003_234, w_000_773, w_002_228);
  and2 I003_235(w_003_235, w_001_053, w_001_953);
  not1 I003_236(w_003_236, w_001_1672);
  nand2 I003_237(w_003_237, w_000_1034, w_000_550);
  and2 I003_238(w_003_238, w_002_471, w_001_498);
  not1 I003_239(w_003_239, w_000_1649);
  nand2 I003_240(w_003_240, w_001_014, w_001_064);
  or2  I003_241(w_003_241, w_002_244, w_002_339);
  not1 I003_242(w_003_242, w_000_1028);
  or2  I003_243(w_003_243, w_001_763, w_000_843);
  not1 I003_244(w_003_244, w_001_188);
  or2  I003_245(w_003_245, w_000_1402, w_002_567);
  and2 I003_246(w_003_246, w_000_1650, w_000_177);
  and2 I003_247(w_003_247, w_002_191, w_001_075);
  and2 I003_248(w_003_248, w_001_1265, w_001_1605);
  nand2 I003_249(w_003_249, w_000_986, w_002_217);
  or2  I003_250(w_003_250, w_002_224, w_002_592);
  not1 I003_251(w_003_251, w_002_094);
  or2  I003_252(w_003_252, w_002_419, w_002_579);
  not1 I003_253(w_003_253, w_002_162);
  not1 I003_254(w_003_254, w_002_135);
  nand2 I003_255(w_003_255, w_002_271, w_001_115);
  and2 I003_256(w_003_256, w_002_351, w_000_819);
  nand2 I003_257(w_003_257, w_002_084, w_000_479);
  nand2 I003_258(w_003_258, w_001_122, w_001_243);
  nand2 I003_259(w_003_259, w_001_946, w_002_081);
  and2 I003_260(w_003_260, w_000_972, w_002_422);
  nand2 I003_261(w_003_261, w_000_460, w_002_130);
  and2 I003_262(w_003_262, w_002_181, w_002_141);
  nand2 I003_263(w_003_263, w_002_396, w_002_105);
  nand2 I003_264(w_003_264, w_002_187, w_001_882);
  and2 I003_265(w_003_265, w_002_008, w_001_307);
  not1 I003_266(w_003_266, w_000_1185);
  not1 I003_267(w_003_267, w_001_1147);
  or2  I003_268(w_003_268, w_001_270, w_001_910);
  and2 I003_269(w_003_269, w_001_1225, w_000_196);
  and2 I003_270(w_003_270, w_000_592, w_002_077);
  and2 I003_271(w_003_271, w_001_1452, w_000_1651);
  and2 I003_272(w_003_272, w_001_124, w_000_035);
  not1 I003_273(w_003_273, w_002_032);
  and2 I003_274(w_003_274, w_000_719, w_000_1652);
  nand2 I003_275(w_003_275, w_002_089, w_001_533);
  and2 I003_276(w_003_276, w_002_136, w_000_300);
  not1 I003_277(w_003_277, w_002_377);
  not1 I003_278(w_003_278, w_001_1369);
  and2 I003_279(w_003_279, w_001_1293, w_002_109);
  or2  I003_280(w_003_280, w_000_591, w_001_309);
  nand2 I003_281(w_003_281, w_001_1380, w_002_332);
  and2 I003_282(w_003_282, w_001_1609, w_002_076);
  or2  I003_283(w_003_283, w_002_212, w_001_366);
  or2  I003_284(w_003_284, w_001_283, w_002_587);
  and2 I003_285(w_003_285, w_000_949, w_001_881);
  not1 I003_286(w_003_286, w_000_1618);
  not1 I003_287(w_003_287, w_001_279);
  or2  I003_288(w_003_288, w_000_1653, w_002_173);
  and2 I003_289(w_003_289, w_000_1654, w_000_1222);
  and2 I003_290(w_003_290, w_002_380, w_002_483);
  or2  I003_291(w_003_291, w_002_172, w_001_1205);
  not1 I003_292(w_003_292, w_002_506);
  and2 I003_293(w_003_293, w_000_1105, w_002_002);
  nand2 I003_294(w_003_294, w_001_064, w_001_400);
  and2 I003_295(w_003_295, w_001_574, w_000_1400);
  and2 I003_296(w_003_296, w_000_974, w_001_275);
  nand2 I003_297(w_003_297, w_002_448, w_002_153);
  nand2 I003_298(w_003_298, w_001_898, w_000_170);
  or2  I003_299(w_003_299, w_002_202, w_002_276);
  and2 I003_300(w_003_300, w_001_617, w_002_075);
  or2  I003_301(w_003_301, w_001_112, w_002_056);
  or2  I003_302(w_003_302, w_000_256, w_001_026);
  or2  I003_303(w_003_303, w_002_439, w_001_1515);
  and2 I003_304(w_003_304, w_002_158, w_002_090);
  not1 I003_305(w_003_305, w_001_035);
  not1 I003_306(w_003_306, w_001_1499);
  nand2 I003_307(w_003_307, w_002_116, w_000_664);
  not1 I003_308(w_003_308, w_000_777);
  or2  I003_309(w_003_309, w_002_290, w_002_136);
  or2  I003_310(w_003_310, w_000_357, w_001_481);
  nand2 I003_311(w_003_311, w_001_112, w_000_427);
  or2  I003_312(w_003_312, w_001_1350, w_001_295);
  and2 I003_313(w_003_313, w_002_054, w_002_126);
  or2  I003_314(w_003_314, w_001_790, w_000_1375);
  nand2 I003_315(w_003_315, w_001_1255, w_001_006);
  and2 I003_316(w_003_316, w_000_508, w_002_311);
  or2  I003_317(w_003_317, w_002_580, w_002_262);
  or2  I003_318(w_003_318, w_002_211, w_002_567);
  not1 I003_319(w_003_319, w_001_1644);
  nand2 I004_000(w_004_000, w_002_448, w_002_077);
  nand2 I004_001(w_004_001, w_001_1184, w_003_209);
  not1 I004_002(w_004_002, w_001_881);
  or2  I004_003(w_004_003, w_001_982, w_000_1207);
  nand2 I004_004(w_004_004, w_002_216, w_003_095);
  nand2 I004_005(w_004_005, w_000_071, w_000_675);
  not1 I004_007(w_004_007, w_001_412);
  or2  I004_008(w_004_008, w_002_167, w_000_927);
  nand2 I004_009(w_004_009, w_002_026, w_000_347);
  or2  I004_011(w_004_011, w_001_593, w_000_1655);
  and2 I004_012(w_004_012, w_000_892, w_003_161);
  not1 I004_013(w_004_013, w_002_269);
  and2 I004_014(w_004_014, w_003_041, w_001_1045);
  not1 I004_015(w_004_015, w_002_191);
  or2  I004_016(w_004_016, w_000_1656, w_001_619);
  and2 I004_017(w_004_017, w_001_174, w_002_515);
  or2  I004_019(w_004_019, w_003_133, w_001_083);
  nand2 I004_021(w_004_021, w_002_183, w_002_332);
  and2 I004_022(w_004_022, w_003_284, w_002_059);
  not1 I004_024(w_004_024, w_000_480);
  nand2 I004_025(w_004_025, w_003_073, w_000_1387);
  not1 I004_027(w_004_027, w_003_254);
  or2  I004_028(w_004_028, w_001_028, w_003_245);
  not1 I004_029(w_004_029, w_003_129);
  and2 I004_030(w_004_030, w_000_025, w_003_294);
  not1 I004_031(w_004_031, w_000_996);
  nand2 I004_032(w_004_032, w_000_1067, w_002_072);
  or2  I004_035(w_004_035, w_001_022, w_000_1630);
  or2  I004_036(w_004_036, w_003_112, w_001_049);
  not1 I004_039(w_004_039, w_001_343);
  nand2 I004_041(w_004_041, w_000_312, w_001_221);
  nand2 I004_042(w_004_042, w_002_388, w_000_004);
  or2  I004_043(w_004_043, w_003_285, w_000_1487);
  nand2 I004_044(w_004_044, w_000_1658, w_003_170);
  nand2 I004_045(w_004_045, w_000_1152, w_002_295);
  not1 I004_046(w_004_046, w_003_304);
  and2 I004_047(w_004_047, w_001_1540, w_000_1297);
  and2 I004_048(w_004_048, w_001_1561, w_003_111);
  or2  I004_049(w_004_049, w_000_1396, w_002_079);
  or2  I004_050(w_004_050, w_003_114, w_000_1411);
  not1 I004_051(w_004_051, w_000_1659);
  or2  I004_054(w_004_054, w_000_749, w_001_254);
  and2 I004_056(w_004_056, w_000_1041, w_002_107);
  nand2 I004_057(w_004_057, w_001_1213, w_003_144);
  nand2 I004_058(w_004_058, w_003_045, w_001_319);
  nand2 I004_059(w_004_059, w_000_128, w_003_271);
  or2  I004_060(w_004_060, w_003_043, w_002_016);
  and2 I004_061(w_004_061, w_003_270, w_003_060);
  nand2 I004_062(w_004_062, w_003_180, w_001_517);
  and2 I004_063(w_004_063, w_000_1660, w_001_1583);
  nand2 I004_064(w_004_064, w_001_631, w_001_358);
  nand2 I004_066(w_004_066, w_003_233, w_000_810);
  and2 I004_068(w_004_068, w_000_850, w_000_1661);
  nand2 I004_070(w_004_070, w_000_1662, w_003_313);
  nand2 I004_071(w_004_071, w_000_1023, w_002_148);
  and2 I004_074(w_004_074, w_001_131, w_000_1663);
  or2  I004_075(w_004_075, w_000_160, w_000_1505);
  and2 I004_076(w_004_076, w_003_018, w_000_1512);
  nand2 I004_077(w_004_077, w_003_177, w_002_205);
  or2  I004_078(w_004_078, w_000_1323, w_003_285);
  not1 I004_079(w_004_079, w_002_027);
  nand2 I004_080(w_004_080, w_002_099, w_003_299);
  not1 I004_081(w_004_081, w_000_636);
  and2 I004_082(w_004_082, w_000_796, w_000_854);
  nand2 I004_084(w_004_084, w_000_1161, w_002_039);
  not1 I004_085(w_004_085, w_002_174);
  or2  I004_086(w_004_086, w_000_012, w_000_1623);
  nand2 I004_087(w_004_087, w_002_074, w_003_294);
  or2  I004_088(w_004_088, w_003_210, w_001_063);
  or2  I004_091(w_004_091, w_001_1511, w_003_008);
  not1 I004_093(w_004_093, w_003_145);
  and2 I004_095(w_004_095, w_003_126, w_001_855);
  or2  I004_096(w_004_096, w_003_124, w_001_1436);
  or2  I004_100(w_004_100, w_003_051, w_000_364);
  and2 I004_101(w_004_101, w_002_536, w_001_1589);
  and2 I004_102(w_004_102, w_000_995, w_002_321);
  not1 I004_104(w_004_104, w_003_307);
  nand2 I004_107(w_004_107, w_002_026, w_003_037);
  or2  I004_108(w_004_108, w_003_222, w_003_215);
  nand2 I004_109(w_004_109, w_000_1664, w_003_232);
  nand2 I004_111(w_004_111, w_003_294, w_000_845);
  or2  I004_112(w_004_112, w_000_1532, w_000_1665);
  or2  I004_114(w_004_114, w_000_536, w_000_1533);
  or2  I004_115(w_004_115, w_000_107, w_000_179);
  not1 I004_116(w_004_116, w_000_511);
  not1 I004_117(w_004_117, w_000_1137);
  or2  I004_118(w_004_118, w_001_086, w_000_391);
  and2 I004_120(w_004_120, w_001_155, w_002_349);
  or2  I004_121(w_004_121, w_002_049, w_001_1135);
  not1 I004_122(w_004_122, w_001_1243);
  not1 I004_123(w_004_123, w_001_1193);
  and2 I004_126(w_004_126, w_003_007, w_002_275);
  nand2 I004_130(w_004_130, w_002_322, w_000_1667);
  or2  I004_132(w_004_132, w_002_326, w_001_593);
  or2  I004_134(w_004_134, w_002_074, w_003_229);
  not1 I004_135(w_004_135, w_002_069);
  not1 I004_136(w_004_136, w_002_166);
  or2  I004_137(w_004_137, w_000_1445, w_000_1124);
  and2 I004_139(w_004_139, w_000_1411, w_001_005);
  nand2 I004_141(w_004_141, w_000_1090, w_002_235);
  and2 I004_142(w_004_142, w_000_086, w_002_538);
  or2  I004_143(w_004_143, w_003_138, w_002_281);
  not1 I004_144(w_004_144, w_000_167);
  not1 I004_146(w_004_146, w_002_170);
  not1 I004_147(w_004_147, w_000_830);
  or2  I004_148(w_004_148, w_002_161, w_001_1056);
  or2  I004_151(w_004_151, w_003_029, w_001_1197);
  or2  I004_152(w_004_152, w_000_801, w_003_143);
  not1 I004_153(w_004_153, w_001_1206);
  nand2 I004_156(w_004_156, w_002_194, w_002_259);
  and2 I004_157(w_004_157, w_003_058, w_001_138);
  or2  I004_159(w_004_159, w_003_206, w_003_128);
  and2 I004_160(w_004_160, w_003_258, w_001_815);
  nand2 I004_162(w_004_162, w_001_073, w_001_298);
  not1 I004_166(w_004_166, w_001_1551);
  nand2 I004_167(w_004_167, w_000_161, w_000_1667);
  not1 I004_170(w_004_170, w_001_1062);
  nand2 I004_171(w_004_171, w_000_704, w_003_037);
  or2  I004_172(w_004_172, w_003_269, w_000_850);
  nand2 I004_173(w_004_173, w_001_754, w_002_122);
  not1 I004_175(w_004_175, w_003_061);
  or2  I004_176(w_004_176, w_002_526, w_002_082);
  nand2 I004_177(w_004_177, w_003_090, w_002_229);
  and2 I004_179(w_004_179, w_001_1081, w_000_384);
  or2  I004_181(w_004_181, w_002_213, w_000_587);
  nand2 I004_182(w_004_182, w_003_008, w_000_693);
  and2 I004_183(w_004_183, w_002_534, w_003_066);
  not1 I004_185(w_004_185, w_003_129);
  nand2 I004_186(w_004_186, w_003_113, w_000_1120);
  nand2 I004_187(w_004_187, w_000_1192, w_001_214);
  or2  I004_188(w_004_188, w_001_801, w_000_668);
  and2 I004_190(w_004_190, w_001_1485, w_000_271);
  not1 I004_191(w_004_191, w_003_179);
  and2 I004_192(w_004_192, w_002_548, w_000_221);
  or2  I004_194(w_004_194, w_000_886, w_002_484);
  nand2 I004_195(w_004_195, w_003_279, w_003_036);
  and2 I004_196(w_004_196, w_003_150, w_002_038);
  not1 I004_197(w_004_197, w_003_243);
  not1 I004_199(w_004_199, w_001_1382);
  and2 I004_200(w_004_200, w_001_1042, w_002_307);
  nand2 I004_201(w_004_201, w_000_925, w_003_286);
  nand2 I004_202(w_004_202, w_002_303, w_003_105);
  not1 I004_206(w_004_206, w_000_1391);
  and2 I004_207(w_004_207, w_002_511, w_003_086);
  or2  I004_209(w_004_209, w_002_480, w_001_007);
  and2 I004_210(w_004_210, w_000_402, w_000_714);
  or2  I004_211(w_004_211, w_003_104, w_003_276);
  not1 I004_213(w_004_213, w_002_420);
  or2  I004_214(w_004_214, w_001_106, w_001_528);
  not1 I004_215(w_004_215, w_000_1177);
  nand2 I004_216(w_004_216, w_003_252, w_000_720);
  and2 I004_217(w_004_217, w_001_1123, w_001_635);
  and2 I004_218(w_004_218, w_000_1091, w_003_177);
  or2  I004_220(w_004_220, w_002_109, w_002_424);
  not1 I004_222(w_004_222, w_001_423);
  not1 I004_223(w_004_223, w_002_307);
  nand2 I004_225(w_004_225, w_002_497, w_000_1518);
  not1 I004_226(w_004_226, w_001_673);
  and2 I004_227(w_004_227, w_000_1233, w_001_186);
  and2 I004_229(w_004_229, w_000_1151, w_000_1442);
  and2 I004_232(w_004_232, w_002_366, w_002_119);
  nand2 I004_233(w_004_233, w_003_116, w_001_416);
  not1 I004_234(w_004_234, w_001_954);
  not1 I004_235(w_004_235, w_001_1599);
  not1 I004_236(w_004_236, w_001_751);
  not1 I004_241(w_004_241, w_000_1673);
  and2 I004_243(w_004_243, w_000_1378, w_000_591);
  nand2 I004_245(w_004_245, w_000_1674, w_003_168);
  nand2 I004_246(w_004_246, w_000_1086, w_000_1675);
  not1 I004_248(w_004_248, w_000_1171);
  not1 I004_249(w_004_249, w_000_293);
  and2 I004_250(w_004_250, w_002_128, w_001_576);
  not1 I004_251(w_004_251, w_000_1676);
  or2  I004_252(w_004_252, w_001_054, w_000_028);
  nand2 I004_254(w_004_254, w_003_001, w_000_1501);
  not1 I004_257(w_004_257, w_001_033);
  and2 I004_258(w_004_258, w_003_152, w_001_1269);
  and2 I004_259(w_004_259, w_001_1502, w_001_1102);
  not1 I004_260(w_004_260, w_002_255);
  and2 I004_261(w_004_261, w_001_888, w_001_765);
  nand2 I004_262(w_004_262, w_003_297, w_000_1417);
  not1 I004_264(w_004_264, w_003_205);
  and2 I004_265(w_004_265, w_002_116, w_003_178);
  nand2 I004_266(w_004_266, w_001_566, w_000_1447);
  and2 I004_269(w_004_269, w_000_792, w_003_185);
  and2 I004_275(w_004_275, w_000_783, w_002_187);
  not1 I004_276(w_004_276, w_003_043);
  not1 I004_277(w_004_277, w_000_1554);
  and2 I004_278(w_004_278, w_001_482, w_000_1218);
  or2  I004_279(w_004_279, w_002_103, w_001_107);
  or2  I004_280(w_004_280, w_000_1307, w_002_349);
  not1 I004_283(w_004_283, w_000_752);
  and2 I004_286(w_004_286, w_001_268, w_001_1202);
  nand2 I004_288(w_004_288, w_000_1266, w_000_594);
  and2 I004_292(w_004_292, w_002_031, w_000_395);
  nand2 I004_293(w_004_293, w_001_260, w_000_1678);
  nand2 I004_296(w_004_296, w_003_081, w_000_281);
  nand2 I004_298(w_004_298, w_002_053, w_002_046);
  not1 I004_300(w_004_300, w_002_103);
  and2 I004_301(w_004_301, w_001_969, w_001_030);
  or2  I004_303(w_004_303, w_003_181, w_002_299);
  or2  I004_305(w_004_305, w_002_469, w_003_304);
  not1 I004_307(w_004_307, w_000_1403);
  nand2 I004_310(w_004_310, w_003_262, w_002_288);
  nand2 I004_312(w_004_312, w_002_110, w_002_436);
  not1 I004_313(w_004_313, w_002_467);
  and2 I004_314(w_004_314, w_003_051, w_000_618);
  not1 I004_315(w_004_315, w_001_005);
  or2  I004_316(w_004_316, w_002_231, w_001_273);
  or2  I004_318(w_004_318, w_003_266, w_001_438);
  or2  I004_319(w_004_319, w_003_229, w_003_153);
  not1 I004_321(w_004_321, w_003_199);
  and2 I004_322(w_004_322, w_000_1680, w_001_794);
  or2  I004_323(w_004_323, w_002_515, w_000_1034);
  not1 I004_324(w_004_324, w_002_550);
  nand2 I004_325(w_004_325, w_001_266, w_000_1119);
  or2  I004_326(w_004_326, w_003_068, w_000_200);
  and2 I004_328(w_004_328, w_001_865, w_000_197);
  or2  I004_331(w_004_331, w_001_194, w_002_321);
  nand2 I004_334(w_004_334, w_003_159, w_000_676);
  or2  I004_337(w_004_337, w_003_172, w_003_077);
  not1 I004_340(w_004_340, w_002_119);
  or2  I004_342(w_004_342, w_001_1320, w_002_119);
  not1 I004_343(w_004_343, w_003_034);
  not1 I004_345(w_004_345, w_000_1454);
  not1 I004_346(w_004_346, w_000_1682);
  and2 I004_352(w_004_352, w_002_215, w_000_980);
  nand2 I004_353(w_004_353, w_001_1289, w_000_1290);
  or2  I004_355(w_004_355, w_002_591, w_002_054);
  and2 I004_356(w_004_356, w_001_988, w_000_424);
  or2  I004_359(w_004_359, w_000_1683, w_000_1684);
  and2 I004_361(w_004_361, w_000_744, w_001_558);
  and2 I004_362(w_004_362, w_001_407, w_000_565);
  and2 I004_364(w_004_364, w_000_509, w_000_171);
  and2 I004_366(w_004_366, w_002_120, w_003_093);
  and2 I004_368(w_004_368, w_000_1522, w_000_120);
  and2 I004_369(w_004_369, w_003_006, w_003_200);
  nand2 I004_371(w_004_371, w_000_1128, w_000_1509);
  nand2 I004_372(w_004_372, w_000_871, w_000_494);
  or2  I004_373(w_004_373, w_003_268, w_000_1559);
  not1 I004_374(w_004_374, w_000_300);
  not1 I004_375(w_004_375, w_000_174);
  not1 I004_377(w_004_377, w_003_093);
  nand2 I004_379(w_004_379, w_001_151, w_003_025);
  not1 I004_380(w_004_380, w_002_019);
  and2 I004_382(w_004_382, w_003_261, w_002_259);
  or2  I004_383(w_004_383, w_000_803, w_003_259);
  nand2 I004_384(w_004_384, w_002_303, w_002_035);
  nand2 I004_385(w_004_385, w_000_068, w_002_465);
  and2 I004_388(w_004_388, w_003_175, w_001_079);
  not1 I004_391(w_004_391, w_003_043);
  or2  I004_394(w_004_394, w_003_264, w_001_1079);
  and2 I004_395(w_004_395, w_000_1254, w_002_266);
  and2 I004_396(w_004_396, w_000_456, w_001_698);
  not1 I004_398(w_004_398, w_000_039);
  not1 I004_399(w_004_399, w_000_663);
  nand2 I004_400(w_004_400, w_002_049, w_001_571);
  and2 I004_402(w_004_402, w_000_461, w_002_226);
  nand2 I004_404(w_004_404, w_003_115, w_002_396);
  nand2 I004_406(w_004_406, w_003_189, w_000_184);
  or2  I004_407(w_004_407, w_003_312, w_000_831);
  not1 I004_409(w_004_409, w_001_1209);
  and2 I004_415(w_004_415, w_001_764, w_000_111);
  nand2 I004_416(w_004_416, w_001_1320, w_000_804);
  not1 I004_417(w_004_417, w_000_443);
  and2 I004_418(w_004_418, w_003_189, w_003_053);
  not1 I004_420(w_004_420, w_002_472);
  not1 I004_422(w_004_422, w_003_010);
  nand2 I004_425(w_004_425, w_000_1434, w_003_133);
  nand2 I004_428(w_004_428, w_002_404, w_002_044);
  not1 I004_429(w_004_429, w_001_458);
  or2  I004_430(w_004_430, w_000_1577, w_002_396);
  or2  I004_433(w_004_433, w_003_170, w_003_021);
  nand2 I004_435(w_004_435, w_001_1179, w_001_1379);
  or2  I004_436(w_004_436, w_003_023, w_002_135);
  nand2 I004_437(w_004_437, w_002_022, w_001_629);
  not1 I004_443(w_004_443, w_000_1567);
  not1 I004_444(w_004_444, w_002_197);
  or2  I004_445(w_004_445, w_003_201, w_001_096);
  and2 I004_446(w_004_446, w_002_038, w_001_954);
  nand2 I004_447(w_004_447, w_003_272, w_001_1332);
  and2 I004_448(w_004_448, w_002_552, w_002_226);
  and2 I004_449(w_004_449, w_002_426, w_001_1207);
  and2 I004_451(w_004_451, w_000_1071, w_001_761);
  or2  I004_452(w_004_452, w_001_543, w_001_442);
  or2  I004_453(w_004_453, w_000_133, w_002_143);
  or2  I004_454(w_004_454, w_002_309, w_000_1220);
  or2  I004_458(w_004_458, w_002_015, w_002_507);
  not1 I004_459(w_004_459, w_003_169);
  and2 I004_460(w_004_460, w_003_303, w_002_182);
  not1 I004_462(w_004_462, w_000_1688);
  or2  I004_469(w_004_469, w_000_1256, w_002_075);
  or2  I004_472(w_004_472, w_002_512, w_002_247);
  not1 I004_476(w_004_476, w_001_421);
  not1 I004_477(w_004_477, w_000_250);
  or2  I004_478(w_004_478, w_000_180, w_002_005);
  or2  I004_481(w_004_481, w_003_183, w_001_209);
  and2 I004_482(w_004_482, w_001_357, w_002_258);
  and2 I004_483(w_004_483, w_000_752, w_001_1269);
  or2  I004_486(w_004_486, w_002_157, w_000_349);
  not1 I004_487(w_004_487, w_001_1084);
  or2  I004_488(w_004_488, w_003_056, w_002_204);
  nand2 I004_490(w_004_490, w_002_131, w_002_243);
  or2  I004_491(w_004_491, w_002_517, w_001_316);
  and2 I004_492(w_004_492, w_003_059, w_001_865);
  and2 I004_493(w_004_493, w_001_1567, w_003_051);
  nand2 I004_494(w_004_494, w_000_1646, w_003_314);
  and2 I004_496(w_004_496, w_001_1402, w_003_307);
  and2 I004_498(w_004_498, w_002_428, w_000_665);
  nand2 I004_501(w_004_501, w_000_1690, w_001_1177);
  not1 I004_503(w_004_503, w_003_291);
  or2  I004_504(w_004_504, w_000_034, w_001_482);
  not1 I004_506(w_004_506, w_002_435);
  not1 I004_507(w_004_507, w_000_479);
  or2  I004_510(w_004_510, w_000_134, w_002_118);
  and2 I004_512(w_004_512, w_003_030, w_001_198);
  and2 I004_513(w_004_513, w_003_299, w_002_205);
  not1 I004_514(w_004_514, w_003_061);
  not1 I004_515(w_004_515, w_000_1399);
  nand2 I004_516(w_004_516, w_002_390, w_000_521);
  nand2 I004_517(w_004_517, w_000_1007, w_001_064);
  and2 I004_518(w_004_518, w_003_061, w_001_1587);
  not1 I004_520(w_004_520, w_001_570);
  nand2 I004_524(w_004_524, w_000_045, w_000_1163);
  not1 I004_527(w_004_527, w_002_005);
  nand2 I004_528(w_004_528, w_002_110, w_002_368);
  or2  I004_529(w_004_529, w_000_144, w_001_270);
  and2 I004_530(w_004_530, w_003_241, w_000_527);
  nand2 I004_534(w_004_534, w_001_1373, w_003_227);
  nand2 I004_535(w_004_535, w_001_195, w_000_1690);
  nand2 I004_537(w_004_537, w_000_737, w_002_258);
  nand2 I004_538(w_004_538, w_000_330, w_000_579);
  not1 I004_540(w_004_540, w_000_1693);
  not1 I004_543(w_004_543, w_000_998);
  not1 I004_544(w_004_544, w_002_378);
  nand2 I004_545(w_004_545, w_003_076, w_003_074);
  or2  I004_546(w_004_546, w_001_1246, w_000_1247);
  not1 I004_547(w_004_547, w_000_776);
  and2 I004_548(w_004_548, w_003_308, w_001_577);
  nand2 I004_550(w_004_550, w_001_209, w_003_271);
  or2  I004_551(w_004_551, w_002_210, w_003_280);
  or2  I004_552(w_004_552, w_002_308, w_000_293);
  or2  I004_553(w_004_553, w_002_351, w_001_549);
  not1 I004_554(w_004_554, w_002_137);
  not1 I004_555(w_004_555, w_001_1266);
  nand2 I004_558(w_004_558, w_000_913, w_002_018);
  nand2 I004_560(w_004_560, w_002_132, w_001_1661);
  and2 I004_561(w_004_561, w_002_021, w_002_311);
  or2  I004_562(w_004_562, w_003_297, w_000_1433);
  or2  I004_563(w_004_563, w_003_233, w_000_1291);
  and2 I004_565(w_004_565, w_000_1684, w_002_277);
  or2  I004_566(w_004_566, w_001_1587, w_003_066);
  not1 I004_571(w_004_571, w_003_220);
  nand2 I004_575(w_004_575, w_003_006, w_001_916);
  nand2 I004_576(w_004_576, w_003_317, w_002_071);
  and2 I004_579(w_004_579, w_001_063, w_003_308);
  or2  I004_581(w_004_581, w_000_1387, w_000_831);
  or2  I004_583(w_004_583, w_003_161, w_001_119);
  nand2 I004_584(w_004_584, w_000_354, w_003_134);
  and2 I004_585(w_004_585, w_003_249, w_001_120);
  or2  I004_587(w_004_587, w_002_003, w_002_342);
  or2  I004_588(w_004_588, w_002_338, w_002_185);
  or2  I004_590(w_004_590, w_000_1084, w_000_1484);
  not1 I004_591(w_004_591, w_003_290);
  nand2 I004_592(w_004_592, w_002_460, w_000_1474);
  not1 I004_593(w_004_593, w_000_926);
  or2  I004_595(w_004_595, w_003_031, w_003_310);
  or2  I004_596(w_004_596, w_003_038, w_003_122);
  nand2 I004_597(w_004_597, w_003_166, w_003_075);
  or2  I004_598(w_004_598, w_002_412, w_000_1485);
  not1 I004_599(w_004_599, w_000_1311);
  nand2 I004_602(w_004_602, w_001_1452, w_002_511);
  or2  I004_603(w_004_603, w_001_1049, w_001_423);
  and2 I004_604(w_004_604, w_000_910, w_003_004);
  nand2 I004_605(w_004_605, w_002_494, w_003_223);
  and2 I004_606(w_004_606, w_003_286, w_000_1187);
  and2 I004_607(w_004_607, w_000_615, w_002_274);
  not1 I004_609(w_004_609, w_002_589);
  and2 I004_610(w_004_610, w_003_201, w_000_951);
  nand2 I004_611(w_004_611, w_000_1627, w_002_216);
  not1 I004_615(w_004_615, w_000_271);
  nand2 I004_616(w_004_616, w_000_1666, w_001_625);
  not1 I004_617(w_004_617, w_000_826);
  not1 I004_618(w_004_618, w_003_289);
  and2 I004_620(w_004_620, w_000_320, w_001_156);
  nand2 I004_624(w_004_624, w_000_961, w_001_1074);
  or2  I004_625(w_004_625, w_003_221, w_000_197);
  nand2 I004_626(w_004_626, w_003_240, w_000_1564);
  not1 I004_628(w_004_628, w_001_091);
  nand2 I004_633(w_004_633, w_003_069, w_003_072);
  not1 I004_635(w_004_635, w_001_1127);
  and2 I004_636(w_004_636, w_001_1023, w_000_1694);
  nand2 I004_637(w_004_637, w_001_1070, w_001_074);
  and2 I004_638(w_004_638, w_003_016, w_003_224);
  nand2 I004_639(w_004_639, w_002_172, w_002_539);
  and2 I004_640(w_004_640, w_001_1125, w_001_1192);
  not1 I004_641(w_004_641, w_000_1695);
  or2  I004_642(w_004_642, w_002_350, w_001_307);
  or2  I004_644(w_004_644, w_000_532, w_002_139);
  and2 I004_645(w_004_645, w_001_832, w_003_079);
  not1 I004_646(w_004_646, w_001_525);
  and2 I004_652(w_004_652, w_000_746, w_001_168);
  or2  I004_653(w_004_653, w_001_1306, w_002_266);
  or2  I004_655(w_004_655, w_001_132, w_003_056);
  nand2 I004_656(w_004_656, w_002_141, w_001_1130);
  not1 I004_657(w_004_657, w_001_524);
  and2 I004_659(w_004_659, w_001_1550, w_001_1578);
  or2  I004_661(w_004_661, w_002_182, w_002_004);
  or2  I004_663(w_004_663, w_001_235, w_003_114);
  nand2 I004_664(w_004_664, w_003_192, w_002_243);
  not1 I004_665(w_004_665, w_002_081);
  or2  I004_670(w_004_670, w_002_116, w_000_1277);
  and2 I004_671(w_004_671, w_002_467, w_003_085);
  not1 I004_672(w_004_672, w_003_281);
  and2 I004_677(w_004_677, w_001_854, w_002_213);
  nand2 I004_678(w_004_678, w_000_1341, w_001_1273);
  and2 I004_680(w_004_680, w_000_400, w_002_153);
  nand2 I004_683(w_004_683, w_003_017, w_002_261);
  or2  I004_687(w_004_687, w_000_700, w_000_1036);
  nand2 I004_694(w_004_694, w_000_366, w_002_224);
  and2 I004_695(w_004_695, w_003_143, w_002_171);
  or2  I004_697(w_004_697, w_000_162, w_003_291);
  and2 I004_700(w_004_700, w_001_031, w_003_294);
  or2  I004_701(w_004_701, w_001_140, w_001_054);
  not1 I004_703(w_004_703, w_001_650);
  nand2 I004_704(w_004_704, w_001_1164, w_003_056);
  nand2 I004_705(w_004_705, w_001_580, w_003_163);
  not1 I004_706(w_004_706, w_003_098);
  not1 I004_710(w_004_710, w_000_1457);
  not1 I004_711(w_004_711, w_002_286);
  and2 I004_713(w_004_713, w_000_622, w_000_039);
  or2  I004_714(w_004_714, w_002_094, w_003_073);
  nand2 I004_715(w_004_715, w_000_179, w_002_256);
  not1 I004_717(w_004_717, w_003_019);
  and2 I004_719(w_004_719, w_002_261, w_002_064);
  not1 I004_721(w_004_721, w_000_823);
  or2  I004_722(w_004_722, w_002_022, w_003_025);
  nand2 I004_723(w_004_723, w_003_030, w_002_093);
  and2 I004_724(w_004_724, w_000_1113, w_002_099);
  and2 I004_725(w_004_725, w_001_1053, w_000_1563);
  not1 I004_726(w_004_726, w_003_084);
  and2 I004_727(w_004_727, w_001_216, w_002_168);
  or2  I004_730(w_004_730, w_000_1703, w_003_289);
  or2  I004_731(w_004_731, w_003_075, w_003_038);
  nand2 I004_732(w_004_732, w_000_1012, w_000_1704);
  not1 I004_733(w_004_733, w_003_156);
  and2 I004_737(w_004_737, w_001_1399, w_003_027);
  and2 I004_738(w_004_738, w_002_342, w_003_313);
  or2  I004_739(w_004_739, w_000_317, w_001_875);
  not1 I004_743(w_004_743, w_003_236);
  not1 I004_744(w_004_744, w_000_948);
  and2 I004_746(w_004_746, w_000_843, w_000_725);
  not1 I004_749(w_004_749, w_000_1303);
  nand2 I004_750(w_004_750, w_001_1497, w_002_560);
  not1 I004_753(w_004_753, w_000_199);
  not1 I004_754(w_004_754, w_001_759);
  not1 I004_755(w_004_755, w_002_020);
  or2  I004_756(w_004_756, w_003_154, w_002_478);
  not1 I004_757(w_004_757, w_000_370);
  or2  I004_758(w_004_758, w_003_008, w_002_078);
  not1 I004_762(w_004_762, w_002_187);
  and2 I004_764(w_004_764, w_002_395, w_000_1465);
  or2  I004_765(w_004_765, w_000_145, w_003_002);
  nand2 I004_766(w_004_766, w_001_147, w_003_238);
  not1 I004_768(w_004_768, w_002_132);
  and2 I004_769(w_004_769, w_002_431, w_002_483);
  nand2 I004_770(w_004_770, w_001_1506, w_003_010);
  not1 I004_771(w_004_771, w_002_083);
  nand2 I004_772(w_004_772, w_003_006, w_003_272);
  nand2 I004_774(w_004_774, w_000_1706, w_001_056);
  nand2 I004_775(w_004_775, w_001_1240, w_002_019);
  and2 I004_777(w_004_777, w_000_853, w_003_086);
  and2 I004_778(w_004_778, w_001_044, w_003_244);
  and2 I004_780(w_004_780, w_003_079, w_003_235);
  not1 I004_782(w_004_782, w_003_267);
  nand2 I004_783(w_004_783, w_003_212, w_002_182);
  and2 I004_785(w_004_785, w_001_393, w_003_141);
  or2  I004_787(w_004_787, w_000_1063, w_003_261);
  and2 I004_788(w_004_788, w_000_1367, w_002_515);
  not1 I004_790(w_004_790, w_000_1096);
  nand2 I004_796(w_004_796, w_000_1707, w_002_452);
  not1 I004_797(w_004_797, w_001_1500);
  and2 I004_798(w_004_798, w_003_252, w_000_038);
  nand2 I004_799(w_004_799, w_001_1428, w_003_305);
  and2 I004_803(w_004_803, w_002_278, w_002_113);
  and2 I004_804(w_004_804, w_002_129, w_000_354);
  or2  I004_805(w_004_805, w_003_227, w_001_000);
  nand2 I004_807(w_004_807, w_003_301, w_001_521);
  and2 I004_809(w_004_809, w_000_1524, w_000_282);
  and2 I004_810(w_004_810, w_000_1709, w_003_284);
  not1 I004_813(w_004_813, w_001_1588);
  or2  I004_814(w_004_814, w_001_200, w_003_242);
  or2  I004_815(w_004_815, w_001_817, w_002_299);
  not1 I004_816(w_004_816, w_002_175);
  not1 I004_817(w_004_817, w_001_257);
  nand2 I004_818(w_004_818, w_001_1146, w_003_284);
  not1 I004_819(w_004_819, w_003_071);
  not1 I004_823(w_004_823, w_003_115);
  or2  I004_824(w_004_824, w_003_285, w_002_086);
  nand2 I004_826(w_004_826, w_003_287, w_003_168);
  or2  I004_827(w_004_827, w_003_271, w_001_110);
  nand2 I004_828(w_004_828, w_002_223, w_003_086);
  not1 I004_830(w_004_830, w_003_318);
  nand2 I004_831(w_004_831, w_001_1076, w_000_977);
  or2  I004_832(w_004_832, w_000_553, w_001_015);
  not1 I004_834(w_004_834, w_003_300);
  nand2 I004_836(w_004_836, w_000_1530, w_002_405);
  and2 I004_837(w_004_837, w_001_1637, w_000_075);
  or2  I004_838(w_004_838, w_000_1052, w_003_188);
  or2  I004_839(w_004_839, w_000_155, w_001_1436);
  not1 I004_840(w_004_840, w_002_575);
  and2 I004_841(w_004_841, w_001_177, w_001_527);
  nand2 I004_842(w_004_842, w_002_092, w_002_010);
  or2  I004_843(w_004_843, w_000_549, w_001_898);
  not1 I004_846(w_004_846, w_002_028);
  not1 I004_848(w_004_848, w_003_289);
  nand2 I004_850(w_004_850, w_000_421, w_003_033);
  not1 I004_852(w_004_852, w_002_421);
  or2  I004_853(w_004_853, w_003_101, w_003_136);
  and2 I004_854(w_004_854, w_002_212, w_002_034);
  not1 I004_856(w_004_856, w_003_075);
  or2  I004_860(w_004_860, w_002_360, w_002_132);
  or2  I004_862(w_004_862, w_002_076, w_003_173);
  or2  I004_866(w_004_866, w_001_649, w_003_235);
  and2 I004_868(w_004_868, w_003_076, w_000_1674);
  and2 I004_870(w_004_870, w_002_330, w_003_018);
  or2  I004_871(w_004_871, w_002_447, w_001_1634);
  not1 I004_872(w_004_872, w_002_037);
  nand2 I004_876(w_004_876, w_003_100, w_003_237);
  or2  I004_877(w_004_877, w_002_267, w_002_257);
  not1 I004_878(w_004_878, w_003_119);
  or2  I004_879(w_004_879, w_002_062, w_001_556);
  or2  I004_881(w_004_881, w_002_453, w_001_711);
  not1 I004_884(w_004_884, w_003_134);
  and2 I004_885(w_004_885, w_003_253, w_001_1441);
  nand2 I004_886(w_004_886, w_002_215, w_003_037);
  not1 I004_888(w_004_888, w_001_227);
  or2  I004_890(w_004_890, w_000_209, w_000_039);
  or2  I004_892(w_004_892, w_000_669, w_000_1562);
  or2  I004_894(w_004_894, w_002_593, w_001_223);
  not1 I004_895(w_004_895, w_000_307);
  nand2 I004_896(w_004_896, w_001_489, w_003_102);
  not1 I004_897(w_004_897, w_003_023);
  nand2 I004_898(w_004_898, w_002_183, w_001_755);
  nand2 I004_899(w_004_899, w_001_1425, w_003_191);
  and2 I004_900(w_004_900, w_001_661, w_001_151);
  not1 I004_901(w_004_901, w_000_1710);
  or2  I004_904(w_004_904, w_003_123, w_001_495);
  not1 I004_905(w_004_905, w_003_172);
  nand2 I004_907(w_004_907, w_000_604, w_000_1711);
  or2  I004_908(w_004_908, w_003_135, w_001_214);
  nand2 I004_909(w_004_909, w_002_059, w_002_390);
  not1 I004_910(w_004_910, w_003_167);
  or2  I004_912(w_004_912, w_000_478, w_001_687);
  or2  I004_914(w_004_914, w_002_005, w_001_1412);
  not1 I004_916(w_004_916, w_000_360);
  or2  I004_917(w_004_917, w_003_174, w_000_1426);
  not1 I004_918(w_004_918, w_003_069);
  not1 I004_920(w_004_920, w_000_1168);
  or2  I004_921(w_004_921, w_002_032, w_000_1283);
  and2 I004_922(w_004_922, w_003_108, w_000_100);
  or2  I004_925(w_004_925, w_000_580, w_000_986);
  nand2 I004_926(w_004_926, w_001_485, w_001_184);
  nand2 I004_929(w_004_929, w_001_1522, w_003_029);
  and2 I004_931(w_004_931, w_002_117, w_002_321);
  or2  I004_933(w_004_933, w_000_1194, w_002_053);
  or2  I004_934(w_004_934, w_003_305, w_002_032);
  and2 I004_935(w_004_935, w_000_1628, w_003_081);
  and2 I004_937(w_004_937, w_002_119, w_000_1712);
  not1 I004_938(w_004_938, w_002_393);
  or2  I004_941(w_004_941, w_001_191, w_000_1391);
  nand2 I004_942(w_004_942, w_000_1019, w_002_533);
  or2  I004_943(w_004_943, w_001_275, w_001_183);
  not1 I004_949(w_004_949, w_001_200);
  or2  I004_950(w_004_950, w_003_073, w_001_069);
  nand2 I004_952(w_004_952, w_000_084, w_002_427);
  or2  I004_953(w_004_953, w_002_119, w_001_123);
  or2  I004_955(w_004_955, w_001_121, w_003_243);
  nand2 I004_957(w_004_957, w_002_180, w_000_1079);
  and2 I004_958(w_004_958, w_003_047, w_000_1374);
  not1 I004_959(w_004_959, w_001_116);
  nand2 I004_960(w_004_960, w_002_239, w_003_142);
  and2 I004_962(w_004_962, w_003_260, w_002_367);
  not1 I004_963(w_004_963, w_000_1024);
  or2  I004_964(w_004_964, w_003_072, w_002_182);
  not1 I004_970(w_004_970, w_003_235);
  and2 I004_973(w_004_973, w_003_138, w_003_071);
  not1 I004_975(w_004_975, w_000_1427);
  or2  I004_977(w_004_977, w_000_923, w_001_244);
  nand2 I004_978(w_004_978, w_003_174, w_000_1716);
  nand2 I004_979(w_004_979, w_001_1134, w_000_152);
  and2 I004_980(w_004_980, w_003_143, w_001_409);
  not1 I004_981(w_004_981, w_000_1717);
  not1 I004_983(w_004_983, w_001_048);
  and2 I004_984(w_004_984, w_001_1324, w_001_556);
  nand2 I004_985(w_004_985, w_001_1050, w_003_316);
  not1 I004_987(w_004_987, w_000_1314);
  and2 I004_989(w_004_989, w_003_058, w_000_1554);
  not1 I004_990(w_004_990, w_000_137);
  nand2 I004_991(w_004_991, w_001_1149, w_000_1649);
  nand2 I004_993(w_004_993, w_003_120, w_003_085);
  and2 I004_994(w_004_994, w_001_1423, w_001_1684);
  and2 I004_996(w_004_996, w_002_117, w_000_320);
  nand2 I004_997(w_004_997, w_000_457, w_002_457);
  not1 I004_1001(w_004_1001, w_000_081);
  or2  I004_1004(w_004_1004, w_002_414, w_000_1219);
  or2  I004_1008(w_004_1008, w_002_105, w_002_344);
  not1 I004_1009(w_004_1009, w_000_816);
  not1 I004_1011(w_004_1011, w_001_779);
  or2  I004_1015(w_004_1015, w_000_667, w_001_1005);
  or2  I004_1016(w_004_1016, w_003_295, w_001_1065);
  nand2 I004_1017(w_004_1017, w_001_349, w_001_1482);
  and2 I004_1020(w_004_1020, w_003_070, w_002_111);
  and2 I004_1021(w_004_1021, w_003_200, w_002_525);
  nand2 I004_1023(w_004_1023, w_002_067, w_003_112);
  not1 I004_1025(w_004_1025, w_003_160);
  not1 I004_1027(w_004_1027, w_003_019);
  and2 I004_1028(w_004_1028, w_002_173, w_003_094);
  or2  I004_1029(w_004_1029, w_002_274, w_001_646);
  nand2 I004_1030(w_004_1030, w_003_090, w_001_057);
  or2  I004_1033(w_004_1033, w_001_034, w_001_1570);
  not1 I004_1035(w_004_1035, w_002_550);
  and2 I004_1037(w_004_1037, w_003_255, w_003_054);
  not1 I004_1038(w_004_1038, w_001_1059);
  or2  I004_1039(w_004_1039, w_002_303, w_001_395);
  and2 I004_1040(w_004_1040, w_003_256, w_002_135);
  and2 I004_1043(w_004_1043, w_001_001, w_001_1431);
  nand2 I004_1046(w_004_1046, w_003_318, w_003_059);
  nand2 I004_1047(w_004_1047, w_002_388, w_001_696);
  and2 I004_1049(w_004_1049, w_002_268, w_000_1439);
  or2  I004_1050(w_004_1050, w_002_277, w_002_268);
  or2  I004_1051(w_004_1051, w_003_273, w_002_102);
  not1 I004_1053(w_004_1053, w_001_1467);
  or2  I004_1054(w_004_1054, w_003_115, w_002_096);
  or2  I004_1056(w_004_1056, w_002_137, w_002_144);
  or2  I004_1061(w_004_1061, w_002_284, w_002_319);
  nand2 I004_1062(w_004_1062, w_003_077, w_000_209);
  or2  I004_1063(w_004_1063, w_000_662, w_000_1598);
  nand2 I004_1065(w_004_1065, w_001_406, w_000_552);
  and2 I004_1066(w_004_1066, w_001_1540, w_002_120);
  or2  I004_1069(w_004_1069, w_000_1722, w_002_233);
  or2  I004_1071(w_004_1071, w_000_1723, w_000_941);
  nand2 I004_1073(w_004_1073, w_002_197, w_001_732);
  and2 I004_1074(w_004_1074, w_000_980, w_000_102);
  nand2 I004_1076(w_004_1076, w_003_150, w_000_193);
  or2  I004_1077(w_004_1077, w_002_119, w_002_214);
  nand2 I004_1078(w_004_1078, w_002_344, w_002_174);
  and2 I004_1080(w_004_1080, w_003_078, w_000_1615);
  or2  I004_1082(w_004_1082, w_000_1443, w_003_060);
  or2  I004_1083(w_004_1083, w_000_1726, w_000_098);
  not1 I004_1085(w_004_1085, w_002_435);
  nand2 I004_1086(w_004_1086, w_001_797, w_003_076);
  and2 I004_1089(w_004_1089, w_000_1137, w_001_012);
  and2 I004_1090(w_004_1090, w_001_110, w_001_1233);
  not1 I004_1091(w_004_1091, w_002_321);
  and2 I004_1092(w_004_1092, w_000_890, w_003_194);
  nand2 I004_1093(w_004_1093, w_003_222, w_003_063);
  not1 I004_1094(w_004_1094, w_003_143);
  not1 I004_1095(w_004_1095, w_001_367);
  nand2 I004_1096(w_004_1096, w_002_545, w_003_080);
  and2 I004_1097(w_004_1097, w_003_308, w_002_221);
  or2  I004_1098(w_004_1098, w_003_287, w_003_139);
  and2 I004_1100(w_004_1100, w_000_1609, w_002_353);
  and2 I004_1101(w_004_1101, w_001_092, w_000_1728);
  nand2 I004_1102(w_004_1102, w_003_056, w_003_184);
  not1 I004_1105(w_004_1105, w_002_162);
  and2 I004_1107(w_004_1107, w_002_276, w_000_1107);
  nand2 I004_1108(w_004_1108, w_000_984, w_002_036);
  and2 I004_1109(w_004_1109, w_001_688, w_003_120);
  not1 I004_1110(w_004_1110, w_000_860);
  nand2 I004_1111(w_004_1111, w_001_459, w_000_1730);
  or2  I004_1112(w_004_1112, w_002_159, w_001_1661);
  not1 I004_1114(w_004_1114, w_000_191);
  or2  I004_1115(w_004_1115, w_001_1527, w_003_221);
  nand2 I004_1116(w_004_1116, w_000_909, w_003_312);
  or2  I004_1120(w_004_1120, w_003_080, w_000_1060);
  nand2 I004_1121(w_004_1121, w_001_015, w_003_289);
  not1 I004_1122(w_004_1122, w_002_221);
  nand2 I004_1123(w_004_1123, w_001_1354, w_002_501);
  not1 I004_1125(w_004_1125, w_003_031);
  not1 I004_1127(w_004_1127, w_001_638);
  not1 I004_1128(w_004_1128, w_001_894);
  nand2 I004_1130(w_004_1130, w_000_1732, w_001_1094);
  and2 I004_1132(w_004_1132, w_002_413, w_003_258);
  not1 I004_1133(w_004_1133, w_001_737);
  or2  I004_1135(w_004_1135, w_001_658, w_003_315);
  and2 I004_1136(w_004_1136, w_001_012, w_003_175);
  nand2 I004_1138(w_004_1138, w_000_714, w_003_016);
  nand2 I004_1140(w_004_1140, w_003_293, w_001_1071);
  not1 I004_1141(w_004_1141, w_002_500);
  or2  I004_1149(w_004_1149, w_000_1659, w_000_610);
  not1 I004_1150(w_004_1150, w_001_453);
  or2  I004_1151(w_004_1151, w_002_352, w_003_247);
  nand2 I004_1152(w_004_1152, w_003_089, w_003_002);
  nand2 I004_1153(w_004_1153, w_002_379, w_002_117);
  and2 I004_1157(w_004_1157, w_003_005, w_002_325);
  or2  I004_1158(w_004_1158, w_001_1212, w_000_984);
  not1 I004_1161(w_004_1161, w_003_100);
  nand2 I004_1164(w_004_1164, w_002_355, w_002_551);
  and2 I004_1166(w_004_1166, w_003_198, w_003_141);
  and2 I004_1169(w_004_1169, w_003_022, w_001_1416);
  nand2 I004_1171(w_004_1171, w_002_569, w_000_170);
  not1 I004_1174(w_004_1174, w_003_107);
  or2  I004_1177(w_004_1177, w_001_894, w_002_040);
  and2 I004_1179(w_004_1179, w_001_977, w_003_027);
  and2 I004_1180(w_004_1180, w_002_123, w_002_035);
  nand2 I004_1181(w_004_1181, w_001_494, w_002_162);
  nand2 I004_1182(w_004_1182, w_003_017, w_001_470);
  and2 I004_1184(w_004_1184, w_001_1402, w_001_850);
  and2 I004_1186(w_004_1186, w_003_065, w_000_1029);
  not1 I004_1187(w_004_1187, w_002_228);
  not1 I004_1188(w_004_1188, w_003_263);
  and2 I004_1189(w_004_1189, w_000_090, w_000_1253);
  nand2 I004_1191(w_004_1191, w_000_520, w_000_1694);
  nand2 I004_1194(w_004_1194, w_003_278, w_001_815);
  not1 I004_1197(w_004_1197, w_002_173);
  and2 I004_1200(w_004_1200, w_002_435, w_003_041);
  or2  I004_1201(w_004_1201, w_000_1176, w_003_173);
  nand2 I004_1202(w_004_1202, w_003_035, w_003_219);
  or2  I004_1204(w_004_1204, w_000_655, w_002_564);
  or2  I004_1206(w_004_1206, w_002_178, w_000_821);
  or2  I004_1207(w_004_1207, w_002_121, w_002_285);
  nand2 I004_1208(w_004_1208, w_001_460, w_002_407);
  and2 I004_1210(w_004_1210, w_002_129, w_003_252);
  nand2 I004_1211(w_004_1211, w_002_048, w_003_200);
  and2 I004_1212(w_004_1212, w_001_527, w_000_1561);
  not1 I004_1215(w_004_1215, w_003_260);
  or2  I004_1216(w_004_1216, w_000_042, w_001_1462);
  or2  I004_1217(w_004_1217, w_000_675, w_000_1558);
  and2 I004_1221(w_004_1221, w_002_498, w_001_1003);
  nand2 I004_1222(w_004_1222, w_000_033, w_002_456);
  and2 I004_1224(w_004_1224, w_001_804, w_000_012);
  not1 I004_1226(w_004_1226, w_002_164);
  nand2 I004_1228(w_004_1228, w_000_1525, w_000_939);
  and2 I004_1229(w_004_1229, w_001_1324, w_002_503);
  not1 I004_1231(w_004_1231, w_003_145);
  nand2 I004_1232(w_004_1232, w_003_262, w_002_031);
  nand2 I004_1234(w_004_1234, w_001_1486, w_001_316);
  or2  I004_1235(w_004_1235, w_001_151, w_002_234);
  or2  I004_1236(w_004_1236, w_003_152, w_003_156);
  and2 I004_1239(w_004_1239, w_002_120, w_003_286);
  and2 I004_1241(w_004_1241, w_000_353, w_002_201);
  nand2 I004_1243(w_004_1243, w_003_081, w_003_107);
  nand2 I004_1244(w_004_1244, w_000_884, w_000_808);
  nand2 I004_1248(w_004_1248, w_003_195, w_003_124);
  not1 I004_1250(w_004_1250, w_000_1736);
  or2  I004_1254(w_004_1254, w_001_674, w_001_011);
  and2 I004_1255(w_004_1255, w_000_692, w_003_107);
  and2 I004_1259(w_004_1259, w_000_529, w_001_075);
  and2 I004_1260(w_004_1260, w_002_492, w_001_1359);
  or2  I004_1263(w_004_1263, w_001_1639, w_001_653);
  not1 I004_1264(w_004_1264, w_003_094);
  not1 I004_1265(w_004_1265, w_000_071);
  and2 I004_1267(w_004_1267, w_001_908, w_003_181);
  nand2 I004_1268(w_004_1268, w_003_302, w_002_436);
  or2  I004_1269(w_004_1269, w_003_096, w_003_183);
  not1 I004_1270(w_004_1270, w_001_133);
  nand2 I004_1271(w_004_1271, w_002_151, w_002_059);
  and2 I004_1272(w_004_1272, w_003_084, w_000_1666);
  nand2 I004_1276(w_004_1276, w_002_120, w_002_209);
  not1 I004_1278(w_004_1278, w_002_329);
  not1 I004_1279(w_004_1279, w_001_1647);
  not1 I004_1280(w_004_1280, w_003_280);
  nand2 I004_1281(w_004_1281, w_000_697, w_001_261);
  or2  I004_1283(w_004_1283, w_003_141, w_003_226);
  and2 I004_1284(w_004_1284, w_000_1022, w_003_141);
  nand2 I004_1287(w_004_1287, w_000_588, w_002_400);
  or2  I004_1288(w_004_1288, w_003_053, w_002_178);
  nand2 I004_1289(w_004_1289, w_000_754, w_000_1627);
  and2 I004_1290(w_004_1290, w_003_205, w_000_1636);
  and2 I004_1291(w_004_1291, w_003_129, w_002_095);
  and2 I004_1292(w_004_1292, w_002_389, w_001_783);
  or2  I004_1293(w_004_1293, w_000_543, w_001_285);
  nand2 I004_1294(w_004_1294, w_002_004, w_000_749);
  not1 I004_1295(w_004_1295, w_000_1701);
  or2  I004_1296(w_004_1296, w_000_1328, w_001_1172);
  not1 I004_1298(w_004_1298, w_000_1609);
  not1 I004_1300(w_004_1300, w_001_068);
  not1 I004_1301(w_004_1301, w_000_1098);
  or2  I004_1302(w_004_1302, w_003_132, w_000_1187);
  or2  I004_1305(w_004_1305, w_000_895, w_002_419);
  nand2 I004_1306(w_004_1306, w_003_234, w_001_016);
  not1 I004_1310(w_004_1310, w_000_1612);
  not1 I004_1311(w_004_1311, w_000_1739);
  and2 I004_1312(w_004_1312, w_000_640, w_002_099);
  and2 I004_1315(w_004_1315, w_001_577, w_001_1085);
  not1 I004_1319(w_004_1319, w_000_452);
  not1 I004_1320(w_004_1320, w_000_1740);
  nand2 I004_1321(w_004_1321, w_000_1576, w_002_178);
  and2 I004_1322(w_004_1322, w_001_261, w_003_298);
  or2  I004_1324(w_004_1324, w_003_021, w_001_1101);
  or2  I004_1326(w_004_1326, w_001_948, w_003_102);
  not1 I004_1328(w_004_1328, w_003_077);
  or2  I004_1329(w_004_1329, w_002_193, w_001_553);
  nand2 I004_1330(w_004_1330, w_002_215, w_001_157);
  and2 I004_1335(w_004_1335, w_003_103, w_003_116);
  nand2 I004_1337(w_004_1337, w_003_032, w_000_280);
  not1 I004_1338(w_004_1338, w_002_108);
  or2  I004_1340(w_004_1340, w_003_069, w_002_138);
  nand2 I004_1344(w_004_1344, w_002_259, w_003_234);
  and2 I004_1348(w_004_1348, w_003_204, w_003_195);
  or2  I004_1349(w_004_1349, w_001_860, w_003_105);
  nand2 I004_1352(w_004_1352, w_003_055, w_000_929);
  nand2 I004_1354(w_004_1354, w_001_287, w_003_032);
  and2 I004_1356(w_004_1356, w_002_275, w_000_1317);
  or2  I004_1357(w_004_1357, w_003_107, w_000_229);
  or2  I004_1358(w_004_1358, w_003_280, w_000_1742);
  not1 I004_1361(w_004_1361, w_003_295);
  nand2 I004_1362(w_004_1362, w_001_395, w_002_493);
  and2 I004_1364(w_004_1364, w_002_180, w_000_1603);
  nand2 I004_1365(w_004_1365, w_000_1516, w_003_068);
  not1 I004_1366(w_004_1366, w_001_1456);
  or2  I004_1374(w_004_1374, w_000_1657, w_003_170);
  and2 I004_1379(w_004_1379, w_003_237, w_003_089);
  or2  I004_1380(w_004_1380, w_001_993, w_002_080);
  nand2 I004_1381(w_004_1381, w_002_123, w_002_534);
  or2  I004_1382(w_004_1382, w_002_580, w_002_523);
  or2  I004_1384(w_004_1384, w_000_422, w_000_1744);
  and2 I004_1388(w_004_1388, w_001_1462, w_001_1199);
  nand2 I004_1390(w_004_1390, w_000_1405, w_003_152);
  not1 I004_1393(w_004_1393, w_002_050);
  and2 I004_1394(w_004_1394, w_003_291, w_003_019);
  nand2 I004_1398(w_004_1398, w_000_1261, w_002_307);
  and2 I004_1399(w_004_1399, w_003_297, w_003_069);
  or2  I004_1401(w_004_1401, w_003_200, w_003_024);
  nand2 I004_1402(w_004_1402, w_003_067, w_000_635);
  or2  I004_1404(w_004_1404, w_000_632, w_002_474);
  nand2 I004_1406(w_004_1406, w_003_219, w_001_1155);
  or2  I004_1409(w_004_1409, w_003_240, w_001_746);
  nand2 I004_1410(w_004_1410, w_001_1646, w_001_589);
  or2  I004_1412(w_004_1412, w_002_030, w_001_363);
  or2  I004_1413(w_004_1413, w_000_1222, w_002_543);
  not1 I004_1414(w_004_1414, w_000_1745);
  or2  I004_1415(w_004_1415, w_002_419, w_000_391);
  not1 I004_1417(w_004_1417, w_003_132);
  nand2 I004_1418(w_004_1418, w_000_042, w_003_280);
  and2 I004_1420(w_004_1420, w_000_711, w_002_410);
  or2  I004_1422(w_004_1422, w_003_000, w_001_1230);
  nand2 I004_1423(w_004_1423, w_003_004, w_001_478);
  nand2 I004_1425(w_004_1425, w_001_225, w_001_1485);
  not1 I004_1427(w_004_1427, w_001_219);
  nand2 I004_1428(w_004_1428, w_000_820, w_000_323);
  not1 I004_1430(w_004_1430, w_000_703);
  not1 I004_1435(w_004_1435, w_002_189);
  not1 I004_1436(w_004_1436, w_002_492);
  or2  I004_1437(w_004_1437, w_002_130, w_002_565);
  and2 I004_1442(w_004_1442, w_000_1747, w_000_874);
  or2  I004_1445(w_004_1445, w_000_1748, w_003_183);
  nand2 I004_1446(w_004_1446, w_002_171, w_000_1362);
  or2  I004_1447(w_004_1447, w_000_1184, w_000_859);
  not1 I004_1448(w_004_1448, w_000_939);
  nand2 I004_1449(w_004_1449, w_001_165, w_002_449);
  and2 I004_1453(w_004_1453, w_003_104, w_001_073);
  and2 I004_1454(w_004_1454, w_001_974, w_002_042);
  not1 I004_1455(w_004_1455, w_001_123);
  nand2 I004_1456(w_004_1456, w_000_1749, w_001_170);
  and2 I004_1458(w_004_1458, w_000_1339, w_003_027);
  and2 I004_1459(w_004_1459, w_002_126, w_000_1597);
  and2 I004_1460(w_004_1460, w_002_524, w_001_221);
  and2 I004_1463(w_004_1463, w_001_1217, w_001_1556);
  or2  I004_1466(w_004_1466, w_002_102, w_001_108);
  not1 I004_1467(w_004_1467, w_002_020);
  and2 I004_1468(w_004_1468, w_002_325, w_001_137);
  not1 I004_1469(w_004_1469, w_001_1184);
  not1 I004_1470(w_004_1470, w_002_159);
  and2 I004_1472(w_004_1472, w_003_254, w_003_083);
  not1 I004_1474(w_004_1474, w_003_124);
  nand2 I004_1478(w_004_1478, w_002_327, w_003_273);
  or2  I004_1480(w_004_1480, w_000_1036, w_003_147);
  and2 I004_1481(w_004_1481, w_000_1326, w_001_822);
  and2 I004_1484(w_004_1484, w_003_192, w_000_1745);
  and2 I004_1485(w_004_1485, w_003_019, w_001_390);
  or2  I004_1487(w_004_1487, w_001_030, w_001_1057);
  and2 I004_1488(w_004_1488, w_002_097, w_002_385);
  or2  I004_1492(w_004_1492, w_001_699, w_001_580);
  nand2 I004_1493(w_004_1493, w_002_283, w_000_1447);
  or2  I004_1494(w_004_1494, w_002_504, w_001_1488);
  and2 I004_1495(w_004_1495, w_000_1061, w_003_063);
  not1 I004_1501(w_004_1501, w_000_999);
  nand2 I004_1502(w_004_1502, w_003_055, w_003_024);
  nand2 I004_1508(w_004_1508, w_003_022, w_002_258);
  not1 I004_1509(w_004_1509, w_002_062);
  or2  I004_1511(w_004_1511, w_003_062, w_001_637);
  nand2 I004_1516(w_004_1516, w_003_287, w_000_417);
  nand2 I004_1517(w_004_1517, w_001_106, w_001_047);
  nand2 I004_1519(w_004_1519, w_000_1385, w_000_431);
  or2  I004_1521(w_004_1521, w_000_1327, w_003_193);
  and2 I004_1523(w_004_1523, w_003_067, w_003_092);
  nand2 I004_1524(w_004_1524, w_001_491, w_001_787);
  or2  I004_1530(w_004_1530, w_003_166, w_000_1752);
  nand2 I004_1532(w_004_1532, w_001_389, w_000_1753);
  and2 I004_1533(w_004_1533, w_000_1754, w_001_1593);
  and2 I004_1534(w_004_1534, w_000_546, w_001_641);
  or2  I004_1535(w_004_1535, w_002_067, w_000_1473);
  or2  I004_1537(w_004_1537, w_001_223, w_003_194);
  and2 I004_1539(w_004_1539, w_003_238, w_000_499);
  and2 I004_1540(w_004_1540, w_002_445, w_000_1450);
  nand2 I004_1543(w_004_1543, w_001_1456, w_001_350);
  nand2 I004_1544(w_004_1544, w_000_1756, w_001_1039);
  not1 I004_1546(w_004_1546, w_002_340);
  nand2 I004_1547(w_004_1547, w_002_384, w_002_054);
  and2 I004_1549(w_004_1549, w_003_021, w_003_036);
  nand2 I004_1552(w_004_1552, w_003_255, w_001_729);
  or2  I004_1553(w_004_1553, w_000_257, w_000_726);
  nand2 I004_1554(w_004_1554, w_002_538, w_000_1757);
  not1 I004_1555(w_004_1555, w_003_005);
  nand2 I004_1558(w_004_1558, w_003_038, w_001_137);
  nand2 I004_1560(w_004_1560, w_003_274, w_003_081);
  not1 I004_1562(w_004_1562, w_000_1073);
  and2 I004_1563(w_004_1563, w_002_183, w_001_1096);
  nand2 I004_1565(w_004_1565, w_003_270, w_000_1175);
  and2 I004_1566(w_004_1566, w_003_152, w_000_1202);
  nand2 I004_1568(w_004_1568, w_001_1076, w_001_1061);
  not1 I004_1570(w_004_1570, w_000_1758);
  nand2 I004_1572(w_004_1572, w_001_316, w_002_211);
  and2 I004_1573(w_004_1573, w_002_288, w_000_554);
  and2 I004_1575(w_004_1575, w_001_1654, w_001_446);
  and2 I004_1576(w_004_1576, w_003_292, w_002_443);
  and2 I004_1578(w_004_1578, w_001_248, w_000_1759);
  nand2 I004_1583(w_004_1583, w_000_757, w_002_044);
  or2  I004_1589(w_004_1589, w_003_187, w_002_527);
  and2 I004_1590(w_004_1590, w_002_118, w_002_503);
  nand2 I004_1592(w_004_1592, w_001_061, w_002_472);
  or2  I004_1593(w_004_1593, w_003_227, w_003_278);
  not1 I004_1594(w_004_1594, w_002_012);
  nand2 I004_1595(w_004_1595, w_003_001, w_001_734);
  or2  I004_1596(w_004_1596, w_003_208, w_001_825);
  not1 I004_1597(w_004_1597, w_003_049);
  not1 I004_1599(w_004_1599, w_003_099);
  and2 I004_1600(w_004_1600, w_003_029, w_003_150);
  and2 I004_1601(w_004_1601, w_001_071, w_003_231);
  and2 I004_1602(w_004_1602, w_002_505, w_001_1508);
  not1 I004_1603(w_004_1603, w_001_026);
  nand2 I004_1604(w_004_1604, w_002_395, w_002_331);
  and2 I004_1605(w_004_1605, w_003_246, w_002_129);
  nand2 I004_1608(w_004_1608, w_003_248, w_000_225);
  not1 I004_1610(w_004_1610, w_002_221);
  or2  I004_1611(w_004_1611, w_000_1740, w_001_883);
  nand2 I004_1612(w_004_1612, w_003_006, w_003_212);
  and2 I004_1613(w_004_1613, w_000_1080, w_000_575);
  nand2 I004_1614(w_004_1614, w_000_1761, w_002_425);
  and2 I004_1615(w_004_1615, w_002_056, w_001_1008);
  or2  I004_1616(w_004_1616, w_000_1762, w_003_050);
  or2  I004_1618(w_004_1618, w_003_037, w_003_298);
  not1 I004_1619(w_004_1619, w_003_066);
  not1 I004_1622(w_004_1622, w_002_278);
  nand2 I004_1624(w_004_1624, w_001_1084, w_000_1587);
  and2 I004_1625(w_004_1625, w_002_340, w_003_099);
  nand2 I004_1626(w_004_1626, w_002_073, w_002_002);
  not1 I004_1631(w_004_1631, w_001_888);
  and2 I004_1633(w_004_1633, w_000_1763, w_003_127);
  not1 I004_1635(w_004_1635, w_001_1088);
  or2  I004_1636(w_004_1636, w_002_241, w_001_1436);
  or2  I004_1637(w_004_1637, w_000_484, w_000_1764);
  not1 I004_1638(w_004_1638, w_002_534);
  not1 I004_1640(w_004_1640, w_002_356);
  not1 I004_1641(w_004_1641, w_002_104);
  and2 I004_1643(w_004_1643, w_003_214, w_003_248);
  nand2 I004_1645(w_004_1645, w_001_486, w_001_1033);
  or2  I004_1647(w_004_1647, w_003_157, w_003_020);
  and2 I004_1648(w_004_1648, w_001_236, w_000_1765);
  or2  I004_1649(w_004_1649, w_001_390, w_003_165);
  and2 I004_1652(w_004_1652, w_003_183, w_001_020);
  or2  I004_1653(w_004_1653, w_002_055, w_002_156);
  and2 I004_1655(w_004_1655, w_001_1386, w_001_1098);
  and2 I004_1656(w_004_1656, w_000_223, w_002_094);
  and2 I004_1659(w_004_1659, w_001_1669, w_001_584);
  and2 I004_1660(w_004_1660, w_000_1334, w_001_965);
  and2 I004_1661(w_004_1661, w_002_496, w_000_1551);
  not1 I004_1663(w_004_1663, w_002_037);
  and2 I004_1664(w_004_1664, w_001_1428, w_000_225);
  nand2 I004_1665(w_004_1665, w_002_080, w_003_042);
  and2 I004_1667(w_004_1667, w_001_246, w_000_831);
  not1 I004_1674(w_004_1674, w_003_034);
  nand2 I004_1675(w_004_1675, w_001_233, w_002_028);
  or2  I004_1678(w_004_1678, w_000_461, w_003_296);
  not1 I004_1679(w_004_1679, w_000_1447);
  or2  I004_1681(w_004_1681, w_001_436, w_001_1515);
  and2 I004_1682(w_004_1682, w_002_560, w_002_568);
  not1 I004_1684(w_004_1684, w_000_028);
  or2  I004_1686(w_004_1686, w_000_1699, w_001_1583);
  or2  I004_1687(w_004_1687, w_003_277, w_003_076);
  not1 I004_1689(w_004_1689, w_002_089);
  and2 I004_1690(w_004_1690, w_002_539, w_000_1261);
  not1 I004_1692(w_004_1692, w_001_234);
  not1 I004_1693(w_004_1693, w_003_074);
  nand2 I004_1694(w_004_1694, w_000_210, w_002_275);
  and2 I004_1696(w_004_1696, w_001_1063, w_003_215);
  nand2 I004_1698(w_004_1698, w_000_1632, w_000_1575);
  not1 I004_1699(w_004_1699, w_002_162);
  nand2 I004_1702(w_004_1702, w_002_320, w_002_367);
  and2 I004_1703(w_004_1703, w_003_024, w_000_1486);
  nand2 I004_1706(w_004_1706, w_000_290, w_003_169);
  not1 I004_1707(w_004_1707, w_003_251);
  and2 I004_1708(w_004_1708, w_001_835, w_000_047);
  nand2 I004_1709(w_004_1709, w_002_172, w_003_234);
  not1 I004_1711(w_004_1711, w_001_1322);
  and2 I004_1712(w_004_1712, w_002_115, w_002_501);
  or2  I004_1714(w_004_1714, w_003_264, w_000_955);
  or2  I004_1716(w_004_1716, w_003_060, w_000_1325);
  and2 I004_1718(w_004_1718, w_003_088, w_000_1669);
  nand2 I004_1719(w_004_1719, w_002_522, w_001_716);
  not1 I004_1720(w_004_1720, w_003_107);
  and2 I004_1727(w_004_1727, w_000_1126, w_001_155);
  not1 I004_1731(w_004_1731, w_002_494);
  and2 I004_1732(w_004_1732, w_000_1768, w_003_106);
  and2 I004_1733(w_004_1733, w_003_022, w_000_682);
  nand2 I004_1734(w_004_1734, w_001_798, w_003_275);
  not1 I004_1737(w_004_1737, w_001_989);
  or2  I004_1739(w_004_1739, w_000_967, w_001_419);
  or2  I004_1740(w_004_1740, w_002_265, w_000_1769);
  nand2 I004_1741(w_004_1741, w_003_170, w_003_140);
  and2 I004_1742(w_004_1742, w_001_113, w_000_429);
  not1 I004_1743(w_004_1743, w_001_086);
  and2 I004_1744(w_004_1744, w_002_523, w_000_1518);
  nand2 I004_1745(w_004_1745, w_001_049, w_001_317);
  not1 I004_1746(w_004_1746, w_002_494);
  nand2 I004_1747(w_004_1747, w_000_893, w_000_187);
  or2  I004_1748(w_004_1748, w_003_070, w_000_1659);
  not1 I004_1749(w_004_1749, w_001_082);
  nand2 I004_1750(w_004_1750, w_002_420, w_000_1770);
  nand2 I004_1752(w_004_1752, w_001_459, w_000_1472);
  and2 I004_1753(w_004_1753, w_002_178, w_003_090);
  or2  I004_1755(w_004_1755, w_001_1593, w_001_276);
  nand2 I004_1756(w_004_1756, w_002_049, w_002_039);
  nand2 I004_1757(w_004_1757, w_002_185, w_002_583);
  and2 I004_1760(w_004_1760, w_002_200, w_001_1470);
  not1 I004_1765(w_004_1765, w_000_1771);
  nand2 I004_1767(w_004_1767, w_003_223, w_001_251);
  and2 I004_1769(w_004_1769, w_000_916, w_002_062);
  not1 I004_1770(w_004_1770, w_002_172);
  nand2 I004_1771(w_004_1771, w_000_1461, w_002_126);
  or2  I004_1773(w_004_1773, w_002_440, w_000_813);
  nand2 I004_1774(w_004_1774, w_001_1107, w_000_1772);
  not1 I004_1776(w_004_1776, w_000_1327);
  and2 I004_1777(w_004_1777, w_002_093, w_003_182);
  not1 I004_1778(w_004_1778, w_001_032);
  or2  I004_1780(w_004_1780, w_000_907, w_001_1430);
  not1 I004_1781(w_004_1781, w_003_249);
  nand2 I004_1782(w_004_1782, w_000_1362, w_003_318);
  and2 I004_1784(w_004_1784, w_002_550, w_003_009);
  nand2 I004_1786(w_004_1786, w_003_159, w_002_203);
  and2 I004_1787(w_004_1787, w_002_298, w_002_204);
  nand2 I004_1788(w_004_1788, w_001_1093, w_002_033);
  and2 I004_1791(w_004_1791, w_002_090, w_002_318);
  and2 I004_1792(w_004_1792, w_002_055, w_003_292);
  nand2 I004_1793(w_004_1793, w_000_026, w_003_022);
  and2 I004_1795(w_004_1795, w_000_814, w_000_217);
  or2  I004_1797(w_004_1797, w_000_1774, w_002_549);
  and2 I004_1798(w_004_1798, w_002_347, w_001_109);
  or2  I004_1799(w_004_1799, w_000_393, w_003_248);
  nand2 I004_1800(w_004_1800, w_002_402, w_002_479);
  nand2 I004_1801(w_004_1801, w_003_003, w_001_041);
  and2 I004_1802(w_004_1802, w_000_178, w_002_206);
  or2  I004_1805(w_004_1805, w_002_385, w_003_161);
  nand2 I004_1807(w_004_1807, w_002_122, w_002_353);
  and2 I004_1809(w_004_1809, w_003_301, w_001_1498);
  nand2 I004_1810(w_004_1810, w_001_677, w_003_282);
  or2  I004_1811(w_004_1811, w_001_1152, w_002_244);
  not1 I004_1812(w_004_1812, w_003_318);
  or2  I004_1814(w_004_1814, w_001_1051, w_003_317);
  not1 I004_1815(w_004_1815, w_002_051);
  nand2 I004_1817(w_004_1817, w_001_279, w_000_850);
  not1 I004_1819(w_004_1819, w_001_1585);
  and2 I004_1821(w_004_1821, w_002_465, w_000_1775);
  or2  I004_1823(w_004_1823, w_000_1648, w_000_1776);
  and2 I004_1827(w_004_1827, w_001_1605, w_003_089);
  and2 I004_1828(w_004_1828, w_000_747, w_000_1142);
  not1 I004_1829(w_004_1829, w_001_1118);
  nand2 I004_1831(w_004_1831, w_003_267, w_000_659);
  not1 I004_1832(w_004_1832, w_003_162);
  nand2 I004_1833(w_004_1833, w_000_243, w_002_122);
  and2 I004_1834(w_004_1834, w_001_696, w_001_1526);
  nand2 I004_1835(w_004_1835, w_002_286, w_000_1769);
  not1 I004_1836(w_004_1836, w_002_547);
  nand2 I004_1837(w_004_1837, w_000_1349, w_001_1456);
  not1 I004_1839(w_004_1839, w_000_1082);
  not1 I004_1840(w_004_1840, w_000_1325);
  and2 I004_1841(w_004_1841, w_001_169, w_001_1573);
  and2 I004_1843(w_004_1843, w_001_885, w_002_127);
  and2 I004_1845(w_004_1845, w_000_679, w_000_972);
  or2  I004_1848(w_004_1848, w_001_028, w_003_012);
  or2  I004_1849(w_004_1849, w_000_229, w_002_480);
  and2 I004_1850(w_004_1850, w_001_767, w_003_048);
  not1 I004_1851(w_004_1851, w_003_256);
  not1 I004_1852(w_004_1852, w_003_188);
  and2 I004_1855(w_004_1855, w_003_282, w_001_1135);
  nand2 I004_1858(w_004_1858, w_003_027, w_000_089);
  or2  I004_1860(w_004_1860, w_001_196, w_001_204);
  or2  I004_1861(w_004_1861, w_002_515, w_002_579);
  nand2 I004_1863(w_004_1863, w_003_074, w_000_694);
  and2 I004_1864(w_004_1864, w_000_822, w_000_891);
  or2  I004_1865(w_004_1865, w_000_980, w_003_232);
  or2  I004_1867(w_004_1867, w_003_032, w_001_1078);
  and2 I004_1868(w_004_1868, w_000_1448, w_001_805);
  and2 I004_1871(w_004_1871, w_003_012, w_000_414);
  and2 I004_1872(w_004_1872, w_000_683, w_002_118);
  or2  I004_1873(w_004_1873, w_003_014, w_002_234);
  and2 I004_1874(w_004_1874, w_002_117, w_000_1127);
  not1 I004_1875(w_004_1875, w_001_080);
  not1 I004_1882(w_004_1882, w_000_479);
  or2  I004_1883(w_004_1883, w_003_021, w_001_530);
  not1 I004_1884(w_004_1884, w_002_444);
  nand2 I004_1885(w_004_1885, w_000_199, w_000_1502);
  not1 I004_1886(w_004_1886, w_001_137);
  nand2 I004_1887(w_004_1887, w_002_496, w_003_206);
  or2  I004_1888(w_004_1888, w_001_901, w_001_1649);
  or2  I004_1893(w_004_1893, w_002_159, w_001_094);
  nand2 I004_1894(w_004_1894, w_002_001, w_000_951);
  or2  I004_1895(w_004_1895, w_001_976, w_000_034);
  and2 I004_1896(w_004_1896, w_001_1526, w_001_172);
  not1 I004_1899(w_004_1899, w_003_019);
  nand2 I004_1900(w_004_1900, w_001_312, w_000_1559);
  and2 I004_1902(w_004_1902, w_001_280, w_000_039);
  nand2 I004_1905(w_004_1905, w_001_253, w_003_181);
  and2 I004_1906(w_004_1906, w_002_552, w_003_127);
  or2  I004_1907(w_004_1907, w_000_359, w_001_943);
  not1 I004_1909(w_004_1909, w_003_308);
  not1 I004_1910(w_004_1910, w_002_522);
  and2 I004_1911(w_004_1911, w_000_1778, w_002_191);
  or2  I005_001(w_005_001, w_002_174, w_004_1164);
  nand2 I005_003(w_005_003, w_002_569, w_002_499);
  or2  I005_004(w_005_004, w_004_548, w_004_042);
  and2 I005_005(w_005_005, w_000_389, w_003_277);
  and2 I005_006(w_005_006, w_004_1543, w_004_1740);
  nand2 I005_008(w_005_008, w_004_451, w_003_138);
  not1 I005_009(w_005_009, w_004_407);
  or2  I005_013(w_005_013, w_000_135, w_000_585);
  not1 I005_014(w_005_014, w_001_070);
  not1 I005_015(w_005_015, w_003_103);
  or2  I005_016(w_005_016, w_004_261, w_002_393);
  not1 I005_017(w_005_017, w_001_1477);
  and2 I005_019(w_005_019, w_000_1779, w_004_596);
  and2 I005_021(w_005_021, w_001_963, w_004_003);
  or2  I005_022(w_005_022, w_004_353, w_004_1712);
  not1 I005_023(w_005_023, w_003_006);
  or2  I005_024(w_005_024, w_002_110, w_000_1574);
  and2 I005_025(w_005_025, w_004_807, w_001_1215);
  and2 I005_026(w_005_026, w_003_112, w_003_084);
  and2 I005_029(w_005_029, w_001_1065, w_002_539);
  nand2 I005_030(w_005_030, w_000_281, w_000_1656);
  and2 I005_032(w_005_032, w_004_1221, w_004_451);
  or2  I005_033(w_005_033, w_002_336, w_003_251);
  not1 I005_034(w_005_034, w_002_037);
  or2  I005_035(w_005_035, w_000_521, w_000_844);
  nand2 I005_036(w_005_036, w_002_571, w_003_204);
  and2 I005_037(w_005_037, w_003_180, w_004_448);
  and2 I005_038(w_005_038, w_001_862, w_001_623);
  nand2 I005_039(w_005_039, w_002_480, w_003_020);
  not1 I005_040(w_005_040, w_001_213);
  or2  I005_041(w_005_041, w_000_1480, w_003_048);
  not1 I005_042(w_005_042, w_000_172);
  nand2 I005_044(w_005_044, w_000_414, w_004_1568);
  nand2 I005_045(w_005_045, w_002_188, w_002_000);
  or2  I005_046(w_005_046, w_004_1427, w_004_1664);
  or2  I005_047(w_005_047, w_002_138, w_003_013);
  and2 I005_048(w_005_048, w_001_1261, w_002_201);
  or2  I005_049(w_005_049, w_003_141, w_000_855);
  nand2 I005_050(w_005_050, w_004_061, w_001_818);
  nand2 I005_051(w_005_051, w_000_548, w_002_396);
  and2 I005_052(w_005_052, w_003_269, w_002_191);
  or2  I005_053(w_005_053, w_000_400, w_000_1603);
  or2  I005_054(w_005_054, w_003_032, w_003_080);
  nand2 I005_055(w_005_055, w_003_096, w_003_003);
  nand2 I005_056(w_005_056, w_000_143, w_001_569);
  or2  I005_057(w_005_057, w_003_041, w_003_202);
  not1 I005_058(w_005_058, w_004_080);
  nand2 I005_059(w_005_059, w_001_053, w_000_498);
  not1 I005_060(w_005_060, w_001_454);
  not1 I005_065(w_005_065, w_002_555);
  or2  I005_066(w_005_066, w_000_1554, w_000_969);
  or2  I005_068(w_005_068, w_002_106, w_001_177);
  and2 I005_069(w_005_069, w_000_1056, w_003_194);
  and2 I005_070(w_005_070, w_001_976, w_000_1780);
  or2  I005_072(w_005_072, w_000_1152, w_004_001);
  or2  I005_073(w_005_073, w_001_336, w_001_568);
  and2 I005_074(w_005_074, w_002_562, w_001_1656);
  not1 I005_075(w_005_075, w_003_068);
  not1 I005_076(w_005_076, w_001_182);
  nand2 I005_077(w_005_077, w_000_1159, w_003_070);
  nand2 I005_078(w_005_078, w_000_010, w_000_412);
  and2 I005_079(w_005_079, w_000_1781, w_003_078);
  not1 I005_080(w_005_080, w_004_415);
  and2 I005_082(w_005_082, w_004_1519, w_004_501);
  nand2 I005_083(w_005_083, w_002_098, w_001_1247);
  nand2 I005_084(w_005_084, w_003_118, w_000_380);
  not1 I005_086(w_005_086, w_000_462);
  not1 I005_087(w_005_087, w_003_244);
  nand2 I005_089(w_005_089, w_003_224, w_004_071);
  and2 I005_090(w_005_090, w_001_677, w_000_650);
  or2  I005_093(w_005_093, w_003_275, w_002_196);
  or2  I005_094(w_005_094, w_003_075, w_004_1560);
  not1 I005_095(w_005_095, w_003_234);
  or2  I005_096(w_005_096, w_002_184, w_004_1189);
  not1 I005_097(w_005_097, w_002_084);
  not1 I005_098(w_005_098, w_003_230);
  and2 I005_100(w_005_100, w_003_242, w_003_158);
  and2 I005_101(w_005_101, w_000_1475, w_001_187);
  and2 I005_103(w_005_103, w_004_1423, w_000_1193);
  and2 I005_105(w_005_105, w_003_281, w_000_424);
  nand2 I005_106(w_005_106, w_002_227, w_004_1090);
  nand2 I005_109(w_005_109, w_000_1783, w_002_203);
  not1 I005_111(w_005_111, w_001_626);
  nand2 I005_112(w_005_112, w_001_1402, w_003_200);
  nand2 I005_114(w_005_114, w_004_1356, w_002_268);
  nand2 I005_115(w_005_115, w_000_985, w_003_056);
  nand2 I005_116(w_005_116, w_001_393, w_004_726);
  nand2 I005_117(w_005_117, w_003_246, w_003_224);
  and2 I005_120(w_005_120, w_002_138, w_003_111);
  not1 I005_121(w_005_121, w_003_187);
  and2 I005_123(w_005_123, w_003_002, w_001_491);
  and2 I005_124(w_005_124, w_002_199, w_002_232);
  and2 I005_125(w_005_125, w_004_1050, w_000_821);
  and2 I005_126(w_005_126, w_003_013, w_003_122);
  and2 I005_127(w_005_127, w_003_153, w_003_301);
  and2 I005_128(w_005_128, w_003_280, w_002_188);
  and2 I005_129(w_005_129, w_002_331, w_004_019);
  or2  I005_131(w_005_131, w_002_152, w_002_097);
  and2 I005_132(w_005_132, w_003_232, w_001_513);
  or2  I005_133(w_005_133, w_004_235, w_001_125);
  and2 I005_134(w_005_134, w_000_1716, w_001_998);
  not1 I005_136(w_005_136, w_002_499);
  and2 I005_137(w_005_137, w_001_1147, w_002_069);
  not1 I005_139(w_005_139, w_002_527);
  and2 I005_140(w_005_140, w_002_168, w_004_194);
  nand2 I005_142(w_005_142, w_004_146, w_004_652);
  and2 I005_143(w_005_143, w_003_051, w_001_691);
  not1 I005_144(w_005_144, w_003_107);
  and2 I005_146(w_005_146, w_003_164, w_002_069);
  or2  I005_148(w_005_148, w_003_065, w_000_1784);
  and2 I005_149(w_005_149, w_000_440, w_000_122);
  and2 I005_150(w_005_150, w_000_1166, w_000_1512);
  and2 I005_151(w_005_151, w_003_291, w_001_285);
  and2 I005_152(w_005_152, w_003_210, w_003_298);
  not1 I005_153(w_005_153, w_002_561);
  and2 I005_154(w_005_154, w_004_958, w_001_689);
  and2 I005_155(w_005_155, w_001_983, w_000_1493);
  and2 I005_156(w_005_156, w_003_048, w_002_031);
  not1 I005_158(w_005_158, w_003_060);
  not1 I005_159(w_005_159, w_003_117);
  nand2 I005_160(w_005_160, w_000_1365, w_003_166);
  and2 I005_162(w_005_162, w_001_1469, w_003_247);
  and2 I005_163(w_005_163, w_003_268, w_001_692);
  not1 I005_165(w_005_165, w_000_578);
  and2 I005_167(w_005_167, w_004_081, w_002_065);
  or2  I005_168(w_005_168, w_000_1536, w_001_162);
  or2  I005_169(w_005_169, w_001_1689, w_002_574);
  or2  I005_170(w_005_170, w_003_019, w_004_437);
  and2 I005_172(w_005_172, w_001_1325, w_003_308);
  nand2 I005_173(w_005_173, w_002_128, w_000_1785);
  nand2 I005_175(w_005_175, w_003_054, w_002_178);
  and2 I005_176(w_005_176, w_004_1201, w_002_420);
  not1 I005_178(w_005_178, w_001_156);
  and2 I005_179(w_005_179, w_001_096, w_001_1170);
  not1 I005_180(w_005_180, w_003_017);
  or2  I005_182(w_005_182, w_003_229, w_000_142);
  or2  I005_183(w_005_183, w_003_130, w_000_1149);
  or2  I005_186(w_005_186, w_004_1096, w_001_715);
  nand2 I005_187(w_005_187, w_001_196, w_004_070);
  and2 I005_188(w_005_188, w_004_1568, w_002_152);
  or2  I005_189(w_005_189, w_002_294, w_001_1627);
  and2 I005_190(w_005_190, w_001_1129, w_004_942);
  or2  I005_191(w_005_191, w_000_652, w_004_843);
  and2 I005_192(w_005_192, w_004_1815, w_000_295);
  and2 I005_194(w_005_194, w_000_1787, w_004_091);
  nand2 I005_195(w_005_195, w_002_243, w_004_1281);
  or2  I005_196(w_005_196, w_000_909, w_002_116);
  not1 I005_197(w_005_197, w_004_841);
  or2  I005_199(w_005_199, w_000_482, w_001_027);
  and2 I005_201(w_005_201, w_003_202, w_000_592);
  or2  I005_202(w_005_202, w_001_183, w_001_223);
  not1 I005_203(w_005_203, w_003_211);
  and2 I005_204(w_005_204, w_002_410, w_004_049);
  or2  I005_205(w_005_205, w_002_037, w_000_1788);
  or2  I005_206(w_005_206, w_003_021, w_002_413);
  not1 I005_207(w_005_207, w_003_158);
  nand2 I005_208(w_005_208, w_003_072, w_001_1250);
  or2  I005_209(w_005_209, w_002_529, w_000_845);
  not1 I005_212(w_005_212, w_002_026);
  and2 I005_213(w_005_213, w_000_1357, w_000_1402);
  not1 I005_216(w_005_216, w_003_292);
  and2 I005_220(w_005_220, w_002_386, w_002_113);
  or2  I005_222(w_005_222, w_000_869, w_004_1850);
  nand2 I005_223(w_005_223, w_002_266, w_004_1905);
  and2 I005_226(w_005_226, w_004_019, w_004_827);
  not1 I005_228(w_005_228, w_000_841);
  nand2 I005_229(w_005_229, w_002_062, w_003_237);
  nand2 I005_232(w_005_232, w_001_662, w_004_1777);
  nand2 I005_234(w_005_234, w_001_1402, w_000_1431);
  not1 I005_236(w_005_236, w_002_129);
  nand2 I005_237(w_005_237, w_004_1554, w_003_263);
  nand2 I005_239(w_005_239, w_002_526, w_002_575);
  nand2 I005_240(w_005_240, w_004_091, w_001_1350);
  not1 I005_242(w_005_242, w_002_556);
  or2  I005_243(w_005_243, w_004_1061, w_004_1008);
  and2 I005_244(w_005_244, w_003_024, w_003_117);
  or2  I005_245(w_005_245, w_003_178, w_003_163);
  or2  I005_246(w_005_246, w_001_1206, w_002_017);
  nand2 I005_248(w_005_248, w_000_853, w_002_480);
  and2 I005_251(w_005_251, w_001_163, w_003_129);
  nand2 I005_252(w_005_252, w_002_016, w_003_185);
  nand2 I005_253(w_005_253, w_002_568, w_001_343);
  nand2 I005_255(w_005_255, w_002_067, w_004_460);
  nand2 I005_256(w_005_256, w_004_245, w_000_1559);
  or2  I005_257(w_005_257, w_000_492, w_001_283);
  not1 I005_258(w_005_258, w_004_1095);
  not1 I005_259(w_005_259, w_000_240);
  or2  I005_260(w_005_260, w_002_214, w_002_577);
  and2 I005_261(w_005_261, w_004_700, w_004_044);
  and2 I005_262(w_005_262, w_003_143, w_002_584);
  not1 I005_263(w_005_263, w_003_175);
  not1 I005_267(w_005_267, w_002_589);
  and2 I005_268(w_005_268, w_002_036, w_003_278);
  or2  I005_269(w_005_269, w_003_009, w_003_066);
  not1 I005_271(w_005_271, w_004_1565);
  nand2 I005_272(w_005_272, w_003_143, w_001_259);
  nand2 I005_273(w_005_273, w_004_1315, w_002_492);
  or2  I005_274(w_005_274, w_001_270, w_004_975);
  and2 I005_275(w_005_275, w_002_533, w_002_040);
  not1 I005_276(w_005_276, w_002_161);
  and2 I005_278(w_005_278, w_000_1624, w_004_1460);
  and2 I005_279(w_005_279, w_000_1719, w_003_101);
  nand2 I005_280(w_005_280, w_002_320, w_000_538);
  not1 I005_281(w_005_281, w_001_1514);
  nand2 I005_283(w_005_283, w_003_254, w_001_1186);
  and2 I005_285(w_005_285, w_000_928, w_004_1125);
  and2 I005_286(w_005_286, w_001_844, w_003_183);
  nand2 I005_287(w_005_287, w_002_135, w_004_711);
  or2  I005_288(w_005_288, w_002_577, w_002_045);
  and2 I005_289(w_005_289, w_001_216, w_002_431);
  and2 I005_290(w_005_290, w_000_864, w_004_588);
  not1 I005_292(w_005_292, w_002_580);
  not1 I005_293(w_005_293, w_003_317);
  not1 I005_294(w_005_294, w_000_312);
  not1 I005_295(w_005_295, w_003_149);
  and2 I005_296(w_005_296, w_002_008, w_004_606);
  not1 I005_298(w_005_298, w_001_718);
  not1 I005_299(w_005_299, w_000_1658);
  nand2 I005_300(w_005_300, w_002_129, w_003_013);
  or2  I005_302(w_005_302, w_001_276, w_001_260);
  and2 I005_303(w_005_303, w_001_1176, w_002_427);
  or2  I005_305(w_005_305, w_003_060, w_002_485);
  not1 I005_306(w_005_306, w_004_737);
  or2  I005_307(w_005_307, w_001_1001, w_004_1841);
  not1 I005_308(w_005_308, w_002_113);
  not1 I005_309(w_005_309, w_004_1750);
  and2 I005_310(w_005_310, w_000_863, w_001_342);
  and2 I005_313(w_005_313, w_000_1464, w_003_169);
  nand2 I005_314(w_005_314, w_003_214, w_001_190);
  not1 I005_315(w_005_315, w_004_101);
  and2 I005_316(w_005_316, w_001_200, w_000_487);
  not1 I005_317(w_005_317, w_002_587);
  nand2 I005_318(w_005_318, w_000_1324, w_004_645);
  or2  I005_319(w_005_319, w_000_1790, w_004_1401);
  nand2 I005_320(w_005_320, w_004_866, w_004_774);
  or2  I005_321(w_005_321, w_004_1660, w_002_019);
  not1 I005_322(w_005_322, w_001_213);
  not1 I005_323(w_005_323, w_000_455);
  or2  I005_328(w_005_328, w_003_271, w_000_1430);
  and2 I005_331(w_005_331, w_000_615, w_003_181);
  nand2 I005_333(w_005_333, w_000_058, w_000_1791);
  nand2 I005_338(w_005_338, w_000_1118, w_004_1809);
  nand2 I005_339(w_005_339, w_003_011, w_001_1130);
  or2  I005_341(w_005_341, w_001_527, w_002_243);
  and2 I005_344(w_005_344, w_004_762, w_001_728);
  not1 I005_346(w_005_346, w_004_804);
  or2  I005_348(w_005_348, w_003_086, w_002_061);
  nand2 I005_357(w_005_357, w_002_154, w_002_346);
  or2  I005_362(w_005_362, w_000_771, w_004_031);
  or2  I005_363(w_005_363, w_000_539, w_004_1675);
  and2 I005_366(w_005_366, w_004_774, w_004_1071);
  or2  I005_368(w_005_368, w_001_1371, w_004_683);
  not1 I005_369(w_005_369, w_000_628);
  not1 I005_371(w_005_371, w_004_534);
  not1 I005_375(w_005_375, w_000_292);
  nand2 I005_376(w_005_376, w_000_1430, w_003_061);
  or2  I005_377(w_005_377, w_003_261, w_002_213);
  or2  I005_378(w_005_378, w_002_108, w_001_1664);
  and2 I005_379(w_005_379, w_002_263, w_001_1628);
  and2 I005_381(w_005_381, w_003_229, w_003_091);
  and2 I005_385(w_005_385, w_002_188, w_002_158);
  nand2 I005_386(w_005_386, w_003_288, w_002_011);
  not1 I005_387(w_005_387, w_004_1043);
  nand2 I005_390(w_005_390, w_002_118, w_002_219);
  and2 I005_394(w_005_394, w_002_472, w_000_297);
  nand2 I005_395(w_005_395, w_000_1382, w_001_1356);
  or2  I005_398(w_005_398, w_000_1713, w_001_115);
  or2  I005_400(w_005_400, w_000_803, w_003_165);
  not1 I005_402(w_005_402, w_004_1469);
  or2  I005_406(w_005_406, w_000_1792, w_002_556);
  not1 I005_408(w_005_408, w_001_026);
  or2  I005_409(w_005_409, w_004_199, w_002_214);
  or2  I005_411(w_005_411, w_003_170, w_000_1453);
  and2 I005_415(w_005_415, w_000_1244, w_002_454);
  not1 I005_420(w_005_420, w_004_201);
  nand2 I005_423(w_005_423, w_000_930, w_003_281);
  and2 I005_425(w_005_425, w_004_778, w_000_1318);
  and2 I005_428(w_005_428, w_001_665, w_000_119);
  and2 I005_430(w_005_430, w_002_114, w_000_1299);
  or2  I005_433(w_005_433, w_002_461, w_001_657);
  and2 I005_434(w_005_434, w_003_260, w_001_1646);
  or2  I005_438(w_005_438, w_004_183, w_004_1774);
  nand2 I005_439(w_005_439, w_004_1837, w_003_048);
  nand2 I005_444(w_005_444, w_001_199, w_003_141);
  and2 I005_446(w_005_446, w_003_201, w_003_122);
  nand2 I005_449(w_005_449, w_001_030, w_004_1572);
  and2 I005_453(w_005_453, w_002_295, w_001_099);
  nand2 I005_457(w_005_457, w_004_503, w_001_890);
  nand2 I005_458(w_005_458, w_001_910, w_004_1300);
  nand2 I005_459(w_005_459, w_002_363, w_000_050);
  and2 I005_460(w_005_460, w_000_375, w_004_1357);
  or2  I005_461(w_005_461, w_001_1200, w_003_274);
  not1 I005_465(w_005_465, w_004_009);
  not1 I005_466(w_005_466, w_001_880);
  and2 I005_472(w_005_472, w_004_078, w_003_318);
  and2 I005_473(w_005_473, w_001_956, w_000_1398);
  nand2 I005_477(w_005_477, w_002_539, w_004_816);
  nand2 I005_478(w_005_478, w_002_220, w_004_345);
  not1 I005_479(w_005_479, w_003_192);
  nand2 I005_484(w_005_484, w_001_1500, w_003_303);
  and2 I005_485(w_005_485, w_004_1289, w_000_1462);
  not1 I005_487(w_005_487, w_000_302);
  not1 I005_488(w_005_488, w_004_1001);
  and2 I005_490(w_005_490, w_000_357, w_002_001);
  nand2 I005_494(w_005_494, w_004_513, w_000_1074);
  not1 I005_496(w_005_496, w_003_158);
  not1 I005_497(w_005_497, w_003_195);
  not1 I005_500(w_005_500, w_002_170);
  not1 I005_501(w_005_501, w_003_049);
  or2  I005_503(w_005_503, w_004_372, w_004_1553);
  nand2 I005_504(w_005_504, w_004_1702, w_001_294);
  and2 I005_505(w_005_505, w_004_1640, w_000_1749);
  not1 I005_506(w_005_506, w_001_1424);
  not1 I005_508(w_005_508, w_002_029);
  and2 I005_511(w_005_511, w_002_449, w_002_026);
  not1 I005_523(w_005_523, w_002_113);
  and2 I005_525(w_005_525, w_004_886, w_002_493);
  not1 I005_527(w_005_527, w_003_052);
  nand2 I005_528(w_005_528, w_002_250, w_004_1656);
  not1 I005_529(w_005_529, w_001_997);
  and2 I005_530(w_005_530, w_000_1403, w_004_931);
  and2 I005_532(w_005_532, w_002_152, w_001_861);
  or2  I005_533(w_005_533, w_003_299, w_004_1241);
  not1 I005_534(w_005_534, w_000_1293);
  or2  I005_535(w_005_535, w_004_1895, w_003_066);
  not1 I005_537(w_005_537, w_000_386);
  and2 I005_538(w_005_538, w_003_109, w_000_1041);
  and2 I005_539(w_005_539, w_000_1425, w_000_553);
  not1 I005_541(w_005_541, w_001_650);
  nand2 I005_542(w_005_542, w_004_120, w_002_477);
  not1 I005_543(w_005_543, w_000_1267);
  not1 I005_544(w_005_544, w_003_157);
  and2 I005_546(w_005_546, w_003_305, w_003_126);
  nand2 I005_548(w_005_548, w_002_010, w_002_489);
  not1 I005_551(w_005_551, w_002_571);
  nand2 I005_555(w_005_555, w_001_104, w_003_185);
  or2  I005_556(w_005_556, w_000_1371, w_003_273);
  nand2 I005_559(w_005_559, w_003_104, w_004_1810);
  or2  I005_560(w_005_560, w_002_022, w_004_1706);
  and2 I005_562(w_005_562, w_001_207, w_001_559);
  or2  I005_564(w_005_564, w_002_200, w_002_353);
  or2  I005_565(w_005_565, w_003_259, w_000_824);
  or2  I005_570(w_005_570, w_001_564, w_001_1159);
  not1 I005_574(w_005_574, w_004_1157);
  not1 I005_576(w_005_576, w_001_681);
  not1 I005_577(w_005_577, w_001_1682);
  or2  I005_578(w_005_578, w_000_081, w_002_184);
  or2  I005_580(w_005_580, w_001_509, w_001_372);
  and2 I005_584(w_005_584, w_003_034, w_004_371);
  and2 I005_585(w_005_585, w_001_804, w_003_022);
  or2  I005_586(w_005_586, w_002_165, w_003_282);
  or2  I005_591(w_005_591, w_001_586, w_004_027);
  nand2 I005_593(w_005_593, w_004_1066, w_004_973);
  or2  I005_594(w_005_594, w_000_1428, w_004_599);
  not1 I005_596(w_005_596, w_001_507);
  or2  I005_597(w_005_597, w_000_1204, w_001_1074);
  not1 I005_598(w_005_598, w_001_519);
  or2  I005_599(w_005_599, w_004_1280, w_003_039);
  or2  I005_600(w_005_600, w_004_246, w_000_681);
  and2 I005_602(w_005_602, w_001_312, w_004_388);
  nand2 I005_605(w_005_605, w_002_132, w_003_016);
  not1 I005_608(w_005_608, w_002_551);
  nand2 I005_610(w_005_610, w_002_371, w_001_792);
  or2  I005_611(w_005_611, w_001_1503, w_004_1047);
  nand2 I005_612(w_005_612, w_004_1773, w_002_028);
  nand2 I005_617(w_005_617, w_000_509, w_002_205);
  nand2 I005_619(w_005_619, w_003_304, w_003_062);
  and2 I005_620(w_005_620, w_004_730, w_002_547);
  and2 I005_622(w_005_622, w_001_1204, w_001_258);
  nand2 I005_623(w_005_623, w_000_1797, w_004_1493);
  or2  I005_624(w_005_624, w_001_1480, w_001_184);
  or2  I005_625(w_005_625, w_002_291, w_000_088);
  or2  I005_627(w_005_627, w_003_257, w_001_805);
  and2 I005_628(w_005_628, w_002_261, w_000_145);
  and2 I005_630(w_005_630, w_000_820, w_002_419);
  or2  I005_632(w_005_632, w_004_1741, w_002_264);
  nand2 I005_633(w_005_633, w_000_1232, w_003_156);
  nand2 I005_636(w_005_636, w_000_287, w_004_130);
  and2 I005_638(w_005_638, w_004_229, w_004_1180);
  not1 I005_640(w_005_640, w_001_174);
  and2 I005_642(w_005_642, w_002_385, w_001_1541);
  not1 I005_643(w_005_643, w_003_028);
  nand2 I005_644(w_005_644, w_003_040, w_004_080);
  and2 I005_645(w_005_645, w_002_234, w_000_1238);
  nand2 I005_647(w_005_647, w_003_068, w_003_023);
  or2  I005_650(w_005_650, w_002_489, w_001_1470);
  or2  I005_651(w_005_651, w_000_1800, w_003_259);
  nand2 I005_652(w_005_652, w_000_778, w_004_257);
  nand2 I005_653(w_005_653, w_000_1421, w_003_188);
  or2  I005_654(w_005_654, w_001_1523, w_004_1534);
  not1 I005_655(w_005_655, w_004_1321);
  nand2 I005_658(w_005_658, w_000_245, w_003_090);
  and2 I005_659(w_005_659, w_000_868, w_004_1742);
  or2  I005_661(w_005_661, w_000_1323, w_003_071);
  or2  I005_662(w_005_662, w_004_352, w_002_368);
  or2  I005_663(w_005_663, w_001_163, w_001_1606);
  not1 I005_665(w_005_665, w_004_905);
  and2 I005_668(w_005_668, w_004_1570, w_001_1550);
  and2 I005_669(w_005_669, w_000_1801, w_004_1222);
  and2 I005_670(w_005_670, w_000_1737, w_000_1802);
  and2 I005_671(w_005_671, w_001_297, w_003_031);
  not1 I005_672(w_005_672, w_004_217);
  and2 I005_673(w_005_673, w_000_1217, w_000_1244);
  and2 I005_674(w_005_674, w_001_1491, w_003_076);
  or2  I005_675(w_005_675, w_004_1226, w_003_280);
  nand2 I005_677(w_005_677, w_002_332, w_004_860);
  nand2 I005_680(w_005_680, w_001_953, w_001_1071);
  not1 I005_682(w_005_682, w_003_289);
  and2 I005_686(w_005_686, w_000_816, w_003_288);
  or2  I005_687(w_005_687, w_001_000, w_003_192);
  and2 I005_694(w_005_694, w_004_483, w_003_162);
  or2  I005_695(w_005_695, w_001_239, w_004_899);
  and2 I005_697(w_005_697, w_000_1142, w_002_003);
  nand2 I005_699(w_005_699, w_000_972, w_000_995);
  and2 I005_702(w_005_702, w_003_083, w_004_876);
  not1 I005_706(w_005_706, w_000_571);
  or2  I005_707(w_005_707, w_003_049, w_004_528);
  not1 I005_708(w_005_708, w_002_349);
  and2 I005_709(w_005_709, w_002_192, w_003_137);
  and2 I005_712(w_005_712, w_003_292, w_004_1025);
  not1 I005_713(w_005_713, w_004_1596);
  nand2 I005_717(w_005_717, w_000_1803, w_002_142);
  or2  I005_722(w_005_722, w_002_152, w_001_414);
  nand2 I005_728(w_005_728, w_001_895, w_003_079);
  and2 I005_729(w_005_729, w_000_1613, w_002_143);
  not1 I005_730(w_005_730, w_001_1513);
  not1 I005_731(w_005_731, w_004_395);
  not1 I005_732(w_005_732, w_004_1485);
  or2  I005_733(w_005_733, w_004_544, w_003_062);
  nand2 I005_734(w_005_734, w_004_1418, w_002_516);
  not1 I005_736(w_005_736, w_001_175);
  or2  I005_738(w_005_738, w_004_973, w_002_069);
  nand2 I005_741(w_005_741, w_004_1747, w_001_1106);
  or2  I005_742(w_005_742, w_003_301, w_003_237);
  nand2 I005_747(w_005_747, w_003_181, w_003_247);
  and2 I005_748(w_005_748, w_002_212, w_000_1060);
  or2  I005_752(w_005_752, w_002_524, w_004_504);
  and2 I005_753(w_005_753, w_002_114, w_004_185);
  nand2 I005_756(w_005_756, w_002_311, w_001_362);
  or2  I005_758(w_005_758, w_001_852, w_001_1028);
  and2 I005_759(w_005_759, w_000_1532, w_001_708);
  not1 I005_760(w_005_760, w_000_1245);
  or2  I005_765(w_005_765, w_002_140, w_000_137);
  or2  I005_766(w_005_766, w_001_1197, w_001_218);
  or2  I005_768(w_005_768, w_004_1232, w_002_147);
  not1 I005_769(w_005_769, w_001_241);
  or2  I005_770(w_005_770, w_004_1509, w_001_807);
  not1 I005_771(w_005_771, w_002_513);
  not1 I005_774(w_005_774, w_000_1394);
  not1 I005_775(w_005_775, w_001_099);
  or2  I005_777(w_005_777, w_002_211, w_004_1208);
  nand2 I005_778(w_005_778, w_001_835, w_001_294);
  or2  I005_780(w_005_780, w_003_123, w_003_037);
  or2  I005_781(w_005_781, w_004_391, w_004_036);
  nand2 I005_782(w_005_782, w_003_076, w_002_031);
  not1 I005_785(w_005_785, w_001_1046);
  not1 I005_786(w_005_786, w_003_259);
  nand2 I005_787(w_005_787, w_004_1294, w_002_096);
  not1 I005_789(w_005_789, w_001_022);
  not1 I005_790(w_005_790, w_003_177);
  not1 I005_791(w_005_791, w_004_1626);
  not1 I005_793(w_005_793, w_002_285);
  or2  I005_794(w_005_794, w_000_1755, w_004_109);
  not1 I005_796(w_005_796, w_004_727);
  or2  I005_797(w_005_797, w_002_535, w_004_1560);
  nand2 I005_798(w_005_798, w_001_655, w_004_1340);
  nand2 I005_800(w_005_800, w_001_1446, w_001_1240);
  not1 I005_801(w_005_801, w_001_1485);
  and2 I005_802(w_005_802, w_003_309, w_002_410);
  nand2 I005_808(w_005_808, w_001_1020, w_002_409);
  or2  I005_809(w_005_809, w_004_1765, w_004_892);
  nand2 I005_811(w_005_811, w_004_1053, w_004_046);
  and2 I005_812(w_005_812, w_001_358, w_004_1077);
  nand2 I005_816(w_005_816, w_004_024, w_001_141);
  or2  I005_817(w_005_817, w_002_559, w_002_513);
  not1 I005_823(w_005_823, w_004_293);
  not1 I005_824(w_005_824, w_003_166);
  or2  I005_825(w_005_825, w_000_1552, w_000_1079);
  or2  I005_830(w_005_830, w_002_389, w_000_1313);
  and2 I005_832(w_005_832, w_000_1386, w_002_531);
  and2 I005_838(w_005_838, w_004_001, w_003_068);
  not1 I005_839(w_005_839, w_003_094);
  or2  I005_840(w_005_840, w_000_840, w_003_276);
  and2 I005_841(w_005_841, w_002_444, w_003_129);
  or2  I005_842(w_005_842, w_004_565, w_000_991);
  or2  I005_844(w_005_844, w_001_1046, w_000_385);
  nand2 I005_845(w_005_845, w_003_085, w_004_264);
  nand2 I005_849(w_005_849, w_003_264, w_002_248);
  nand2 I005_850(w_005_850, w_001_019, w_004_1056);
  or2  I005_851(w_005_851, w_002_546, w_002_278);
  nand2 I005_853(w_005_853, w_002_100, w_000_803);
  and2 I005_856(w_005_856, w_002_088, w_001_985);
  nand2 I005_857(w_005_857, w_004_1004, w_003_025);
  or2  I005_858(w_005_858, w_002_249, w_004_560);
  or2  I005_860(w_005_860, w_002_178, w_002_131);
  not1 I005_862(w_005_862, w_001_265);
  not1 I005_863(w_005_863, w_000_395);
  and2 I005_864(w_005_864, w_000_1619, w_004_175);
  not1 I005_872(w_005_872, w_001_1483);
  nand2 I005_873(w_005_873, w_000_719, w_001_1439);
  and2 I005_875(w_005_875, w_001_511, w_001_1365);
  and2 I005_876(w_005_876, w_001_1109, w_004_1494);
  and2 I005_880(w_005_880, w_003_277, w_001_122);
  nand2 I005_882(w_005_882, w_002_166, w_001_1023);
  or2  I005_883(w_005_883, w_002_349, w_000_1804);
  and2 I005_886(w_005_886, w_001_752, w_001_1582);
  nand2 I005_890(w_005_890, w_001_049, w_001_937);
  and2 I005_891(w_005_891, w_001_915, w_001_1532);
  nand2 I005_893(w_005_893, w_002_473, w_003_224);
  not1 I005_894(w_005_894, w_002_168);
  nand2 I005_897(w_005_897, w_000_1705, w_002_208);
  not1 I005_898(w_005_898, w_000_1717);
  nand2 I005_901(w_005_901, w_003_166, w_004_1232);
  nand2 I005_905(w_005_905, w_004_1181, w_003_001);
  and2 I005_907(w_005_907, w_000_720, w_001_1514);
  and2 I005_910(w_005_910, w_004_216, w_003_166);
  or2  I005_911(w_005_911, w_000_324, w_000_124);
  nand2 I005_912(w_005_912, w_002_117, w_003_268);
  and2 I005_914(w_005_914, w_003_197, w_003_008);
  not1 I005_915(w_005_915, w_004_1664);
  nand2 I005_917(w_005_917, w_001_1585, w_001_1441);
  or2  I005_919(w_005_919, w_000_1222, w_004_022);
  nand2 I005_922(w_005_922, w_002_276, w_004_991);
  not1 I005_924(w_005_924, w_002_589);
  and2 I005_926(w_005_926, w_001_1143, w_002_413);
  not1 I005_929(w_005_929, w_004_021);
  not1 I005_930(w_005_930, w_004_1636);
  not1 I005_932(w_005_932, w_004_316);
  not1 I005_933(w_005_933, w_000_849);
  not1 I005_934(w_005_934, w_000_028);
  not1 I005_937(w_005_937, w_001_624);
  or2  I005_943(w_005_943, w_000_047, w_002_131);
  or2  I005_944(w_005_944, w_002_074, w_003_086);
  or2  I005_949(w_005_949, w_000_1674, w_004_900);
  or2  I005_951(w_005_951, w_001_776, w_003_178);
  and2 I005_952(w_005_952, w_002_164, w_003_114);
  or2  I005_953(w_005_953, w_000_260, w_003_117);
  not1 I005_954(w_005_954, w_002_044);
  nand2 I005_955(w_005_955, w_002_065, w_004_797);
  not1 I005_959(w_005_959, w_001_526);
  nand2 I005_960(w_005_960, w_001_786, w_002_205);
  and2 I005_961(w_005_961, w_000_1789, w_000_842);
  or2  I005_962(w_005_962, w_001_302, w_004_827);
  nand2 I005_965(w_005_965, w_000_031, w_004_195);
  or2  I005_966(w_005_966, w_000_721, w_002_140);
  nand2 I005_967(w_005_967, w_004_722, w_001_1661);
  and2 I005_970(w_005_970, w_004_409, w_003_071);
  not1 I005_971(w_005_971, w_004_446);
  not1 I005_973(w_005_973, w_004_1107);
  or2  I005_974(w_005_974, w_001_181, w_003_237);
  and2 I005_975(w_005_975, w_002_373, w_004_1784);
  nand2 I005_977(w_005_977, w_001_961, w_003_244);
  nand2 I005_979(w_005_979, w_003_152, w_003_034);
  not1 I005_982(w_005_982, w_001_685);
  nand2 I005_984(w_005_984, w_003_315, w_001_722);
  and2 I005_986(w_005_986, w_001_683, w_001_511);
  and2 I005_988(w_005_988, w_000_1417, w_002_252);
  not1 I005_993(w_005_993, w_004_898);
  or2  I005_994(w_005_994, w_002_463, w_004_908);
  or2  I005_995(w_005_995, w_001_264, w_000_365);
  nand2 I005_997(w_005_997, w_001_1061, w_004_472);
  or2  I005_999(w_005_999, w_001_308, w_003_057);
  not1 I005_1002(w_005_1002, w_000_954);
  and2 I005_1005(w_005_1005, w_001_597, w_004_319);
  not1 I005_1006(w_005_1006, w_002_075);
  not1 I005_1007(w_005_1007, w_004_003);
  not1 I005_1010(w_005_1010, w_000_1730);
  or2  I005_1011(w_005_1011, w_004_176, w_002_070);
  and2 I005_1015(w_005_1015, w_004_135, w_002_120);
  nand2 I005_1019(w_005_1019, w_000_1809, w_000_901);
  not1 I005_1022(w_005_1022, w_002_357);
  or2  I005_1023(w_005_1023, w_002_119, w_000_1551);
  not1 I005_1025(w_005_1025, w_002_202);
  not1 I005_1026(w_005_1026, w_004_1910);
  and2 I005_1027(w_005_1027, w_000_1553, w_002_306);
  and2 I005_1028(w_005_1028, w_003_246, w_002_423);
  or2  I005_1033(w_005_1033, w_000_1392, w_000_1021);
  nand2 I005_1034(w_005_1034, w_002_330, w_002_052);
  not1 I005_1035(w_005_1035, w_000_776);
  or2  I005_1038(w_005_1038, w_001_1097, w_003_111);
  nand2 I005_1041(w_005_1041, w_000_1810, w_000_1811);
  or2  I005_1043(w_005_1043, w_001_1559, w_002_314);
  nand2 I005_1044(w_005_1044, w_000_165, w_004_1171);
  not1 I005_1045(w_005_1045, w_002_172);
  nand2 I005_1047(w_005_1047, w_002_108, w_001_1488);
  not1 I005_1050(w_005_1050, w_000_273);
  or2  I005_1052(w_005_1052, w_004_343, w_001_700);
  not1 I005_1056(w_005_1056, w_004_328);
  and2 I005_1057(w_005_1057, w_003_247, w_000_1671);
  and2 I005_1058(w_005_1058, w_000_456, w_003_136);
  or2  I005_1059(w_005_1059, w_004_1120, w_003_009);
  nand2 I005_1061(w_005_1061, w_003_279, w_000_1647);
  not1 I005_1065(w_005_1065, w_000_482);
  not1 I005_1070(w_005_1070, w_000_643);
  or2  I005_1074(w_005_1074, w_001_096, w_002_528);
  and2 I005_1075(w_005_1075, w_000_1480, w_004_975);
  not1 I005_1076(w_005_1076, w_004_1863);
  or2  I005_1077(w_005_1077, w_004_506, w_004_1459);
  or2  I005_1078(w_005_1078, w_001_345, w_003_205);
  or2  I005_1079(w_005_1079, w_003_290, w_002_168);
  nand2 I005_1080(w_005_1080, w_004_1733, w_003_122);
  and2 I005_1081(w_005_1081, w_000_1565, w_003_260);
  or2  I005_1082(w_005_1082, w_004_868, w_003_038);
  or2  I005_1087(w_005_1087, w_004_300, w_002_400);
  and2 I005_1088(w_005_1088, w_004_963, w_002_039);
  or2  I005_1090(w_005_1090, w_004_406, w_003_072);
  nand2 I005_1092(w_005_1092, w_000_250, w_001_567);
  nand2 I005_1093(w_005_1093, w_000_1812, w_000_337);
  nand2 I005_1094(w_005_1094, w_003_176, w_000_660);
  nand2 I005_1098(w_005_1098, w_003_316, w_004_921);
  and2 I005_1099(w_005_1099, w_002_176, w_004_1592);
  or2  I005_1100(w_005_1100, w_002_246, w_004_107);
  or2  I005_1101(w_005_1101, w_000_623, w_001_232);
  and2 I005_1102(w_005_1102, w_000_1813, w_001_008);
  not1 I005_1103(w_005_1103, w_000_650);
  not1 I005_1105(w_005_1105, w_003_026);
  not1 I005_1106(w_005_1106, w_000_1814);
  and2 I005_1109(w_005_1109, w_000_984, w_003_067);
  or2  I005_1112(w_005_1112, w_002_130, w_004_1544);
  not1 I005_1113(w_005_1113, w_001_303);
  and2 I005_1114(w_005_1114, w_002_142, w_001_370);
  and2 I005_1115(w_005_1115, w_003_314, w_001_629);
  not1 I005_1116(w_005_1116, w_001_145);
  or2  I005_1117(w_005_1117, w_003_303, w_003_065);
  not1 I005_1118(w_005_1118, w_004_987);
  and2 I005_1119(w_005_1119, w_000_992, w_004_060);
  nand2 I005_1121(w_005_1121, w_000_1069, w_002_106);
  or2  I005_1123(w_005_1123, w_001_005, w_004_017);
  nand2 I005_1125(w_005_1125, w_004_1097, w_002_387);
  or2  I005_1126(w_005_1126, w_004_1379, w_003_094);
  and2 I005_1129(w_005_1129, w_000_210, w_003_187);
  nand2 I005_1130(w_005_1130, w_004_220, w_000_1815);
  or2  I005_1132(w_005_1132, w_000_1103, w_000_1816);
  and2 I005_1133(w_005_1133, w_004_1576, w_003_279);
  not1 I005_1134(w_005_1134, w_002_456);
  not1 I005_1136(w_005_1136, w_003_227);
  or2  I005_1137(w_005_1137, w_000_1119, w_003_106);
  not1 I005_1138(w_005_1138, w_001_1240);
  and2 I005_1139(w_005_1139, w_000_1138, w_004_1384);
  and2 I005_1140(w_005_1140, w_000_908, w_001_698);
  nand2 I005_1141(w_005_1141, w_002_105, w_001_303);
  or2  I005_1142(w_005_1142, w_001_059, w_000_1066);
  or2  I005_1143(w_005_1143, w_003_045, w_003_213);
  not1 I005_1147(w_005_1147, w_002_378);
  or2  I005_1149(w_005_1149, w_000_114, w_001_321);
  nand2 I005_1150(w_005_1150, w_004_166, w_000_1378);
  not1 I005_1151(w_005_1151, w_001_904);
  nand2 I005_1152(w_005_1152, w_001_1063, w_004_269);
  not1 I005_1153(w_005_1153, w_004_633);
  or2  I005_1157(w_005_1157, w_001_078, w_002_180);
  or2  I005_1158(w_005_1158, w_000_1695, w_004_711);
  and2 I005_1159(w_005_1159, w_004_1638, w_002_405);
  nand2 I005_1160(w_005_1160, w_001_268, w_003_051);
  and2 I005_1163(w_005_1163, w_003_064, w_003_030);
  or2  I005_1165(w_005_1165, w_003_213, w_001_440);
  or2  I005_1166(w_005_1166, w_001_499, w_003_294);
  not1 I005_1167(w_005_1167, w_003_145);
  or2  I005_1168(w_005_1168, w_002_257, w_001_1120);
  or2  I005_1171(w_005_1171, w_000_585, w_004_493);
  nand2 I005_1173(w_005_1173, w_001_095, w_003_055);
  or2  I005_1175(w_005_1175, w_004_1633, w_001_342);
  or2  I005_1178(w_005_1178, w_000_1302, w_000_1817);
  nand2 I005_1180(w_005_1180, w_004_315, w_003_077);
  and2 I005_1181(w_005_1181, w_004_671, w_001_1235);
  or2  I005_1182(w_005_1182, w_001_1290, w_004_1906);
  and2 I005_1185(w_005_1185, w_003_122, w_003_040);
  and2 I005_1186(w_005_1186, w_004_1404, w_003_064);
  or2  I005_1187(w_005_1187, w_003_073, w_004_1409);
  not1 I005_1189(w_005_1189, w_004_012);
  not1 I005_1190(w_005_1190, w_000_609);
  and2 I005_1197(w_005_1197, w_004_054, w_001_241);
  nand2 I005_1199(w_005_1199, w_003_241, w_002_338);
  nand2 I005_1205(w_005_1205, w_002_593, w_002_055);
  nand2 I005_1209(w_005_1209, w_004_292, w_004_1123);
  or2  I005_1211(w_005_1211, w_000_1343, w_002_051);
  or2  I005_1213(w_005_1213, w_001_308, w_001_1278);
  or2  I005_1216(w_005_1216, w_000_1818, w_000_026);
  not1 I005_1217(w_005_1217, w_004_1435);
  nand2 I005_1218(w_005_1218, w_000_778, w_001_068);
  or2  I005_1219(w_005_1219, w_002_536, w_003_060);
  and2 I005_1220(w_005_1220, w_004_1291, w_003_178);
  nand2 I005_1222(w_005_1222, w_000_1609, w_002_033);
  or2  I005_1223(w_005_1223, w_002_194, w_001_1312);
  or2  I005_1224(w_005_1224, w_003_309, w_001_044);
  or2  I005_1228(w_005_1228, w_000_663, w_003_127);
  nand2 I005_1229(w_005_1229, w_001_422, w_000_1819);
  nand2 I005_1233(w_005_1233, w_002_056, w_002_389);
  or2  I005_1234(w_005_1234, w_003_101, w_001_1066);
  or2  I005_1235(w_005_1235, w_001_505, w_001_1617);
  nand2 I005_1237(w_005_1237, w_000_448, w_003_126);
  nand2 I005_1239(w_005_1239, w_001_237, w_004_048);
  or2  I005_1243(w_005_1243, w_001_300, w_004_1150);
  or2  I005_1251(w_005_1251, w_003_124, w_004_276);
  or2  I005_1252(w_005_1252, w_001_264, w_001_815);
  and2 I005_1254(w_005_1254, w_000_1821, w_004_818);
  not1 I005_1255(w_005_1255, w_002_297);
  or2  I005_1257(w_005_1257, w_000_455, w_003_134);
  nand2 I005_1258(w_005_1258, w_002_214, w_004_453);
  and2 I005_1259(w_005_1259, w_000_1621, w_001_530);
  or2  I005_1261(w_005_1261, w_001_200, w_002_242);
  not1 I005_1264(w_005_1264, w_002_062);
  and2 I005_1265(w_005_1265, w_003_228, w_001_214);
  or2  I005_1266(w_005_1266, w_004_1096, w_000_1822);
  and2 I005_1267(w_005_1267, w_004_1063, w_003_197);
  not1 I005_1268(w_005_1268, w_002_587);
  or2  I005_1271(w_005_1271, w_003_256, w_004_213);
  and2 I005_1274(w_005_1274, w_004_1290, w_000_073);
  or2  I005_1276(w_005_1276, w_000_1677, w_004_1909);
  nand2 I005_1278(w_005_1278, w_004_1608, w_003_214);
  or2  I005_1281(w_005_1281, w_000_1318, w_003_072);
  and2 I005_1283(w_005_1283, w_001_733, w_000_421);
  nand2 I005_1285(w_005_1285, w_003_283, w_003_126);
  not1 I005_1286(w_005_1286, w_001_137);
  and2 I005_1288(w_005_1288, w_001_734, w_004_1098);
  and2 I005_1289(w_005_1289, w_003_038, w_004_346);
  and2 I005_1292(w_005_1292, w_000_1296, w_002_336);
  nand2 I005_1293(w_005_1293, w_000_913, w_003_195);
  not1 I005_1296(w_005_1296, w_001_897);
  and2 I005_1297(w_005_1297, w_004_1311, w_000_821);
  nand2 I005_1298(w_005_1298, w_001_455, w_004_261);
  and2 I005_1300(w_005_1300, w_001_1314, w_001_1547);
  and2 I005_1303(w_005_1303, w_001_004, w_001_416);
  or2  I005_1304(w_005_1304, w_000_1118, w_002_236);
  and2 I005_1307(w_005_1307, w_002_330, w_001_1575);
  or2  I005_1308(w_005_1308, w_000_548, w_001_482);
  not1 I005_1309(w_005_1309, w_004_066);
  nand2 I005_1310(w_005_1310, w_000_396, w_000_632);
  not1 I005_1315(w_005_1315, w_000_1430);
  or2  I005_1317(w_005_1317, w_000_350, w_000_1823);
  nand2 I005_1321(w_005_1321, w_000_1824, w_003_100);
  and2 I005_1322(w_005_1322, w_003_105, w_001_1019);
  or2  I005_1324(w_005_1324, w_000_818, w_001_419);
  not1 I005_1328(w_005_1328, w_001_1203);
  not1 I005_1329(w_005_1329, w_004_1648);
  not1 I005_1330(w_005_1330, w_000_106);
  nand2 I005_1331(w_005_1331, w_003_197, w_003_124);
  or2  I005_1336(w_005_1336, w_004_088, w_004_1141);
  not1 I005_1337(w_005_1337, w_001_605);
  nand2 I005_1346(w_005_1346, w_003_021, w_004_1534);
  and2 I005_1347(w_005_1347, w_000_1168, w_002_135);
  or2  I005_1348(w_005_1348, w_003_298, w_003_074);
  nand2 I005_1349(w_005_1349, w_002_131, w_002_313);
  nand2 I005_1353(w_005_1353, w_000_334, w_003_120);
  and2 I005_1355(w_005_1355, w_003_185, w_002_141);
  or2  I005_1357(w_005_1357, w_002_036, w_000_1063);
  and2 I005_1358(w_005_1358, w_001_715, w_001_165);
  not1 I005_1360(w_005_1360, w_002_194);
  or2  I005_1362(w_005_1362, w_000_1192, w_000_1739);
  nand2 I005_1364(w_005_1364, w_001_746, w_003_073);
  nand2 I005_1366(w_005_1366, w_002_146, w_002_294);
  not1 I005_1368(w_005_1368, w_000_1158);
  nand2 I005_1369(w_005_1369, w_002_566, w_003_175);
  not1 I005_1370(w_005_1370, w_002_218);
  and2 I005_1374(w_005_1374, w_003_053, w_003_138);
  nand2 I005_1376(w_005_1376, w_003_019, w_001_655);
  and2 I005_1379(w_005_1379, w_001_617, w_000_843);
  not1 I005_1380(w_005_1380, w_000_671);
  nand2 I005_1381(w_005_1381, w_003_121, w_004_1111);
  and2 I005_1384(w_005_1384, w_000_1397, w_003_022);
  nand2 I005_1385(w_005_1385, w_000_511, w_002_386);
  nand2 I005_1392(w_005_1392, w_001_525, w_003_028);
  nand2 I005_1393(w_005_1393, w_001_899, w_001_003);
  or2  I005_1394(w_005_1394, w_002_199, w_004_908);
  nand2 I005_1397(w_005_1397, w_002_274, w_003_150);
  not1 I005_1398(w_005_1398, w_003_006);
  and2 I005_1404(w_005_1404, w_003_037, w_004_611);
  nand2 I005_1408(w_005_1408, w_000_482, w_004_1595);
  and2 I005_1409(w_005_1409, w_003_273, w_002_562);
  and2 I005_1410(w_005_1410, w_001_466, w_001_1633);
  and2 I005_1415(w_005_1415, w_002_540, w_003_292);
  and2 I005_1418(w_005_1418, w_002_249, w_002_547);
  not1 I005_1420(w_005_1420, w_000_1262);
  not1 I005_1421(w_005_1421, w_002_125);
  not1 I005_1422(w_005_1422, w_004_1428);
  and2 I005_1424(w_005_1424, w_003_263, w_004_477);
  not1 I005_1426(w_005_1426, w_002_396);
  and2 I005_1428(w_005_1428, w_002_374, w_004_1158);
  not1 I005_1429(w_005_1429, w_003_270);
  and2 I005_1430(w_005_1430, w_001_142, w_002_344);
  and2 I005_1431(w_005_1431, w_002_227, w_000_650);
  or2  I005_1436(w_005_1436, w_002_473, w_001_1413);
  nand2 I005_1439(w_005_1439, w_003_201, w_003_004);
  or2  I005_1440(w_005_1440, w_001_054, w_001_668);
  and2 I005_1441(w_005_1441, w_001_539, w_003_196);
  and2 I005_1443(w_005_1443, w_003_003, w_000_1103);
  nand2 I005_1445(w_005_1445, w_000_1076, w_004_215);
  and2 I005_1446(w_005_1446, w_001_481, w_004_1480);
  or2  I005_1447(w_005_1447, w_002_465, w_003_161);
  or2  I005_1448(w_005_1448, w_002_008, w_004_388);
  nand2 I005_1449(w_005_1449, w_003_006, w_000_1826);
  not1 I005_1450(w_005_1450, w_000_119);
  nand2 I005_1451(w_005_1451, w_000_1362, w_001_1350);
  and2 I005_1461(w_005_1461, w_002_220, w_004_1792);
  or2  I005_1464(w_005_1464, w_003_028, w_001_231);
  not1 I005_1467(w_005_1467, w_004_1745);
  or2  I005_1469(w_005_1469, w_001_045, w_000_1250);
  nand2 I005_1470(w_005_1470, w_002_313, w_004_1896);
  or2  I005_1473(w_005_1473, w_004_1302, w_002_049);
  or2  I005_1478(w_005_1478, w_003_004, w_002_100);
  nand2 I005_1480(w_005_1480, w_004_1867, w_003_288);
  not1 I005_1485(w_005_1485, w_002_138);
  nand2 I005_1487(w_005_1487, w_000_715, w_004_616);
  and2 I005_1491(w_005_1491, w_000_116, w_002_030);
  not1 I005_1492(w_005_1492, w_002_352);
  not1 I005_1493(w_005_1493, w_004_054);
  or2  I005_1494(w_005_1494, w_001_683, w_003_002);
  or2  I005_1495(w_005_1495, w_003_158, w_002_172);
  and2 I005_1499(w_005_1499, w_001_856, w_004_1902);
  nand2 I005_1501(w_005_1501, w_004_694, w_003_228);
  nand2 I005_1505(w_005_1505, w_001_1215, w_002_126);
  and2 I005_1511(w_005_1511, w_000_557, w_004_1043);
  not1 I005_1513(w_005_1513, w_004_162);
  or2  I005_1519(w_005_1519, w_004_117, w_000_1705);
  nand2 I005_1522(w_005_1522, w_003_108, w_002_397);
  nand2 I005_1523(w_005_1523, w_001_059, w_001_709);
  or2  I005_1525(w_005_1525, w_004_1819, w_003_070);
  and2 I005_1526(w_005_1526, w_003_007, w_001_1101);
  or2  I005_1528(w_005_1528, w_004_396, w_001_538);
  and2 I005_1529(w_005_1529, w_002_394, w_001_110);
  or2  I005_1533(w_005_1533, w_002_434, w_001_1317);
  and2 I005_1534(w_005_1534, w_000_661, w_000_591);
  and2 I005_1536(w_005_1536, w_000_1470, w_002_559);
  or2  I005_1538(w_005_1538, w_002_582, w_002_300);
  or2  I005_1540(w_005_1540, w_000_1058, w_003_075);
  and2 I005_1542(w_005_1542, w_004_1745, w_003_111);
  or2  I005_1548(w_005_1548, w_000_1381, w_004_305);
  and2 I005_1549(w_005_1549, w_001_998, w_003_097);
  or2  I005_1550(w_005_1550, w_003_285, w_000_615);
  nand2 I005_1551(w_005_1551, w_004_042, w_002_537);
  nand2 I005_1553(w_005_1553, w_000_1106, w_000_1830);
  not1 I005_1554(w_005_1554, w_004_1260);
  nand2 I005_1557(w_005_1557, w_000_232, w_004_1884);
  or2  I005_1558(w_005_1558, w_003_087, w_000_295);
  nand2 I005_1560(w_005_1560, w_003_037, w_003_279);
  not1 I005_1561(w_005_1561, w_002_120);
  and2 I005_1562(w_005_1562, w_000_1035, w_002_302);
  nand2 I005_1566(w_005_1566, w_003_172, w_002_370);
  nand2 I005_1569(w_005_1569, w_002_460, w_002_137);
  and2 I005_1572(w_005_1572, w_001_704, w_002_149);
  nand2 I005_1574(w_005_1574, w_003_068, w_003_033);
  and2 I005_1575(w_005_1575, w_004_785, w_003_111);
  nand2 I005_1576(w_005_1576, w_002_396, w_004_925);
  or2  I005_1577(w_005_1577, w_002_122, w_001_217);
  not1 I005_1579(w_005_1579, w_000_172);
  nand2 I005_1580(w_005_1580, w_000_1044, w_004_609);
  nand2 I005_1581(w_005_1581, w_004_277, w_003_232);
  or2  I005_1582(w_005_1582, w_002_055, w_003_109);
  and2 I005_1584(w_005_1584, w_002_313, w_000_1566);
  not1 I005_1587(w_005_1587, w_002_374);
  or2  I005_1588(w_005_1588, w_002_191, w_004_096);
  nand2 I005_1591(w_005_1591, w_000_419, w_000_1685);
  not1 I005_1592(w_005_1592, w_001_1529);
  or2  I005_1593(w_005_1593, w_001_270, w_002_210);
  and2 I005_1596(w_005_1596, w_002_540, w_002_548);
  nand2 I005_1597(w_005_1597, w_000_209, w_003_267);
  nand2 I005_1602(w_005_1602, w_002_153, w_002_088);
  or2  I005_1603(w_005_1603, w_001_411, w_003_239);
  and2 I005_1605(w_005_1605, w_003_068, w_001_1028);
  and2 I005_1609(w_005_1609, w_003_063, w_000_1831);
  nand2 I005_1610(w_005_1610, w_003_008, w_000_1560);
  and2 I005_1612(w_005_1612, w_004_031, w_000_324);
  or2  I005_1613(w_005_1613, w_003_318, w_003_143);
  not1 I005_1616(w_005_1616, w_000_415);
  or2  I005_1617(w_005_1617, w_000_424, w_001_247);
  and2 I005_1619(w_005_1619, w_000_930, w_001_349);
  nand2 I005_1620(w_005_1620, w_000_1832, w_002_038);
  and2 I005_1622(w_005_1622, w_004_1049, w_003_216);
  nand2 I005_1624(w_005_1624, w_004_807, w_004_803);
  or2  I005_1626(w_005_1626, w_004_1409, w_003_056);
  nand2 I005_1628(w_005_1628, w_002_413, w_003_228);
  nand2 I005_1631(w_005_1631, w_002_397, w_003_180);
  and2 I005_1636(w_005_1636, w_002_365, w_002_154);
  or2  I005_1637(w_005_1637, w_000_1833, w_004_1202);
  not1 I005_1638(w_005_1638, w_002_374);
  or2  I005_1639(w_005_1639, w_000_1278, w_003_184);
  and2 I005_1641(w_005_1641, w_003_220, w_003_307);
  nand2 I005_1645(w_005_1645, w_002_430, w_003_057);
  nand2 I005_1646(w_005_1646, w_002_316, w_004_1295);
  or2  I005_1650(w_005_1650, w_003_069, w_003_036);
  nand2 I005_1651(w_005_1651, w_002_219, w_001_889);
  not1 I005_1652(w_005_1652, w_004_546);
  or2  I005_1653(w_005_1653, w_004_862, w_001_994);
  not1 I005_1656(w_005_1656, w_000_459);
  and2 I005_1658(w_005_1658, w_003_208, w_004_1324);
  and2 I005_1662(w_005_1662, w_002_382, w_002_202);
  not1 I005_1663(w_005_1663, w_002_419);
  or2  I005_1664(w_005_1664, w_002_580, w_002_056);
  not1 I005_1666(w_005_1666, w_004_772);
  or2  I005_1667(w_005_1667, w_004_1858, w_004_1840);
  nand2 I005_1668(w_005_1668, w_001_485, w_003_018);
  or2  I005_1669(w_005_1669, w_003_034, w_002_539);
  and2 I005_1672(w_005_1672, w_003_186, w_001_1044);
  and2 I005_1674(w_005_1674, w_003_013, w_002_322);
  not1 I006_000(w_006_000, w_005_226);
  and2 I006_001(w_006_001, w_002_394, w_001_049);
  and2 I006_002(w_006_002, w_005_316, w_000_1350);
  nand2 I006_003(w_006_003, w_003_242, w_000_1756);
  or2  I006_004(w_006_004, w_004_1707, w_000_307);
  and2 I006_005(w_006_005, w_005_1639, w_004_766);
  or2  I006_006(w_006_006, w_002_444, w_005_1056);
  and2 I006_007(w_006_007, w_001_606, w_000_1835);
  nand2 I006_008(w_006_008, w_005_890, w_003_007);
  and2 I006_009(w_006_009, w_003_249, w_002_087);
  or2  I006_010(w_006_010, w_001_1035, w_004_1532);
  not1 I006_011(w_006_011, w_004_1357);
  not1 I006_012(w_006_012, w_000_124);
  nand2 I006_013(w_006_013, w_000_1514, w_000_1808);
  not1 I006_014(w_006_014, w_000_767);
  and2 I006_015(w_006_015, w_002_586, w_001_520);
  or2  I006_017(w_006_017, w_000_619, w_000_085);
  not1 I006_018(w_006_018, w_003_149);
  not1 I006_019(w_006_019, w_000_081);
  and2 I006_020(w_006_020, w_002_437, w_004_977);
  or2  I006_021(w_006_021, w_002_193, w_002_142);
  or2  I006_022(w_006_022, w_001_228, w_002_351);
  and2 I006_023(w_006_023, w_002_395, w_001_881);
  not1 I006_024(w_006_024, w_001_1500);
  and2 I006_025(w_006_025, w_000_226, w_002_181);
  or2  I006_026(w_006_026, w_002_020, w_005_984);
  nand2 I006_027(w_006_027, w_001_313, w_000_1447);
  and2 I006_028(w_006_028, w_000_535, w_000_059);
  nand2 I006_029(w_006_029, w_000_1836, w_001_218);
  and2 I006_030(w_006_030, w_002_263, w_001_373);
  nand2 I006_031(w_006_031, w_001_405, w_000_085);
  not1 I006_032(w_006_032, w_005_1587);
  and2 I006_033(w_006_033, w_004_571, w_003_309);
  and2 I006_034(w_006_034, w_004_108, w_003_194);
  nand2 I006_035(w_006_035, w_001_254, w_004_233);
  or2  I006_036(w_006_036, w_000_803, w_001_040);
  nand2 I006_038(w_006_038, w_004_1793, w_002_509);
  or2  I006_039(w_006_039, w_002_383, w_004_1674);
  and2 I006_040(w_006_040, w_003_006, w_002_582);
  and2 I006_041(w_006_041, w_001_1201, w_004_1094);
  not1 I006_042(w_006_042, w_005_708);
  or2  I006_043(w_006_043, w_005_1100, w_000_109);
  not1 I006_044(w_006_044, w_001_127);
  not1 I006_045(w_006_045, w_005_288);
  and2 I006_046(w_006_046, w_001_006, w_000_1222);
  and2 I006_047(w_006_047, w_004_1455, w_005_170);
  nand2 I006_048(w_006_048, w_003_003, w_005_245);
  or2  I006_049(w_006_049, w_003_106, w_005_1285);
  and2 I006_050(w_006_050, w_004_385, w_000_1543);
  and2 I006_051(w_006_051, w_001_023, w_000_203);
  and2 I006_052(w_006_052, w_004_206, w_004_064);
  and2 I006_053(w_006_053, w_000_309, w_001_1026);
  nand2 I006_054(w_006_054, w_005_070, w_002_162);
  not1 I006_055(w_006_055, w_002_145);
  and2 I006_056(w_006_056, w_001_024, w_004_1635);
  or2  I006_057(w_006_057, w_005_1178, w_001_1280);
  nand2 I006_058(w_006_058, w_005_160, w_005_501);
  or2  I006_059(w_006_059, w_003_278, w_004_1776);
  nand2 I006_060(w_006_060, w_003_194, w_002_548);
  nand2 I006_061(w_006_061, w_003_250, w_003_153);
  or2  I006_062(w_006_062, w_000_1634, w_005_1366);
  or2  I006_063(w_006_063, w_003_031, w_005_1492);
  and2 I006_064(w_006_064, w_005_500, w_005_1666);
  or2  I006_065(w_006_065, w_005_662, w_001_323);
  not1 I006_066(w_006_066, w_004_1380);
  and2 I006_067(w_006_067, w_001_1469, w_003_178);
  nand2 I006_068(w_006_068, w_005_283, w_003_083);
  or2  I006_069(w_006_069, w_002_581, w_002_553);
  or2  I006_070(w_006_070, w_005_046, w_003_156);
  not1 I006_071(w_006_071, w_000_1103);
  nand2 I006_072(w_006_072, w_005_117, w_001_1020);
  nand2 I006_073(w_006_073, w_005_753, w_001_986);
  not1 I006_074(w_006_074, w_002_054);
  or2  I006_075(w_006_075, w_001_119, w_002_210);
  and2 I006_076(w_006_076, w_003_012, w_004_334);
  or2  I006_077(w_006_077, w_004_732, w_000_1108);
  not1 I006_078(w_006_078, w_000_211);
  not1 I006_079(w_006_079, w_000_328);
  or2  I006_080(w_006_080, w_004_1235, w_000_201);
  not1 I006_081(w_006_081, w_005_423);
  or2  I006_082(w_006_082, w_005_717, w_004_777);
  nand2 I006_083(w_006_083, w_003_237, w_004_1187);
  and2 I006_084(w_006_084, w_005_632, w_004_1271);
  not1 I006_085(w_006_085, w_000_1254);
  and2 I006_086(w_006_086, w_004_1136, w_000_1820);
  or2  I006_087(w_006_087, w_003_128, w_003_006);
  not1 I006_088(w_006_088, w_002_508);
  nand2 I006_089(w_006_089, w_002_037, w_004_1279);
  not1 I006_090(w_006_090, w_001_1148);
  nand2 I006_091(w_006_091, w_004_1296, w_004_706);
  and2 I006_092(w_006_092, w_003_232, w_003_263);
  and2 I006_093(w_006_093, w_001_1351, w_001_061);
  and2 I006_094(w_006_094, w_004_1821, w_002_004);
  and2 I006_095(w_006_095, w_002_294, w_001_726);
  or2  I006_096(w_006_096, w_003_037, w_004_918);
  not1 I006_097(w_006_097, w_003_032);
  not1 I006_098(w_006_098, w_005_023);
  nand2 I006_099(w_006_099, w_002_328, w_000_1318);
  nand2 I006_100(w_006_100, w_005_669, w_004_1322);
  not1 I006_101(w_006_101, w_000_1496);
  not1 I006_102(w_006_102, w_004_1868);
  not1 I006_103(w_006_103, w_003_283);
  or2  I006_104(w_006_104, w_004_1659, w_004_1366);
  or2  I006_105(w_006_105, w_000_873, w_002_263);
  not1 I006_106(w_006_106, w_000_886);
  or2  I006_107(w_006_107, w_001_216, w_003_298);
  nand2 I006_108(w_006_108, w_000_1722, w_005_1426);
  and2 I006_109(w_006_109, w_005_045, w_002_205);
  nand2 I006_110(w_006_110, w_003_201, w_000_1770);
  and2 I006_111(w_006_111, w_004_1488, w_003_243);
  not1 I006_112(w_006_112, w_003_138);
  and2 I006_113(w_006_113, w_002_156, w_001_267);
  not1 I006_114(w_006_114, w_002_017);
  or2  I006_115(w_006_115, w_001_1279, w_000_1837);
  nand2 I006_116(w_006_116, w_000_052, w_001_153);
  nand2 I006_117(w_006_117, w_003_034, w_003_243);
  not1 I006_118(w_006_118, w_001_051);
  and2 I006_119(w_006_119, w_004_765, w_003_170);
  not1 I006_120(w_006_120, w_003_154);
  nand2 I006_121(w_006_121, w_004_1756, w_004_1791);
  or2  I006_122(w_006_122, w_005_1070, w_002_134);
  or2  I006_123(w_006_123, w_000_780, w_001_589);
  nand2 I006_124(w_006_124, w_004_576, w_002_165);
  not1 I006_125(w_006_125, w_002_216);
  not1 I006_126(w_006_126, w_004_014);
  not1 I006_127(w_006_127, w_005_1126);
  or2  I006_128(w_006_128, w_005_1577, w_004_078);
  or2  I006_129(w_006_129, w_003_315, w_002_538);
  nand2 I006_130(w_006_130, w_001_503, w_005_004);
  not1 I006_131(w_006_131, w_003_111);
  not1 I006_132(w_006_132, w_003_285);
  or2  I006_133(w_006_133, w_001_207, w_002_462);
  not1 I006_134(w_006_134, w_000_068);
  or2  I006_135(w_006_135, w_000_345, w_004_655);
  nand2 I006_137(w_006_137, w_005_1163, w_000_094);
  nand2 I006_138(w_006_138, w_004_353, w_002_039);
  nand2 I006_139(w_006_139, w_003_230, w_003_136);
  and2 I006_140(w_006_140, w_003_230, w_002_349);
  not1 I006_141(w_006_141, w_003_179);
  and2 I006_142(w_006_142, w_005_786, w_003_238);
  nand2 I006_143(w_006_143, w_002_082, w_005_013);
  or2  I006_144(w_006_144, w_005_460, w_002_117);
  or2  I006_145(w_006_145, w_004_884, w_004_1305);
  nand2 I006_146(w_006_146, w_001_1074, w_003_102);
  and2 I006_147(w_006_147, w_005_1443, w_003_052);
  not1 I006_148(w_006_148, w_003_165);
  or2  I006_149(w_006_149, w_004_355, w_002_149);
  or2  I006_150(w_006_150, w_001_296, w_001_113);
  and2 I006_151(w_006_151, w_001_364, w_001_636);
  or2  I006_152(w_006_152, w_000_1838, w_004_1295);
  nand2 I006_153(w_006_153, w_001_038, w_000_1288);
  or2  I006_154(w_006_154, w_001_012, w_000_634);
  or2  I006_155(w_006_155, w_003_174, w_005_049);
  or2  I006_156(w_006_156, w_002_145, w_004_265);
  not1 I006_157(w_006_157, w_002_021);
  not1 I006_158(w_006_158, w_004_1845);
  nand2 I006_159(w_006_159, w_002_138, w_001_1053);
  not1 I006_160(w_006_160, w_000_1443);
  not1 I006_161(w_006_161, w_002_089);
  or2  I006_162(w_006_162, w_004_1037, w_001_776);
  not1 I006_163(w_006_163, w_001_653);
  nand2 I006_164(w_006_164, w_001_507, w_004_249);
  or2  I006_165(w_006_165, w_004_783, w_000_1289);
  nand2 I006_166(w_006_166, w_005_189, w_005_317);
  and2 I006_167(w_006_167, w_005_175, w_000_550);
  or2  I006_168(w_006_168, w_003_179, w_002_177);
  and2 I006_169(w_006_169, w_001_735, w_000_515);
  and2 I006_170(w_006_170, w_000_1338, w_000_1839);
  nand2 I006_171(w_006_171, w_005_305, w_000_1355);
  not1 I006_172(w_006_172, w_002_346);
  not1 I006_173(w_006_173, w_005_176);
  not1 I006_174(w_006_174, w_004_379);
  or2  I006_175(w_006_175, w_005_1436, w_004_1260);
  nand2 I006_176(w_006_176, w_003_189, w_002_047);
  nand2 I006_177(w_006_177, w_003_289, w_003_133);
  or2  I006_178(w_006_178, w_000_1672, w_000_489);
  nand2 I006_179(w_006_179, w_005_787, w_003_127);
  or2  I006_180(w_006_180, w_000_1840, w_000_1367);
  not1 I006_182(w_006_182, w_005_060);
  or2  I006_183(w_006_183, w_000_1241, w_004_1809);
  or2  I006_184(w_006_184, w_005_1379, w_004_815);
  and2 I006_185(w_006_185, w_002_487, w_003_015);
  not1 I006_186(w_006_186, w_002_208);
  nand2 I006_187(w_006_187, w_004_1752, w_002_591);
  and2 I006_188(w_006_188, w_001_1253, w_005_707);
  nand2 I006_189(w_006_189, w_002_525, w_003_304);
  or2  I006_190(w_006_190, w_005_1394, w_000_980);
  or2  I006_191(w_006_191, w_002_013, w_001_027);
  nand2 I006_192(w_006_192, w_002_394, w_005_1289);
  or2  I006_193(w_006_193, w_001_259, w_005_086);
  and2 I006_194(w_006_194, w_003_020, w_003_102);
  nand2 I006_195(w_006_195, w_002_456, w_004_1061);
  not1 I006_196(w_006_196, w_003_000);
  and2 I006_197(w_006_197, w_001_293, w_001_1274);
  and2 I006_198(w_006_198, w_001_1653, w_001_1239);
  nand2 I006_199(w_006_199, w_001_528, w_002_032);
  or2  I006_200(w_006_200, w_005_252, w_003_218);
  nand2 I006_201(w_006_201, w_004_1312, w_000_067);
  not1 I006_202(w_006_202, w_004_1480);
  or2  I006_203(w_006_203, w_000_793, w_001_1261);
  not1 I006_204(w_006_204, w_003_215);
  not1 I006_205(w_006_205, w_002_540);
  not1 I006_206(w_006_206, w_003_268);
  nand2 I006_207(w_006_207, w_002_184, w_003_043);
  not1 I006_208(w_006_208, w_000_085);
  and2 I006_209(w_006_209, w_003_031, w_005_1317);
  not1 I006_210(w_006_210, w_005_893);
  nand2 I006_211(w_006_211, w_004_1733, w_000_406);
  nand2 I006_212(w_006_212, w_000_1841, w_004_046);
  or2  I006_214(w_006_214, w_004_1547, w_004_1718);
  or2  I006_215(w_006_215, w_002_021, w_000_697);
  not1 I006_216(w_006_216, w_003_014);
  or2  I006_217(w_006_217, w_002_072, w_002_063);
  or2  I006_218(w_006_218, w_002_009, w_000_110);
  not1 I006_219(w_006_219, w_003_102);
  or2  I006_220(w_006_220, w_004_985, w_003_041);
  not1 I006_221(w_006_221, w_002_260);
  or2  I006_222(w_006_222, w_000_1242, w_005_457);
  and2 I006_223(w_006_223, w_003_243, w_001_387);
  and2 I006_224(w_006_224, w_003_047, w_004_1652);
  or2  I006_225(w_006_225, w_000_013, w_003_258);
  nand2 I006_226(w_006_226, w_000_633, w_004_1610);
  not1 I006_227(w_006_227, w_002_323);
  and2 I006_228(w_006_228, w_002_584, w_005_1652);
  not1 I006_229(w_006_229, w_005_461);
  not1 I006_230(w_006_230, w_002_430);
  or2  I006_231(w_006_231, w_005_065, w_004_1009);
  or2  I006_232(w_006_232, w_001_354, w_004_300);
  nand2 I006_233(w_006_233, w_002_316, w_004_377);
  and2 I006_234(w_006_234, w_000_347, w_000_1290);
  and2 I006_235(w_006_235, w_000_226, w_005_564);
  and2 I006_236(w_006_236, w_002_431, w_004_264);
  not1 I006_237(w_006_237, w_005_1626);
  nand2 I006_238(w_006_238, w_003_027, w_004_1612);
  or2  I006_239(w_006_239, w_000_1842, w_004_1883);
  or2  I006_240(w_006_240, w_000_612, w_003_103);
  and2 I006_241(w_006_241, w_004_993, w_000_204);
  nand2 I006_242(w_006_242, w_003_161, w_001_352);
  not1 I006_243(w_006_243, w_003_296);
  and2 I006_244(w_006_244, w_002_242, w_005_1505);
  or2  I006_245(w_006_245, w_002_524, w_002_462);
  nand2 I006_246(w_006_246, w_005_697, w_004_095);
  not1 I006_247(w_006_247, w_001_150);
  not1 I006_248(w_006_248, w_003_215);
  not1 I006_249(w_006_249, w_000_714);
  nand2 I006_250(w_006_250, w_003_081, w_003_265);
  not1 I006_251(w_006_251, w_000_1118);
  not1 I006_252(w_006_252, w_002_001);
  and2 I006_253(w_006_253, w_000_1513, w_000_826);
  and2 I006_254(w_006_254, w_001_143, w_005_1385);
  or2  I006_255(w_006_255, w_001_1430, w_001_1309);
  and2 I006_256(w_006_256, w_001_303, w_002_399);
  nand2 I006_257(w_006_257, w_005_387, w_004_246);
  or2  I006_258(w_006_258, w_002_528, w_000_1521);
  not1 I006_259(w_006_259, w_004_1425);
  nand2 I006_260(w_006_260, w_002_251, w_001_359);
  or2  I006_261(w_006_261, w_001_096, w_002_460);
  not1 I006_262(w_006_262, w_001_080);
  not1 I006_263(w_006_263, w_002_425);
  and2 I006_264(w_006_264, w_000_1136, w_003_201);
  nand2 I006_265(w_006_265, w_000_078, w_003_036);
  not1 I006_266(w_006_266, w_004_1614);
  not1 I006_267(w_006_267, w_005_386);
  and2 I006_268(w_006_268, w_005_1485, w_005_496);
  not1 I006_269(w_006_269, w_003_286);
  nand2 I006_270(w_006_270, w_002_473, w_001_876);
  and2 I006_271(w_006_271, w_002_537, w_000_107);
  not1 I006_272(w_006_272, w_001_1418);
  not1 I006_273(w_006_273, w_005_1575);
  nand2 I006_274(w_006_274, w_004_044, w_005_934);
  or2  I006_275(w_006_275, w_001_831, w_004_1413);
  not1 I006_276(w_006_276, w_000_1023);
  not1 I006_277(w_006_277, w_004_1446);
  and2 I006_278(w_006_278, w_002_209, w_000_154);
  not1 I006_279(w_006_279, w_005_101);
  or2  I006_280(w_006_280, w_002_317, w_001_1582);
  and2 I006_281(w_006_281, w_002_563, w_004_1076);
  nand2 I006_282(w_006_282, w_005_842, w_000_570);
  not1 I006_283(w_006_283, w_001_008);
  nand2 I006_284(w_006_284, w_001_502, w_003_221);
  not1 I006_285(w_006_285, w_005_1205);
  nand2 I006_286(w_006_286, w_001_519, w_004_813);
  and2 I006_287(w_006_287, w_004_076, w_001_1263);
  or2  I006_288(w_006_288, w_001_420, w_005_003);
  nand2 I006_289(w_006_289, w_004_520, w_002_018);
  not1 I006_290(w_006_290, w_001_379);
  or2  I006_291(w_006_291, w_000_881, w_003_110);
  and2 I006_292(w_006_292, w_002_321, w_003_040);
  not1 I006_293(w_006_293, w_005_133);
  not1 I006_294(w_006_294, w_004_210);
  or2  I006_295(w_006_295, w_003_155, w_000_1615);
  and2 I006_296(w_006_296, w_000_735, w_001_712);
  or2  I006_297(w_006_297, w_001_251, w_002_428);
  and2 I006_298(w_006_298, w_003_256, w_001_079);
  and2 I006_299(w_006_299, w_002_090, w_003_162);
  not1 I006_300(w_006_300, w_002_021);
  and2 I006_301(w_006_301, w_000_1177, w_005_058);
  and2 I006_302(w_006_302, w_003_069, w_003_208);
  and2 I006_303(w_006_303, w_002_232, w_003_097);
  nand2 I006_304(w_006_304, w_005_112, w_000_538);
  and2 I006_305(w_006_305, w_005_307, w_004_1301);
  nand2 I006_306(w_006_306, w_001_135, w_003_045);
  nand2 I006_307(w_006_307, w_003_264, w_002_096);
  or2  I006_308(w_006_308, w_003_214, w_004_394);
  not1 I006_309(w_006_309, w_002_488);
  not1 I006_310(w_006_310, w_005_1577);
  not1 I006_311(w_006_311, w_003_089);
  not1 I006_312(w_006_312, w_003_089);
  or2  I006_313(w_006_313, w_005_170, w_001_392);
  and2 I006_314(w_006_314, w_004_558, w_000_1733);
  nand2 I006_315(w_006_315, w_000_366, w_004_1287);
  nand2 I006_316(w_006_316, w_002_470, w_003_122);
  and2 I006_317(w_006_317, w_005_013, w_004_102);
  not1 I006_318(w_006_318, w_005_144);
  and2 I006_319(w_006_319, w_002_553, w_000_1477);
  nand2 I006_320(w_006_320, w_001_180, w_003_199);
  and2 I006_321(w_006_321, w_003_285, w_001_053);
  nand2 I006_322(w_006_322, w_003_103, w_002_481);
  or2  I006_323(w_006_323, w_005_1103, w_005_808);
  and2 I006_324(w_006_324, w_001_1262, w_004_084);
  not1 I006_325(w_006_325, w_001_513);
  and2 I006_326(w_006_326, w_001_300, w_001_1246);
  and2 I006_327(w_006_327, w_002_209, w_000_928);
  not1 I006_328(w_006_328, w_000_1023);
  or2  I006_329(w_006_329, w_003_086, w_001_1083);
  nand2 I006_330(w_006_330, w_004_186, w_001_1222);
  not1 I006_331(w_006_331, w_002_485);
  or2  I006_332(w_006_332, w_001_243, w_000_300);
  nand2 I006_333(w_006_333, w_005_642, w_000_1035);
  nand2 I006_334(w_006_334, w_003_144, w_001_1405);
  nand2 I006_335(w_006_335, w_005_428, w_002_173);
  nand2 I006_336(w_006_336, w_004_444, w_000_850);
  not1 I006_337(w_006_337, w_001_425);
  or2  I006_338(w_006_338, w_002_074, w_002_133);
  or2  I006_339(w_006_339, w_002_433, w_001_081);
  nand2 I006_340(w_006_340, w_005_1158, w_004_860);
  not1 I006_341(w_006_341, w_004_617);
  or2  I006_342(w_006_342, w_003_118, w_004_142);
  or2  I006_343(w_006_343, w_000_586, w_001_656);
  nand2 I007_000(w_007_000, w_004_234, w_003_055);
  and2 I007_001(w_007_001, w_001_553, w_002_183);
  not1 I007_002(w_007_002, w_002_422);
  or2  I007_003(w_007_003, w_002_111, w_002_521);
  or2  I007_005(w_007_005, w_001_218, w_001_589);
  nand2 I007_009(w_007_009, w_002_573, w_004_1166);
  and2 I007_013(w_007_013, w_000_1805, w_006_099);
  or2  I007_014(w_007_014, w_006_124, w_001_1027);
  or2  I007_015(w_007_015, w_001_300, w_003_084);
  not1 I007_017(w_007_017, w_005_627);
  or2  I007_018(w_007_018, w_004_1719, w_006_343);
  not1 I007_019(w_007_019, w_006_261);
  not1 I007_020(w_007_020, w_005_111);
  and2 I007_021(w_007_021, w_001_1040, w_002_430);
  not1 I007_022(w_007_022, w_001_014);
  not1 I007_023(w_007_023, w_003_061);
  not1 I007_024(w_007_024, w_004_935);
  or2  I007_025(w_007_025, w_001_104, w_002_416);
  nand2 I007_026(w_007_026, w_001_750, w_000_558);
  or2  I007_027(w_007_027, w_000_1671, w_002_185);
  not1 I007_028(w_007_028, w_006_255);
  not1 I007_030(w_007_030, w_004_1085);
  nand2 I007_031(w_007_031, w_004_724, w_004_743);
  or2  I007_032(w_007_032, w_003_239, w_005_318);
  not1 I007_033(w_007_033, w_006_055);
  or2  I007_034(w_007_034, w_000_180, w_001_1171);
  not1 I007_035(w_007_035, w_005_1493);
  nand2 I007_036(w_007_036, w_006_285, w_005_1404);
  and2 I007_037(w_007_037, w_002_066, w_005_1441);
  not1 I007_038(w_007_038, w_002_165);
  nand2 I007_039(w_007_039, w_001_738, w_006_233);
  and2 I007_042(w_007_042, w_000_474, w_005_760);
  not1 I007_043(w_007_043, w_002_209);
  not1 I007_044(w_007_044, w_006_094);
  not1 I007_045(w_007_045, w_005_1257);
  nand2 I007_046(w_007_046, w_006_237, w_000_1691);
  and2 I007_048(w_007_048, w_001_444, w_005_094);
  and2 I007_049(w_007_049, w_002_350, w_003_259);
  nand2 I007_051(w_007_051, w_002_411, w_005_1658);
  not1 I007_053(w_007_053, w_001_622);
  not1 I007_054(w_007_054, w_005_1175);
  not1 I007_055(w_007_055, w_006_243);
  nand2 I007_057(w_007_057, w_004_1484, w_003_227);
  and2 I007_058(w_007_058, w_005_651, w_001_1263);
  and2 I007_059(w_007_059, w_002_095, w_003_246);
  or2  I007_060(w_007_060, w_000_1240, w_006_164);
  not1 I007_061(w_007_061, w_002_473);
  or2  I007_062(w_007_062, w_001_686, w_006_340);
  not1 I007_063(w_007_063, w_005_112);
  not1 I007_064(w_007_064, w_001_1597);
  not1 I007_066(w_007_066, w_003_125);
  nand2 I007_068(w_007_068, w_006_118, w_004_1278);
  not1 I007_069(w_007_069, w_001_1687);
  not1 I007_071(w_007_071, w_003_181);
  and2 I007_072(w_007_072, w_005_490, w_005_1349);
  and2 I007_074(w_007_074, w_001_929, w_000_831);
  not1 I007_077(w_007_077, w_000_1447);
  nand2 I007_079(w_007_079, w_005_1579, w_004_854);
  not1 I007_080(w_007_080, w_003_257);
  not1 I007_081(w_007_081, w_004_147);
  or2  I007_082(w_007_082, w_003_304, w_005_232);
  or2  I007_084(w_007_084, w_005_1186, w_004_315);
  nand2 I007_085(w_007_085, w_006_224, w_001_346);
  not1 I007_088(w_007_088, w_006_083);
  nand2 I007_090(w_007_090, w_000_1350, w_004_765);
  nand2 I007_091(w_007_091, w_001_261, w_000_861);
  not1 I007_092(w_007_092, w_004_469);
  and2 I007_095(w_007_095, w_002_110, w_006_224);
  not1 I007_097(w_007_097, w_003_211);
  and2 I007_098(w_007_098, w_003_105, w_006_238);
  not1 I007_101(w_007_101, w_006_327);
  nand2 I007_102(w_007_102, w_006_247, w_002_564);
  not1 I007_103(w_007_103, w_006_116);
  not1 I007_104(w_007_104, w_000_563);
  and2 I007_105(w_007_105, w_005_840, w_001_1303);
  and2 I007_106(w_007_106, w_003_037, w_002_112);
  nand2 I007_107(w_007_107, w_000_551, w_004_1828);
  not1 I007_108(w_007_108, w_001_999);
  and2 I007_109(w_007_109, w_006_030, w_006_200);
  and2 I007_110(w_007_110, w_005_1094, w_000_525);
  and2 I007_111(w_007_111, w_005_1440, w_000_1005);
  or2  I007_113(w_007_113, w_006_111, w_000_205);
  not1 I007_114(w_007_114, w_002_386);
  or2  I007_115(w_007_115, w_004_1737, w_000_1031);
  nand2 I007_118(w_007_118, w_002_346, w_000_640);
  not1 I007_119(w_007_119, w_002_112);
  not1 I007_120(w_007_120, w_006_326);
  or2  I007_121(w_007_121, w_004_1235, w_005_169);
  and2 I007_124(w_007_124, w_001_035, w_002_022);
  and2 I007_125(w_007_125, w_002_203, w_005_1223);
  or2  I007_126(w_007_126, w_002_201, w_001_1249);
  and2 I007_127(w_007_127, w_005_244, w_005_1651);
  not1 I007_128(w_007_128, w_001_131);
  nand2 I007_130(w_007_130, w_004_1454, w_004_885);
  or2  I007_131(w_007_131, w_004_447, w_004_1390);
  or2  I007_132(w_007_132, w_002_019, w_006_066);
  nand2 I007_135(w_007_135, w_006_068, w_004_975);
  or2  I007_136(w_007_136, w_004_659, w_006_140);
  not1 I007_137(w_007_137, w_003_066);
  or2  I007_138(w_007_138, w_004_1508, w_006_215);
  or2  I007_141(w_007_141, w_006_019, w_003_172);
  and2 I007_144(w_007_144, w_003_007, w_002_071);
  or2  I007_146(w_007_146, w_003_183, w_005_1234);
  or2  I007_147(w_007_147, w_000_1539, w_004_1362);
  not1 I007_148(w_007_148, w_000_174);
  and2 I007_149(w_007_149, w_001_783, w_003_267);
  nand2 I007_151(w_007_151, w_004_1239, w_000_1411);
  not1 I007_152(w_007_152, w_005_1310);
  not1 I007_154(w_007_154, w_004_137);
  or2  I007_155(w_007_155, w_003_167, w_001_862);
  nand2 I007_157(w_007_157, w_002_033, w_000_651);
  not1 I007_158(w_007_158, w_005_242);
  not1 I007_159(w_007_159, w_004_953);
  and2 I007_162(w_007_162, w_001_487, w_002_030);
  nand2 I007_164(w_007_164, w_003_027, w_000_966);
  nand2 I007_166(w_007_166, w_002_400, w_002_224);
  not1 I007_168(w_007_168, w_005_368);
  or2  I007_170(w_007_170, w_002_589, w_002_528);
  and2 I007_171(w_007_171, w_005_1422, w_000_1843);
  not1 I007_174(w_007_174, w_001_1331);
  and2 I007_175(w_007_175, w_006_027, w_005_1646);
  not1 I007_176(w_007_176, w_004_1232);
  or2  I007_181(w_007_181, w_000_1385, w_006_320);
  or2  I007_182(w_007_182, w_003_052, w_002_583);
  not1 I007_183(w_007_183, w_004_167);
  or2  I007_186(w_007_186, w_004_324, w_004_973);
  not1 I007_187(w_007_187, w_003_260);
  nand2 I007_188(w_007_188, w_002_131, w_005_293);
  not1 I007_189(w_007_189, w_003_274);
  nand2 I007_190(w_007_190, w_005_844, w_005_593);
  nand2 I007_193(w_007_193, w_000_785, w_006_114);
  and2 I007_194(w_007_194, w_002_226, w_001_1670);
  not1 I007_199(w_007_199, w_002_212);
  or2  I007_200(w_007_200, w_006_261, w_000_331);
  or2  I007_202(w_007_202, w_005_083, w_000_1410);
  or2  I007_203(w_007_203, w_001_1617, w_000_333);
  nand2 I007_205(w_007_205, w_000_596, w_000_891);
  or2  I007_206(w_007_206, w_002_108, w_004_1399);
  nand2 I007_207(w_007_207, w_001_348, w_003_063);
  not1 I007_208(w_007_208, w_005_538);
  nand2 I007_209(w_007_209, w_003_013, w_006_030);
  not1 I007_210(w_007_210, w_005_1023);
  or2  I007_211(w_007_211, w_005_1233, w_003_026);
  and2 I007_212(w_007_212, w_003_222, w_005_378);
  nand2 I007_213(w_007_213, w_005_1080, w_002_323);
  nand2 I007_214(w_007_214, w_001_1617, w_002_183);
  nand2 I007_215(w_007_215, w_000_1074, w_006_268);
  nand2 I007_216(w_007_216, w_003_066, w_003_120);
  or2  I007_218(w_007_218, w_000_075, w_001_018);
  and2 I007_221(w_007_221, w_001_1369, w_003_083);
  not1 I007_222(w_007_222, w_006_245);
  and2 I007_223(w_007_223, w_002_059, w_006_222);
  and2 I007_224(w_007_224, w_000_1499, w_006_260);
  nand2 I007_225(w_007_225, w_005_294, w_001_575);
  and2 I007_228(w_007_228, w_004_550, w_003_207);
  nand2 I007_229(w_007_229, w_000_843, w_000_1505);
  or2  I007_230(w_007_230, w_002_146, w_000_1837);
  nand2 I007_232(w_007_232, w_004_301, w_004_530);
  or2  I007_233(w_007_233, w_004_1337, w_002_475);
  nand2 I007_235(w_007_235, w_005_894, w_004_814);
  or2  I007_236(w_007_236, w_002_077, w_004_476);
  or2  I007_237(w_007_237, w_002_071, w_004_1684);
  nand2 I007_238(w_007_238, w_000_1844, w_003_082);
  nand2 I007_241(w_007_241, w_005_999, w_006_165);
  and2 I007_243(w_007_243, w_004_750, w_006_105);
  not1 I007_244(w_007_244, w_006_316);
  not1 I007_245(w_007_245, w_000_694);
  nand2 I007_247(w_007_247, w_005_707, w_000_1046);
  and2 I007_251(w_007_251, w_000_033, w_005_019);
  nand2 I007_252(w_007_252, w_006_052, w_003_256);
  not1 I007_253(w_007_253, w_004_1832);
  not1 I007_255(w_007_255, w_003_083);
  or2  I007_257(w_007_257, w_003_094, w_002_094);
  nand2 I007_258(w_007_258, w_004_004, w_000_1845);
  or2  I007_261(w_007_261, w_002_064, w_002_507);
  not1 I007_264(w_007_264, w_000_1387);
  nand2 I007_266(w_007_266, w_006_009, w_001_1117);
  nand2 I007_267(w_007_267, w_006_207, w_000_142);
  and2 I007_268(w_007_268, w_000_800, w_001_644);
  not1 I007_269(w_007_269, w_002_038);
  and2 I007_270(w_007_270, w_004_213, w_004_488);
  and2 I007_271(w_007_271, w_002_227, w_001_1398);
  or2  I007_272(w_007_272, w_006_086, w_003_289);
  not1 I007_275(w_007_275, w_005_1501);
  and2 I007_277(w_007_277, w_005_748, w_004_1827);
  and2 I007_278(w_007_278, w_006_054, w_004_342);
  nand2 I007_279(w_007_279, w_001_148, w_000_1260);
  nand2 I007_280(w_007_280, w_002_425, w_001_1500);
  not1 I007_283(w_007_283, w_004_227);
  nand2 I007_285(w_007_285, w_003_141, w_002_235);
  and2 I007_288(w_007_288, w_005_1223, w_006_192);
  nand2 I007_289(w_007_289, w_002_319, w_002_369);
  not1 I007_290(w_007_290, w_002_391);
  and2 I007_292(w_007_292, w_005_970, w_004_554);
  nand2 I007_293(w_007_293, w_005_477, w_004_1191);
  nand2 I007_294(w_007_294, w_006_325, w_001_816);
  or2  I007_295(w_007_295, w_005_728, w_000_1104);
  and2 I007_298(w_007_298, w_001_1515, w_003_114);
  or2  I007_299(w_007_299, w_006_070, w_005_275);
  or2  I007_304(w_007_304, w_005_640, w_000_1356);
  nand2 I007_305(w_007_305, w_000_1354, w_006_000);
  and2 I007_306(w_007_306, w_003_110, w_004_904);
  and2 I007_307(w_007_307, w_000_1232, w_005_1298);
  and2 I007_309(w_007_309, w_004_486, w_004_458);
  or2  I007_311(w_007_311, w_001_856, w_004_1797);
  and2 I007_313(w_007_313, w_002_387, w_006_064);
  nand2 I007_314(w_007_314, w_005_205, w_000_1846);
  not1 I007_315(w_007_315, w_001_1661);
  or2  I007_316(w_007_316, w_003_120, w_006_105);
  and2 I007_317(w_007_317, w_001_548, w_002_164);
  and2 I007_318(w_007_318, w_005_286, w_000_429);
  nand2 I007_320(w_007_320, w_001_921, w_005_672);
  or2  I007_322(w_007_322, w_005_995, w_002_466);
  or2  I007_325(w_007_325, w_001_273, w_003_031);
  or2  I007_327(w_007_327, w_000_144, w_006_002);
  or2  I007_329(w_007_329, w_006_032, w_006_119);
  and2 I007_330(w_007_330, w_001_100, w_000_1408);
  nand2 I007_337(w_007_337, w_002_040, w_003_315);
  not1 I007_338(w_007_338, w_004_1210);
  or2  I007_340(w_007_340, w_005_785, w_005_139);
  or2  I007_342(w_007_342, w_001_1256, w_000_686);
  or2  I007_346(w_007_346, w_000_782, w_004_1033);
  and2 I007_348(w_007_348, w_000_734, w_003_286);
  and2 I007_349(w_007_349, w_000_1630, w_002_290);
  or2  I007_351(w_007_351, w_000_339, w_001_966);
  and2 I007_353(w_007_353, w_005_709, w_005_015);
  or2  I007_354(w_007_354, w_000_693, w_003_129);
  and2 I007_357(w_007_357, w_004_1468, w_000_1847);
  nand2 I007_358(w_007_358, w_000_017, w_003_189);
  or2  I007_359(w_007_359, w_006_005, w_000_1265);
  and2 I007_360(w_007_360, w_005_965, w_004_905);
  not1 I007_364(w_007_364, w_000_1645);
  and2 I007_366(w_007_366, w_003_232, w_000_1428);
  and2 I007_367(w_007_367, w_003_074, w_004_824);
  and2 I007_368(w_007_368, w_002_238, w_003_049);
  or2  I007_370(w_007_370, w_000_278, w_003_176);
  not1 I007_373(w_007_373, w_003_092);
  not1 I007_377(w_007_377, w_002_239);
  or2  I007_378(w_007_378, w_001_1109, w_002_516);
  and2 I007_379(w_007_379, w_001_702, w_000_586);
  not1 I007_380(w_007_380, w_004_088);
  nand2 I007_381(w_007_381, w_003_064, w_002_127);
  and2 I007_382(w_007_382, w_001_055, w_003_173);
  nand2 I007_384(w_007_384, w_006_160, w_001_1675);
  not1 I007_388(w_007_388, w_001_1464);
  not1 I007_391(w_007_391, w_005_774);
  nand2 I007_393(w_007_393, w_002_291, w_004_929);
  or2  I007_398(w_007_398, w_005_1140, w_006_312);
  not1 I007_399(w_007_399, w_003_048);
  not1 I007_401(w_007_401, w_001_1034);
  nand2 I007_402(w_007_402, w_003_189, w_006_085);
  and2 I007_405(w_007_405, w_000_961, w_000_171);
  nand2 I007_406(w_007_406, w_001_571, w_006_198);
  not1 I007_411(w_007_411, w_002_016);
  not1 I007_415(w_007_415, w_003_091);
  nand2 I007_417(w_007_417, w_005_1652, w_005_274);
  or2  I007_418(w_007_418, w_002_109, w_001_357);
  nand2 I007_421(w_007_421, w_003_238, w_003_262);
  and2 I007_423(w_007_423, w_005_376, w_000_166);
  nand2 I007_434(w_007_434, w_005_236, w_002_540);
  nand2 I007_436(w_007_436, w_001_895, w_003_068);
  or2  I007_438(w_007_438, w_002_078, w_000_1051);
  and2 I007_439(w_007_439, w_002_239, w_004_1674);
  and2 I007_441(w_007_441, w_001_833, w_002_530);
  or2  I007_442(w_007_442, w_000_1343, w_006_116);
  nand2 I007_443(w_007_443, w_002_082, w_006_235);
  nand2 I007_444(w_007_444, w_006_231, w_003_065);
  and2 I007_446(w_007_446, w_005_1622, w_006_193);
  nand2 I007_447(w_007_447, w_003_066, w_003_119);
  and2 I007_449(w_007_449, w_001_077, w_005_997);
  and2 I007_451(w_007_451, w_003_268, w_003_170);
  or2  I007_453(w_007_453, w_002_456, w_004_1741);
  or2  I007_458(w_007_458, w_003_207, w_002_100);
  nand2 I007_463(w_007_463, w_005_611, w_003_241);
  and2 I007_466(w_007_466, w_003_318, w_001_1039);
  nand2 I007_475(w_007_475, w_002_101, w_002_177);
  nand2 I007_477(w_007_477, w_002_057, w_002_478);
  and2 I007_478(w_007_478, w_004_595, w_004_852);
  nand2 I007_479(w_007_479, w_001_228, w_003_172);
  or2  I007_482(w_007_482, w_006_227, w_000_1286);
  and2 I007_483(w_007_483, w_001_170, w_003_247);
  and2 I007_484(w_007_484, w_005_1092, w_004_602);
  and2 I007_485(w_007_485, w_001_1197, w_000_407);
  nand2 I007_490(w_007_490, w_005_068, w_005_139);
  and2 I007_491(w_007_491, w_000_741, w_005_857);
  or2  I007_498(w_007_498, w_004_1412, w_002_089);
  nand2 I007_503(w_007_503, w_006_264, w_000_1848);
  not1 I007_509(w_007_509, w_001_1011);
  nand2 I007_515(w_007_515, w_005_674, w_006_194);
  or2  I007_517(w_007_517, w_001_545, w_000_937);
  nand2 I007_518(w_007_518, w_002_301, w_003_251);
  nand2 I007_520(w_007_520, w_004_144, w_005_315);
  and2 I007_523(w_007_523, w_006_139, w_004_1269);
  and2 I007_524(w_007_524, w_004_558, w_001_813);
  nand2 I007_525(w_007_525, w_004_1065, w_006_137);
  and2 I007_526(w_007_526, w_004_1874, w_005_313);
  or2  I007_531(w_007_531, w_006_143, w_004_207);
  and2 I007_532(w_007_532, w_003_096, w_000_1610);
  or2  I007_534(w_007_534, w_004_606, w_001_1484);
  nand2 I007_539(w_007_539, w_004_853, w_005_839);
  nand2 I007_540(w_007_540, w_006_133, w_002_495);
  nand2 I007_543(w_007_543, w_004_1501, w_001_053);
  or2  I007_544(w_007_544, w_001_1100, w_005_485);
  not1 I007_546(w_007_546, w_004_433);
  and2 I007_547(w_007_547, w_005_199, w_003_315);
  and2 I007_549(w_007_549, w_005_444, w_004_610);
  or2  I007_550(w_007_550, w_005_663, w_003_031);
  not1 I007_555(w_007_555, w_001_824);
  nand2 I007_559(w_007_559, w_005_1569, w_004_373);
  and2 I007_561(w_007_561, w_006_025, w_000_946);
  not1 I007_563(w_007_563, w_000_1849);
  nand2 I007_564(w_007_564, w_002_253, w_003_172);
  nand2 I007_567(w_007_567, w_006_019, w_003_090);
  nand2 I007_568(w_007_568, w_002_527, w_004_404);
  nand2 I007_569(w_007_569, w_002_284, w_000_1629);
  not1 I007_573(w_007_573, w_004_114);
  nand2 I007_576(w_007_576, w_005_1588, w_000_949);
  nand2 I007_577(w_007_577, w_001_405, w_003_029);
  nand2 I007_579(w_007_579, w_000_1220, w_004_314);
  not1 I007_580(w_007_580, w_001_780);
  or2  I007_583(w_007_583, w_000_1187, w_006_303);
  not1 I007_586(w_007_586, w_003_164);
  nand2 I007_589(w_007_589, w_004_1436, w_001_274);
  or2  I007_590(w_007_590, w_006_128, w_006_097);
  or2  I007_592(w_007_592, w_005_929, w_006_215);
  or2  I007_597(w_007_597, w_003_011, w_006_143);
  nand2 I007_598(w_007_598, w_000_1106, w_002_567);
  and2 I007_599(w_007_599, w_000_1377, w_006_097);
  or2  I007_601(w_007_601, w_006_142, w_001_807);
  and2 I007_603(w_007_603, w_000_603, w_001_111);
  nand2 I007_604(w_007_604, w_001_960, w_000_1764);
  not1 I007_605(w_007_605, w_002_324);
  not1 I007_609(w_007_609, w_006_330);
  nand2 I007_610(w_007_610, w_006_245, w_002_201);
  not1 I007_612(w_007_612, w_003_070);
  or2  I007_613(w_007_613, w_003_244, w_006_010);
  and2 I007_618(w_007_618, w_002_151, w_004_605);
  not1 I007_622(w_007_622, w_004_1858);
  and2 I007_623(w_007_623, w_000_1332, w_001_602);
  and2 I007_624(w_007_624, w_002_052, w_004_116);
  or2  I007_627(w_007_627, w_000_1726, w_004_118);
  or2  I007_628(w_007_628, w_000_1176, w_006_265);
  or2  I007_632(w_007_632, w_003_000, w_000_1024);
  and2 I007_634(w_007_634, w_003_074, w_003_312);
  nand2 I007_636(w_007_636, w_003_290, w_001_561);
  or2  I007_637(w_007_637, w_001_1376, w_001_1568);
  not1 I007_638(w_007_638, w_004_1487);
  nand2 I007_639(w_007_639, w_001_479, w_005_577);
  or2  I007_640(w_007_640, w_004_1174, w_004_008);
  or2  I007_646(w_007_646, w_000_501, w_005_1561);
  not1 I007_652(w_007_652, w_002_027);
  or2  I007_654(w_007_654, w_001_1288, w_001_134);
  nand2 I007_655(w_007_655, w_000_1851, w_002_432);
  and2 I007_656(w_007_656, w_002_526, w_004_498);
  or2  I007_657(w_007_657, w_003_086, w_002_013);
  or2  I007_660(w_007_660, w_005_201, w_004_603);
  not1 I007_663(w_007_663, w_006_120);
  nand2 I007_664(w_007_664, w_000_1190, w_004_1583);
  nand2 I007_666(w_007_666, w_001_590, w_003_120);
  or2  I007_673(w_007_673, w_001_873, w_005_782);
  nand2 I007_676(w_007_676, w_000_1649, w_005_149);
  nand2 I007_680(w_007_680, w_006_268, w_006_252);
  and2 I007_682(w_007_682, w_006_046, w_004_250);
  or2  I007_687(w_007_687, w_006_128, w_002_581);
  not1 I007_689(w_007_689, w_000_398);
  and2 I007_691(w_007_691, w_000_1852, w_005_766);
  nand2 I007_697(w_007_697, w_001_409, w_006_302);
  or2  I007_698(w_007_698, w_004_796, w_001_230);
  nand2 I007_699(w_007_699, w_005_1285, w_003_074);
  not1 I007_701(w_007_701, w_002_094);
  and2 I007_703(w_007_703, w_002_030, w_006_210);
  nand2 I007_704(w_007_704, w_006_240, w_005_668);
  not1 I007_712(w_007_712, w_005_303);
  not1 I007_713(w_007_713, w_001_103);
  nand2 I007_714(w_007_714, w_005_276, w_002_270);
  nand2 I007_715(w_007_715, w_001_161, w_001_352);
  and2 I007_720(w_007_720, w_001_051, w_004_1328);
  or2  I007_722(w_007_722, w_004_1523, w_002_088);
  nand2 I007_725(w_007_725, w_002_356, w_005_541);
  not1 I007_726(w_007_726, w_006_273);
  or2  I007_729(w_007_729, w_002_191, w_006_024);
  not1 I007_732(w_007_732, w_005_286);
  or2  I007_734(w_007_734, w_005_1268, w_001_079);
  nand2 I007_738(w_007_738, w_004_298, w_003_161);
  not1 I007_740(w_007_740, w_006_165);
  not1 I007_741(w_007_741, w_003_162);
  nand2 I007_742(w_007_742, w_006_092, w_004_1358);
  not1 I007_744(w_007_744, w_005_825);
  or2  I007_746(w_007_746, w_005_1523, w_002_136);
  nand2 I007_747(w_007_747, w_003_218, w_006_222);
  and2 I007_750(w_007_750, w_000_193, w_005_208);
  not1 I007_752(w_007_752, w_001_1153);
  or2  I007_755(w_007_755, w_002_120, w_006_046);
  nand2 I007_756(w_007_756, w_002_140, w_003_110);
  not1 I007_757(w_007_757, w_001_303);
  or2  I007_761(w_007_761, w_003_187, w_006_116);
  or2  I007_763(w_007_763, w_001_836, w_002_422);
  nand2 I007_768(w_007_768, w_003_288, w_004_001);
  not1 I007_769(w_007_769, w_003_307);
  or2  I007_772(w_007_772, w_001_416, w_000_472);
  and2 I007_774(w_007_774, w_004_179, w_001_757);
  nand2 I007_778(w_007_778, w_002_565, w_002_219);
  not1 I007_779(w_007_779, w_003_176);
  not1 I007_781(w_007_781, w_004_211);
  nand2 I007_782(w_007_782, w_002_238, w_003_257);
  nand2 I007_784(w_007_784, w_004_1043, w_006_171);
  or2  I007_785(w_007_785, w_006_050, w_004_878);
  nand2 I007_786(w_007_786, w_005_170, w_004_1521);
  and2 I007_790(w_007_790, w_001_984, w_004_1481);
  or2  I007_793(w_007_793, w_003_003, w_001_066);
  not1 I007_796(w_007_796, w_000_1253);
  not1 I007_798(w_007_798, w_002_022);
  and2 I007_800(w_007_800, w_002_074, w_003_136);
  not1 I007_802(w_007_802, w_000_367);
  not1 I007_803(w_007_803, w_003_110);
  nand2 I007_804(w_007_804, w_006_128, w_002_369);
  or2  I007_805(w_007_805, w_005_127, w_004_978);
  nand2 I007_808(w_007_808, w_002_343, w_004_838);
  or2  I007_811(w_007_811, w_006_093, w_006_115);
  not1 I007_814(w_007_814, w_001_1293);
  or2  I007_816(w_007_816, w_005_1220, w_004_011);
  nand2 I007_817(w_007_817, w_005_306, w_001_707);
  and2 I007_822(w_007_822, w_001_692, w_006_052);
  or2  I007_823(w_007_823, w_002_170, w_006_305);
  or2  I007_828(w_007_828, w_005_1261, w_005_056);
  or2  I007_829(w_007_829, w_001_431, w_000_1687);
  nand2 I007_834(w_007_834, w_006_042, w_002_096);
  or2  I007_837(w_007_837, w_002_344, w_004_732);
  nand2 I007_838(w_007_838, w_002_530, w_004_1288);
  or2  I007_839(w_007_839, w_002_312, w_004_955);
  nand2 I007_840(w_007_840, w_006_015, w_001_1586);
  and2 I007_847(w_007_847, w_006_052, w_004_1210);
  not1 I007_849(w_007_849, w_002_108);
  not1 I007_850(w_007_850, w_002_171);
  not1 I007_851(w_007_851, w_004_514);
  nand2 I007_855(w_007_855, w_004_1855, w_005_798);
  or2  I007_858(w_007_858, w_002_427, w_001_1670);
  or2  I007_860(w_007_860, w_006_286, w_002_044);
  or2  I007_862(w_007_862, w_004_721, w_005_893);
  or2  I007_863(w_007_863, w_003_181, w_004_1188);
  or2  I007_865(w_007_865, w_005_986, w_006_046);
  not1 I007_869(w_007_869, w_003_006);
  nand2 I007_871(w_007_871, w_001_900, w_004_241);
  nand2 I007_873(w_007_873, w_006_078, w_002_423);
  not1 I007_874(w_007_874, w_002_570);
  nand2 I007_875(w_007_875, w_004_1631, w_006_195);
  nand2 I007_879(w_007_879, w_005_882, w_003_277);
  and2 I007_880(w_007_880, w_003_208, w_001_1113);
  nand2 I007_881(w_007_881, w_005_390, w_006_164);
  and2 I007_883(w_007_883, w_001_472, w_004_1381);
  or2  I007_884(w_007_884, w_004_443, w_004_1101);
  nand2 I007_887(w_007_887, w_004_755, w_000_1538);
  or2  I007_889(w_007_889, w_004_488, w_004_170);
  nand2 I007_891(w_007_891, w_001_1631, w_006_201);
  and2 I007_892(w_007_892, w_004_356, w_006_168);
  or2  I007_894(w_007_894, w_003_226, w_005_1307);
  and2 I007_900(w_007_900, w_005_197, w_004_1040);
  nand2 I007_903(w_007_903, w_001_013, w_004_1882);
  not1 I007_904(w_007_904, w_001_271);
  nand2 I007_905(w_007_905, w_003_111, w_003_310);
  not1 I007_907(w_007_907, w_001_016);
  nand2 I007_915(w_007_915, w_003_037, w_000_014);
  nand2 I007_916(w_007_916, w_002_328, w_003_027);
  or2  I007_920(w_007_920, w_002_529, w_000_390);
  nand2 I007_921(w_007_921, w_004_243, w_002_310);
  and2 I007_924(w_007_924, w_001_250, w_002_223);
  or2  I007_925(w_007_925, w_004_870, w_001_365);
  nand2 I007_927(w_007_927, w_003_061, w_005_1322);
  and2 I007_928(w_007_928, w_005_226, w_005_731);
  and2 I007_929(w_007_929, w_006_205, w_000_1194);
  and2 I007_931(w_007_931, w_005_117, w_006_159);
  nand2 I007_934(w_007_934, w_000_906, w_000_386);
  and2 I007_935(w_007_935, w_005_1470, w_000_272);
  or2  I007_941(w_007_941, w_002_201, w_000_778);
  or2  I007_944(w_007_944, w_002_081, w_004_1105);
  or2  I007_945(w_007_945, w_002_535, w_006_089);
  nand2 I007_946(w_007_946, w_006_328, w_000_022);
  not1 I007_947(w_007_947, w_005_505);
  nand2 I007_948(w_007_948, w_000_247, w_001_1053);
  not1 I007_951(w_007_951, w_001_234);
  and2 I007_953(w_007_953, w_003_304, w_001_1049);
  not1 I007_954(w_007_954, w_004_1907);
  not1 I007_957(w_007_957, w_001_417);
  and2 I007_961(w_007_961, w_006_265, w_002_303);
  not1 I007_963(w_007_963, w_006_201);
  or2  I007_964(w_007_964, w_002_450, w_000_773);
  nand2 I007_966(w_007_966, w_004_1757, w_006_041);
  not1 I007_967(w_007_967, w_000_1720);
  not1 I007_969(w_007_969, w_003_224);
  nand2 I007_975(w_007_975, w_001_1373, w_004_687);
  or2  I007_977(w_007_977, w_001_1638, w_006_233);
  not1 I007_979(w_007_979, w_005_506);
  and2 I007_980(w_007_980, w_001_864, w_002_039);
  not1 I007_981(w_007_981, w_006_188);
  or2  I007_987(w_007_987, w_006_150, w_001_1030);
  or2  I007_996(w_007_996, w_001_1408, w_000_837);
  or2  I007_997(w_007_997, w_005_1580, w_001_659);
  and2 I007_999(w_007_999, w_002_075, w_001_1358);
  nand2 I007_1002(w_007_1002, w_004_288, w_004_1692);
  not1 I007_1003(w_007_1003, w_003_172);
  or2  I007_1010(w_007_1010, w_002_092, w_003_078);
  and2 I007_1020(w_007_1020, w_001_1547, w_005_048);
  nand2 I007_1022(w_007_1022, w_003_116, w_004_422);
  not1 I007_1026(w_007_1026, w_006_126);
  or2  I007_1033(w_007_1033, w_005_321, w_001_461);
  nand2 I007_1036(w_007_1036, w_003_182, w_005_790);
  nand2 I007_1042(w_007_1042, w_003_189, w_002_333);
  and2 I007_1043(w_007_1043, w_000_069, w_005_216);
  nand2 I007_1044(w_007_1044, w_000_817, w_000_1571);
  and2 I007_1045(w_007_1045, w_003_112, w_000_018);
  or2  I007_1046(w_007_1046, w_001_1495, w_000_055);
  not1 I007_1047(w_007_1047, w_002_214);
  and2 I007_1048(w_007_1048, w_005_065, w_002_562);
  or2  I007_1049(w_007_1049, w_004_1029, w_000_229);
  and2 I007_1054(w_007_1054, w_000_1859, w_000_082);
  or2  I007_1060(w_007_1060, w_000_1651, w_004_084);
  and2 I007_1061(w_007_1061, w_002_080, w_001_835);
  nand2 I007_1063(w_007_1063, w_005_472, w_004_312);
  or2  I007_1065(w_007_1065, w_001_810, w_006_341);
  or2  I007_1068(w_007_1068, w_001_272, w_002_177);
  or2  I007_1069(w_007_1069, w_006_170, w_002_259);
  or2  I007_1077(w_007_1077, w_002_087, w_002_063);
  and2 I007_1078(w_007_1078, w_005_366, w_003_135);
  nand2 I007_1080(w_007_1080, w_006_184, w_002_305);
  or2  I007_1083(w_007_1083, w_003_262, w_005_731);
  or2  I007_1084(w_007_1084, w_000_1862, w_003_304);
  or2  I007_1085(w_007_1085, w_006_343, w_004_1030);
  nand2 I007_1086(w_007_1086, w_004_1361, w_003_180);
  not1 I007_1087(w_007_1087, w_006_250);
  not1 I007_1089(w_007_1089, w_002_478);
  nand2 I007_1090(w_007_1090, w_005_280, w_003_132);
  and2 I007_1094(w_007_1094, w_006_219, w_000_1101);
  nand2 I007_1095(w_007_1095, w_001_480, w_002_230);
  not1 I007_1097(w_007_1097, w_006_321);
  and2 I007_1101(w_007_1101, w_006_187, w_000_1685);
  nand2 I007_1103(w_007_1103, w_004_665, w_001_836);
  and2 I007_1104(w_007_1104, w_003_058, w_006_112);
  not1 I007_1110(w_007_1110, w_002_307);
  or2  I007_1117(w_007_1117, w_000_1488, w_002_410);
  nand2 I007_1118(w_007_1118, w_005_190, w_006_068);
  or2  I007_1119(w_007_1119, w_004_1748, w_006_123);
  nand2 I007_1120(w_007_1120, w_005_823, w_001_169);
  not1 I007_1123(w_007_1123, w_006_116);
  or2  I007_1127(w_007_1127, w_003_052, w_006_240);
  and2 I007_1129(w_007_1129, w_006_262, w_000_369);
  or2  I007_1130(w_007_1130, w_004_837, w_000_1195);
  not1 I007_1132(w_007_1132, w_005_276);
  and2 I007_1134(w_007_1134, w_003_025, w_005_1493);
  nand2 I007_1137(w_007_1137, w_000_563, w_006_326);
  nand2 I007_1138(w_007_1138, w_000_707, w_000_536);
  not1 I007_1140(w_007_1140, w_006_253);
  and2 I007_1141(w_007_1141, w_000_689, w_006_116);
  not1 I007_1142(w_007_1142, w_000_1865);
  or2  I007_1148(w_007_1148, w_006_259, w_003_137);
  not1 I007_1151(w_007_1151, w_005_1636);
  not1 I007_1153(w_007_1153, w_004_046);
  and2 I007_1157(w_007_1157, w_000_670, w_006_076);
  or2  I007_1159(w_007_1159, w_003_010, w_003_008);
  and2 I007_1160(w_007_1160, w_000_764, w_005_1550);
  nand2 I007_1161(w_007_1161, w_000_1866, w_001_250);
  and2 I007_1168(w_007_1168, w_003_002, w_001_1242);
  not1 I007_1173(w_007_1173, w_005_1151);
  nand2 I007_1175(w_007_1175, w_006_257, w_002_260);
  and2 I007_1176(w_007_1176, w_000_931, w_005_105);
  not1 I007_1178(w_007_1178, w_006_059);
  not1 I007_1179(w_007_1179, w_001_180);
  not1 I007_1182(w_007_1182, w_005_1576);
  and2 I007_1184(w_007_1184, w_004_111, w_000_419);
  and2 I007_1187(w_007_1187, w_000_701, w_001_276);
  not1 I007_1189(w_007_1189, w_001_1228);
  nand2 I007_1190(w_007_1190, w_006_005, w_004_1615);
  not1 I007_1194(w_007_1194, w_004_1234);
  or2  I007_1197(w_007_1197, w_000_319, w_001_019);
  and2 I007_1198(w_007_1198, w_002_556, w_003_066);
  nand2 I007_1204(w_007_1204, w_002_046, w_002_272);
  not1 I007_1206(w_007_1206, w_004_1709);
  not1 I007_1208(w_007_1208, w_004_917);
  nand2 I007_1209(w_007_1209, w_006_177, w_001_107);
  nand2 I007_1211(w_007_1211, w_002_244, w_001_090);
  nand2 I007_1214(w_007_1214, w_004_841, w_004_013);
  nand2 I007_1215(w_007_1215, w_006_130, w_002_299);
  nand2 I007_1219(w_007_1219, w_006_196, w_001_890);
  not1 I007_1223(w_007_1223, w_004_1413);
  not1 I007_1227(w_007_1227, w_000_1395);
  and2 I007_1229(w_007_1229, w_001_1393, w_003_177);
  nand2 I007_1230(w_007_1230, w_005_1591, w_002_211);
  or2  I007_1231(w_007_1231, w_001_1146, w_003_137);
  or2  I007_1233(w_007_1233, w_002_084, w_001_859);
  not1 I007_1234(w_007_1234, w_001_254);
  not1 I007_1235(w_007_1235, w_001_160);
  or2  I007_1243(w_007_1243, w_001_1479, w_006_192);
  or2  I007_1244(w_007_1244, w_004_236, w_004_583);
  not1 I007_1245(w_007_1245, w_006_027);
  not1 I007_1246(w_007_1246, w_002_128);
  nand2 I007_1247(w_007_1247, w_006_322, w_005_1534);
  not1 I007_1248(w_007_1248, w_005_075);
  nand2 I007_1250(w_007_1250, w_000_820, w_003_185);
  and2 I007_1251(w_007_1251, w_002_132, w_000_1261);
  or2  I007_1256(w_007_1256, w_004_653, w_006_056);
  or2  I007_1257(w_007_1257, w_000_953, w_005_619);
  and2 I007_1258(w_007_1258, w_003_280, w_002_150);
  and2 I007_1259(w_007_1259, w_006_007, w_002_144);
  nand2 I007_1261(w_007_1261, w_006_103, w_002_410);
  or2  I007_1263(w_007_1263, w_006_038, w_005_922);
  and2 I007_1264(w_007_1264, w_004_1893, w_004_293);
  and2 I007_1269(w_007_1269, w_005_1082, w_006_311);
  or2  I007_1276(w_007_1276, w_001_066, w_003_053);
  nand2 I007_1279(w_007_1279, w_002_558, w_005_699);
  or2  I007_1281(w_007_1281, w_005_1061, w_002_457);
  and2 I007_1284(w_007_1284, w_002_476, w_004_1653);
  not1 I007_1292(w_007_1292, w_001_939);
  not1 I007_1294(w_007_1294, w_000_1406);
  not1 I007_1295(w_007_1295, w_004_002);
  nand2 I007_1298(w_007_1298, w_006_178, w_003_001);
  and2 I007_1299(w_007_1299, w_003_311, w_006_018);
  and2 I007_1302(w_007_1302, w_001_123, w_002_434);
  or2  I007_1303(w_007_1303, w_003_162, w_001_1131);
  nand2 I007_1304(w_007_1304, w_000_268, w_002_172);
  and2 I007_1307(w_007_1307, w_002_562, w_001_869);
  and2 I007_1310(w_007_1310, w_002_438, w_003_241);
  or2  I007_1313(w_007_1313, w_004_1517, w_004_1492);
  nand2 I007_1315(w_007_1315, w_002_589, w_002_587);
  not1 I007_1316(w_007_1316, w_006_100);
  not1 I007_1318(w_007_1318, w_006_309);
  or2  I007_1321(w_007_1321, w_005_863, w_000_1340);
  and2 I007_1323(w_007_1323, w_003_245, w_006_299);
  not1 I007_1326(w_007_1326, w_000_1868);
  or2  I007_1328(w_007_1328, w_005_645, w_005_511);
  or2  I007_1331(w_007_1331, w_005_712, w_005_030);
  nand2 I007_1333(w_007_1333, w_003_036, w_003_153);
  and2 I007_1334(w_007_1334, w_003_211, w_003_164);
  not1 I007_1337(w_007_1337, w_005_1033);
  not1 I007_1338(w_007_1338, w_003_135);
  and2 I007_1340(w_007_1340, w_002_356, w_001_806);
  and2 I007_1341(w_007_1341, w_005_014, w_004_1840);
  and2 I007_1343(w_007_1343, w_006_195, w_006_242);
  nand2 I007_1345(w_007_1345, w_006_332, w_002_090);
  nand2 I007_1347(w_007_1347, w_001_796, w_000_1399);
  or2  I007_1349(w_007_1349, w_001_290, w_004_1248);
  or2  I007_1350(w_007_1350, w_006_270, w_002_395);
  and2 I007_1351(w_007_1351, w_004_813, w_003_215);
  nand2 I007_1353(w_007_1353, w_004_062, w_003_249);
  and2 I007_1355(w_007_1355, w_000_1726, w_006_124);
  or2  I007_1358(w_007_1358, w_002_145, w_001_161);
  or2  I007_1360(w_007_1360, w_001_313, w_002_354);
  and2 I007_1365(w_007_1365, w_003_139, w_000_1430);
  and2 I007_1366(w_007_1366, w_004_025, w_004_144);
  or2  I007_1368(w_007_1368, w_000_732, w_000_463);
  or2  I007_1374(w_007_1374, w_004_005, w_004_1563);
  and2 I007_1377(w_007_1377, w_004_011, w_001_073);
  nand2 I007_1378(w_007_1378, w_000_927, w_006_301);
  and2 I007_1379(w_007_1379, w_003_264, w_005_204);
  or2  I007_1384(w_007_1384, w_001_1265, w_003_312);
  not1 I007_1388(w_007_1388, w_002_398);
  or2  I007_1390(w_007_1390, w_003_113, w_002_186);
  or2  I007_1393(w_007_1393, w_004_1393, w_005_303);
  nand2 I007_1397(w_007_1397, w_002_332, w_000_006);
  nand2 I007_1402(w_007_1402, w_002_505, w_000_1131);
  not1 I007_1405(w_007_1405, w_004_1575);
  or2  I007_1406(w_007_1406, w_005_280, w_001_169);
  and2 I007_1407(w_007_1407, w_003_233, w_002_541);
  or2  I007_1412(w_007_1412, w_004_1894, w_001_274);
  nand2 I007_1415(w_007_1415, w_005_453, w_006_144);
  not1 I007_1420(w_007_1420, w_002_220);
  and2 I007_1423(w_007_1423, w_004_1083, w_002_249);
  or2  I007_1435(w_007_1435, w_000_1536, w_001_1199);
  not1 I007_1436(w_007_1436, w_004_301);
  not1 I007_1442(w_007_1442, w_002_235);
  and2 I007_1443(w_007_1443, w_003_313, w_006_087);
  or2  I007_1444(w_007_1444, w_005_1613, w_002_448);
  and2 I007_1446(w_007_1446, w_002_532, w_003_261);
  and2 I007_1449(w_007_1449, w_004_196, w_004_749);
  or2  I007_1450(w_007_1450, w_003_276, w_003_224);
  not1 I007_1451(w_007_1451, w_003_212);
  nand2 I007_1454(w_007_1454, w_000_1380, w_002_100);
  not1 I007_1455(w_007_1455, w_004_1843);
  nand2 I007_1456(w_007_1456, w_000_391, w_002_591);
  or2  I007_1458(w_007_1458, w_006_308, w_004_1692);
  nand2 I007_1459(w_007_1459, w_002_225, w_002_217);
  not1 I007_1460(w_007_1460, w_001_857);
  and2 I007_1462(w_007_1462, w_003_130, w_003_094);
  and2 I007_1465(w_007_1465, w_002_588, w_004_472);
  nand2 I007_1467(w_007_1467, w_001_087, w_000_235);
  not1 I007_1468(w_007_1468, w_005_1480);
  and2 I007_1469(w_007_1469, w_006_214, w_001_1386);
  and2 I007_1470(w_007_1470, w_002_382, w_002_161);
  not1 I007_1472(w_007_1472, w_001_615);
  not1 I007_1473(w_007_1473, w_003_283);
  or2  I007_1474(w_007_1474, w_001_1012, w_004_064);
  not1 I007_1477(w_007_1477, w_002_207);
  and2 I007_1478(w_007_1478, w_005_1542, w_006_277);
  or2  I007_1479(w_007_1479, w_006_188, w_000_1488);
  not1 I007_1480(w_007_1480, w_002_457);
  and2 I007_1481(w_007_1481, w_001_063, w_001_1566);
  not1 I007_1482(w_007_1482, w_001_033);
  nand2 I007_1484(w_007_1484, w_003_191, w_001_549);
  or2  I007_1486(w_007_1486, w_000_034, w_006_031);
  and2 I007_1487(w_007_1487, w_001_1082, w_005_128);
  not1 I007_1488(w_007_1488, w_006_337);
  nand2 I007_1492(w_007_1492, w_006_219, w_004_618);
  not1 I007_1493(w_007_1493, w_002_371);
  or2  I007_1494(w_007_1494, w_003_299, w_003_084);
  not1 I007_1495(w_007_1495, w_006_204);
  and2 I007_1497(w_007_1497, w_004_1647, w_003_183);
  or2  I007_1500(w_007_1500, w_000_207, w_000_1871);
  and2 I007_1502(w_007_1502, w_001_901, w_006_144);
  not1 I007_1504(w_007_1504, w_004_482);
  nand2 I007_1506(w_007_1506, w_004_1860, w_002_003);
  or2  I007_1507(w_007_1507, w_005_880, w_005_047);
  or2  I007_1508(w_007_1508, w_000_621, w_003_002);
  and2 I007_1510(w_007_1510, w_004_1289, w_002_491);
  and2 I007_1511(w_007_1511, w_004_973, w_005_674);
  nand2 I007_1512(w_007_1512, w_001_091, w_003_100);
  and2 I007_1513(w_007_1513, w_005_1078, w_002_430);
  and2 I007_1515(w_007_1515, w_003_190, w_004_1624);
  nand2 I007_1519(w_007_1519, w_000_236, w_001_067);
  not1 I007_1520(w_007_1520, w_002_540);
  nand2 I007_1522(w_007_1522, w_006_144, w_005_707);
  not1 I007_1524(w_007_1524, w_002_111);
  and2 I007_1527(w_007_1527, w_001_1337, w_005_853);
  and2 I007_1530(w_007_1530, w_006_039, w_006_206);
  or2  I007_1531(w_007_1531, w_006_317, w_003_088);
  not1 I007_1533(w_007_1533, w_005_444);
  and2 I007_1536(w_007_1536, w_001_691, w_002_287);
  not1 I007_1538(w_007_1538, w_005_444);
  nand2 I007_1543(w_007_1543, w_004_1354, w_003_042);
  and2 I007_1551(w_007_1551, w_000_1504, w_006_313);
  and2 I007_1554(w_007_1554, w_001_438, w_001_603);
  not1 I007_1555(w_007_1555, w_000_841);
  not1 I007_1562(w_007_1562, w_002_220);
  nand2 I007_1565(w_007_1565, w_004_1298, w_006_210);
  nand2 I007_1566(w_007_1566, w_002_198, w_005_075);
  or2  I007_1567(w_007_1567, w_002_592, w_006_020);
  or2  I007_1570(w_007_1570, w_003_150, w_002_196);
  nand2 I007_1574(w_007_1574, w_001_416, w_000_105);
  not1 I007_1579(w_007_1579, w_005_789);
  nand2 I007_1583(w_007_1583, w_006_111, w_004_973);
  and2 I007_1584(w_007_1584, w_003_143, w_006_278);
  nand2 I007_1588(w_007_1588, w_002_121, w_002_251);
  nand2 I007_1590(w_007_1590, w_006_044, w_005_1268);
  and2 I007_1592(w_007_1592, w_000_1359, w_006_040);
  or2  I007_1593(w_007_1593, w_005_1293, w_004_1626);
  nand2 I007_1594(w_007_1594, w_001_398, w_004_1546);
  nand2 I007_1595(w_007_1595, w_006_047, w_004_916);
  or2  I007_1596(w_007_1596, w_004_1743, w_004_656);
  nand2 I007_1597(w_007_1597, w_003_005, w_004_894);
  nand2 I007_1598(w_007_1598, w_003_315, w_004_991);
  nand2 I007_1599(w_007_1599, w_000_1873, w_003_045);
  and2 I007_1600(w_007_1600, w_004_1016, w_003_117);
  not1 I007_1601(w_007_1601, w_003_049);
  nand2 I007_1603(w_007_1603, w_002_192, w_001_137);
  nand2 I007_1605(w_007_1605, w_004_1092, w_002_405);
  nand2 I007_1606(w_007_1606, w_000_383, w_002_553);
  or2  I007_1615(w_007_1615, w_002_239, w_004_1073);
  nand2 I007_1616(w_007_1616, w_006_088, w_002_493);
  nand2 I007_1617(w_007_1617, w_002_310, w_006_042);
  and2 I007_1618(w_007_1618, w_006_060, w_006_067);
  or2  I007_1619(w_007_1619, w_006_142, w_003_224);
  and2 I007_1620(w_007_1620, w_006_171, w_000_1875);
  nand2 I008_002(w_008_002, w_007_393, w_001_206);
  not1 I008_003(w_008_003, w_004_1184);
  nand2 I008_005(w_008_005, w_001_1462, w_000_552);
  not1 I008_006(w_008_006, w_004_015);
  not1 I008_008(w_008_008, w_003_157);
  nand2 I008_009(w_008_009, w_001_768, w_002_339);
  or2  I008_010(w_008_010, w_002_277, w_005_1610);
  and2 I008_011(w_008_011, w_007_1508, w_004_1540);
  or2  I008_013(w_008_013, w_004_415, w_006_018);
  not1 I008_014(w_008_014, w_004_1116);
  and2 I008_015(w_008_015, w_007_290, w_007_417);
  not1 I008_016(w_008_016, w_001_756);
  and2 I008_017(w_008_017, w_003_105, w_001_1141);
  or2  I008_018(w_008_018, w_000_1002, w_006_261);
  not1 I008_019(w_008_019, w_003_064);
  not1 I008_020(w_008_020, w_001_1521);
  nand2 I008_021(w_008_021, w_000_463, w_001_292);
  nand2 I008_022(w_008_022, w_005_346, w_003_175);
  or2  I008_023(w_008_023, w_004_1850, w_002_050);
  not1 I008_024(w_008_024, w_005_1217);
  nand2 I008_025(w_008_025, w_002_358, w_000_1108);
  and2 I008_026(w_008_026, w_005_1358, w_004_765);
  or2  I008_027(w_008_027, w_005_638, w_000_1669);
  or2  I008_028(w_008_028, w_001_003, w_001_398);
  or2  I008_031(w_008_031, w_005_100, w_003_309);
  and2 I008_032(w_008_032, w_004_082, w_002_288);
  not1 I008_034(w_008_034, w_003_228);
  or2  I008_035(w_008_035, w_004_259, w_002_176);
  or2  I008_036(w_008_036, w_000_496, w_001_288);
  and2 I008_038(w_008_038, w_004_1618, w_000_1504);
  and2 I008_039(w_008_039, w_003_144, w_004_454);
  or2  I008_040(w_008_040, w_001_114, w_007_1084);
  not1 I008_041(w_008_041, w_004_1664);
  and2 I008_043(w_008_043, w_003_150, w_000_082);
  nand2 I008_044(w_008_044, w_001_1039, w_000_1454);
  nand2 I008_046(w_008_046, w_001_426, w_004_1755);
  and2 I008_047(w_008_047, w_004_839, w_002_092);
  or2  I008_049(w_008_049, w_001_064, w_004_1425);
  or2  I008_051(w_008_051, w_004_744, w_007_1298);
  nand2 I008_052(w_008_052, w_006_227, w_005_891);
  not1 I008_053(w_008_053, w_001_847);
  not1 I008_056(w_008_056, w_006_028);
  nand2 I008_058(w_008_058, w_004_1272, w_007_181);
  or2  I008_059(w_008_059, w_007_188, w_007_162);
  nand2 I008_060(w_008_060, w_002_092, w_006_065);
  or2  I008_061(w_008_061, w_005_316, w_005_169);
  or2  I008_062(w_008_062, w_005_539, w_003_300);
  or2  I008_064(w_008_064, w_006_024, w_002_195);
  or2  I008_065(w_008_065, w_007_236, w_001_1102);
  nand2 I008_066(w_008_066, w_004_1872, w_007_1506);
  or2  I008_067(w_008_067, w_000_871, w_000_214);
  nand2 I008_069(w_008_069, w_006_204, w_004_989);
  and2 I008_070(w_008_070, w_005_1099, w_000_1695);
  or2  I008_071(w_008_071, w_005_1638, w_005_1574);
  or2  I008_073(w_008_073, w_006_012, w_005_975);
  not1 I008_074(w_008_074, w_001_732);
  or2  I008_076(w_008_076, w_001_1475, w_001_478);
  not1 I008_077(w_008_077, w_001_526);
  nand2 I008_078(w_008_078, w_006_172, w_005_845);
  or2  I008_079(w_008_079, w_001_1408, w_006_085);
  nand2 I008_081(w_008_081, w_003_040, w_000_395);
  or2  I008_082(w_008_082, w_005_1233, w_007_214);
  nand2 I008_084(w_008_084, w_002_142, w_007_1127);
  or2  I008_085(w_008_085, w_000_1201, w_005_246);
  nand2 I008_087(w_008_087, w_005_1374, w_002_127);
  not1 I008_088(w_008_088, w_002_522);
  and2 I008_089(w_008_089, w_000_702, w_003_166);
  not1 I008_090(w_008_090, w_003_227);
  not1 I008_092(w_008_092, w_007_1043);
  not1 I008_093(w_008_093, w_000_385);
  or2  I008_094(w_008_094, w_006_188, w_000_541);
  or2  I008_095(w_008_095, w_006_247, w_002_213);
  not1 I008_096(w_008_096, w_007_1513);
  and2 I008_098(w_008_098, w_007_351, w_004_957);
  and2 I008_100(w_008_100, w_006_095, w_005_1591);
  or2  I008_102(w_008_102, w_002_212, w_007_063);
  not1 I008_103(w_008_103, w_006_176);
  and2 I008_104(w_008_104, w_003_268, w_005_1315);
  or2  I008_106(w_008_106, w_004_252, w_001_272);
  or2  I008_108(w_008_108, w_003_147, w_002_557);
  nand2 I008_109(w_008_109, w_002_003, w_006_056);
  or2  I008_110(w_008_110, w_002_016, w_002_091);
  nand2 I008_111(w_008_111, w_006_216, w_007_663);
  and2 I008_112(w_008_112, w_004_1771, w_000_581);
  not1 I008_114(w_008_114, w_005_314);
  or2  I008_115(w_008_115, w_007_546, w_004_1177);
  not1 I008_117(w_008_117, w_007_612);
  or2  I008_119(w_008_119, w_000_567, w_001_1221);
  or2  I008_122(w_008_122, w_005_1610, w_005_1255);
  and2 I008_123(w_008_123, w_002_346, w_002_005);
  or2  I008_124(w_008_124, w_007_1326, w_006_283);
  not1 I008_125(w_008_125, w_007_1603);
  or2  I008_126(w_008_126, w_000_1176, w_005_036);
  not1 I008_127(w_008_127, w_001_786);
  or2  I008_128(w_008_128, w_002_579, w_002_215);
  not1 I008_129(w_008_129, w_007_1365);
  nand2 I008_130(w_008_130, w_006_225, w_001_907);
  not1 I008_132(w_008_132, w_005_1362);
  or2  I008_133(w_008_133, w_000_755, w_001_880);
  or2  I008_134(w_008_134, w_005_1346, w_002_587);
  not1 I008_136(w_008_136, w_005_1229);
  nand2 I008_139(w_008_139, w_002_546, w_000_941);
  or2  I008_143(w_008_143, w_002_002, w_003_061);
  and2 I008_144(w_008_144, w_002_106, w_005_196);
  and2 I008_147(w_008_147, w_007_944, w_006_194);
  nand2 I008_148(w_008_148, w_002_149, w_002_511);
  not1 I008_151(w_008_151, w_006_139);
  nand2 I008_152(w_008_152, w_002_549, w_003_049);
  not1 I008_154(w_008_154, w_004_1107);
  or2  I008_156(w_008_156, w_005_623, w_001_1177);
  nand2 I008_157(w_008_157, w_002_379, w_003_097);
  or2  I008_158(w_008_158, w_001_1220, w_004_1115);
  not1 I008_160(w_008_160, w_002_554);
  and2 I008_162(w_008_162, w_002_443, w_006_325);
  or2  I008_163(w_008_163, w_003_060, w_002_124);
  and2 I008_164(w_008_164, w_004_503, w_007_158);
  and2 I008_165(w_008_165, w_000_1378, w_004_1243);
  and2 I008_166(w_008_166, w_003_072, w_003_309);
  nand2 I008_167(w_008_167, w_002_566, w_007_750);
  nand2 I008_168(w_008_168, w_004_552, w_002_232);
  not1 I008_170(w_008_170, w_006_042);
  not1 I008_172(w_008_172, w_005_1650);
  not1 I008_174(w_008_174, w_000_1260);
  and2 I008_175(w_008_175, w_002_097, w_006_165);
  nand2 I008_176(w_008_176, w_006_152, w_002_014);
  nand2 I008_177(w_008_177, w_000_1686, w_001_1642);
  and2 I008_180(w_008_180, w_000_1863, w_006_320);
  nand2 I008_181(w_008_181, w_007_1235, w_007_1245);
  and2 I008_182(w_008_182, w_006_100, w_000_224);
  nand2 I008_184(w_008_184, w_002_044, w_007_003);
  nand2 I008_185(w_008_185, w_006_009, w_000_1748);
  nand2 I008_186(w_008_186, w_001_013, w_007_927);
  or2  I008_187(w_008_187, w_002_002, w_000_1873);
  and2 I008_188(w_008_188, w_001_480, w_000_1876);
  not1 I008_190(w_008_190, w_004_1056);
  or2  I008_192(w_008_192, w_002_304, w_006_006);
  nand2 I008_193(w_008_193, w_007_019, w_002_302);
  or2  I008_195(w_008_195, w_002_258, w_001_1092);
  nand2 I008_196(w_008_196, w_001_745, w_000_511);
  and2 I008_197(w_008_197, w_004_005, w_006_031);
  not1 I008_198(w_008_198, w_004_009);
  not1 I008_199(w_008_199, w_002_016);
  or2  I008_200(w_008_200, w_001_387, w_004_1151);
  and2 I008_201(w_008_201, w_001_644, w_006_039);
  or2  I008_202(w_008_202, w_000_870, w_006_324);
  or2  I008_203(w_008_203, w_007_446, w_005_686);
  and2 I008_205(w_008_205, w_000_287, w_004_826);
  or2  I008_206(w_008_206, w_006_154, w_007_1103);
  or2  I008_207(w_008_207, w_003_255, w_002_424);
  nand2 I008_208(w_008_208, w_000_1035, w_001_504);
  or2  I008_209(w_008_209, w_007_205, w_006_111);
  nand2 I008_210(w_008_210, w_003_229, w_005_273);
  nand2 I008_211(w_008_211, w_005_765, w_002_214);
  nand2 I008_212(w_008_212, w_000_1656, w_001_1367);
  and2 I008_213(w_008_213, w_006_186, w_007_768);
  not1 I008_216(w_008_216, w_001_986);
  or2  I008_217(w_008_217, w_005_180, w_006_273);
  not1 I008_218(w_008_218, w_003_126);
  or2  I008_219(w_008_219, w_005_709, w_005_766);
  nand2 I008_222(w_008_222, w_006_013, w_003_223);
  not1 I008_224(w_008_224, w_007_415);
  and2 I008_225(w_008_225, w_000_098, w_007_1151);
  not1 I008_228(w_008_228, w_005_1002);
  and2 I008_230(w_008_230, w_006_247, w_002_162);
  or2  I008_231(w_008_231, w_001_076, w_001_401);
  or2  I008_233(w_008_233, w_003_193, w_000_1877);
  not1 I008_234(w_008_234, w_000_1457);
  and2 I008_235(w_008_235, w_005_459, w_005_937);
  not1 I008_236(w_008_236, w_006_195);
  not1 I008_237(w_008_237, w_004_171);
  and2 I008_238(w_008_238, w_003_208, w_005_246);
  nand2 I008_240(w_008_240, w_007_032, w_001_1276);
  nand2 I008_241(w_008_241, w_002_022, w_006_124);
  and2 I008_242(w_008_242, w_007_124, w_002_542);
  or2  I008_243(w_008_243, w_003_316, w_007_1046);
  nand2 I008_244(w_008_244, w_004_1217, w_003_263);
  not1 I008_245(w_008_245, w_001_126);
  and2 I008_246(w_008_246, w_000_657, w_007_935);
  or2  I008_247(w_008_247, w_000_564, w_004_130);
  and2 I008_248(w_008_248, w_002_012, w_005_897);
  nand2 I008_250(w_008_250, w_002_255, w_003_192);
  not1 I008_251(w_008_251, w_007_402);
  not1 I008_252(w_008_252, w_006_140);
  nand2 I008_253(w_008_253, w_006_208, w_003_023);
  nand2 I008_254(w_008_254, w_002_414, w_007_1142);
  and2 I008_256(w_008_256, w_007_905, w_003_050);
  and2 I008_257(w_008_257, w_005_577, w_007_1533);
  and2 I008_258(w_008_258, w_006_287, w_002_152);
  nand2 I008_259(w_008_259, w_005_1026, w_003_200);
  or2  I008_260(w_008_260, w_002_262, w_001_1089);
  or2  I008_261(w_008_261, w_005_658, w_000_347);
  or2  I008_262(w_008_262, w_004_1690, w_002_185);
  and2 I008_263(w_008_263, w_007_316, w_006_142);
  or2  I008_264(w_008_264, w_006_237, w_001_1264);
  or2  I008_266(w_008_266, w_005_1346, w_007_1487);
  and2 I008_268(w_008_268, w_000_1878, w_002_128);
  nand2 I008_269(w_008_269, w_007_097, w_007_1085);
  and2 I008_270(w_008_270, w_001_001, w_005_1650);
  nand2 I008_271(w_008_271, w_006_222, w_000_170);
  or2  I008_273(w_008_273, w_004_063, w_005_797);
  not1 I008_275(w_008_275, w_006_246);
  or2  I008_276(w_008_276, w_005_1007, w_005_1602);
  nand2 I008_277(w_008_277, w_006_261, w_004_104);
  and2 I008_278(w_008_278, w_003_102, w_000_1061);
  or2  I008_279(w_008_279, w_005_314, w_006_009);
  and2 I008_280(w_008_280, w_003_198, w_000_1350);
  and2 I008_281(w_008_281, w_003_314, w_006_121);
  and2 I008_282(w_008_282, w_003_286, w_007_544);
  or2  I008_285(w_008_285, w_005_1492, w_002_320);
  or2  I008_286(w_008_286, w_000_1276, w_006_283);
  not1 I008_288(w_008_288, w_001_587);
  and2 I008_289(w_008_289, w_003_187, w_000_1305);
  nand2 I008_290(w_008_290, w_000_1879, w_002_539);
  and2 I008_293(w_008_293, w_005_369, w_004_1105);
  nand2 I008_294(w_008_294, w_007_267, w_005_041);
  not1 I008_296(w_008_296, w_002_174);
  not1 I008_297(w_008_297, w_003_123);
  nand2 I008_298(w_008_298, w_005_189, w_006_325);
  not1 I008_300(w_008_300, w_006_196);
  not1 I008_301(w_008_301, w_002_377);
  not1 I008_303(w_008_303, w_005_591);
  nand2 I008_306(w_008_306, w_004_962, w_004_798);
  nand2 I008_308(w_008_308, w_006_300, w_003_237);
  and2 I008_310(w_008_310, w_000_1379, w_004_012);
  nand2 I008_312(w_008_312, w_002_572, w_002_498);
  nand2 I008_314(w_008_314, w_004_1833, w_007_1567);
  or2  I008_315(w_008_315, w_005_555, w_000_1306);
  or2  I008_316(w_008_316, w_003_093, w_006_011);
  and2 I008_317(w_008_317, w_002_125, w_007_405);
  or2  I008_318(w_008_318, w_002_547, w_005_460);
  or2  I008_319(w_008_319, w_007_498, w_007_1294);
  and2 I008_324(w_008_324, w_006_273, w_001_771);
  and2 I008_326(w_008_326, w_007_805, w_003_135);
  nand2 I008_327(w_008_327, w_004_213, w_006_329);
  nand2 I008_330(w_008_330, w_005_121, w_004_1487);
  and2 I008_332(w_008_332, w_002_239, w_002_193);
  not1 I008_336(w_008_336, w_006_084);
  not1 I008_342(w_008_342, w_004_941);
  nand2 I008_343(w_008_343, w_001_1066, w_001_1476);
  and2 I008_344(w_008_344, w_006_018, w_003_318);
  and2 I008_345(w_008_345, w_006_166, w_001_522);
  nand2 I008_346(w_008_346, w_007_315, w_002_229);
  nand2 I008_348(w_008_348, w_003_036, w_007_1303);
  not1 I008_349(w_008_349, w_003_245);
  nand2 I008_351(w_008_351, w_005_1467, w_002_511);
  nand2 I008_352(w_008_352, w_000_1241, w_000_915);
  and2 I008_353(w_008_353, w_000_1230, w_002_579);
  not1 I008_355(w_008_355, w_007_359);
  nand2 I008_359(w_008_359, w_004_552, w_004_516);
  nand2 I008_360(w_008_360, w_006_283, w_004_555);
  not1 I008_362(w_008_362, w_000_1462);
  nand2 I008_364(w_008_364, w_005_1235, w_003_170);
  or2  I008_365(w_008_365, w_007_1407, w_000_1019);
  nand2 I008_368(w_008_368, w_007_673, w_006_130);
  nand2 I008_369(w_008_369, w_007_969, w_002_554);
  nand2 I008_370(w_008_370, w_005_790, w_007_698);
  nand2 I008_372(w_008_372, w_007_124, w_003_107);
  nand2 I008_373(w_008_373, w_002_340, w_005_1109);
  and2 I008_374(w_008_374, w_000_1588, w_005_1431);
  and2 I008_376(w_008_376, w_007_1168, w_006_310);
  not1 I008_379(w_008_379, w_005_223);
  or2  I008_380(w_008_380, w_001_234, w_000_927);
  and2 I008_381(w_008_381, w_005_1276, w_000_786);
  or2  I008_382(w_008_382, w_007_233, w_002_021);
  and2 I008_384(w_008_384, w_007_1049, w_004_624);
  or2  I008_386(w_008_386, w_007_793, w_004_191);
  nand2 I008_390(w_008_390, w_001_213, w_003_280);
  and2 I008_393(w_008_393, w_006_170, w_000_1701);
  nand2 I008_394(w_008_394, w_004_1089, w_007_632);
  and2 I008_395(w_008_395, w_005_1052, w_007_1302);
  not1 I008_396(w_008_396, w_000_332);
  nand2 I008_399(w_008_399, w_004_042, w_007_778);
  and2 I008_400(w_008_400, w_007_479, w_007_1251);
  and2 I008_401(w_008_401, w_007_236, w_000_068);
  and2 I008_402(w_008_402, w_000_1722, w_006_288);
  not1 I008_404(w_008_404, w_000_346);
  not1 I008_407(w_008_407, w_001_673);
  not1 I008_408(w_008_408, w_000_909);
  not1 I008_412(w_008_412, w_005_1065);
  nand2 I008_413(w_008_413, w_000_767, w_004_1349);
  and2 I008_415(w_008_415, w_004_1108, w_000_1401);
  not1 I008_417(w_008_417, w_005_537);
  not1 I008_418(w_008_418, w_001_1288);
  or2  I008_419(w_008_419, w_007_230, w_002_206);
  not1 I008_420(w_008_420, w_003_319);
  not1 I008_421(w_008_421, w_000_669);
  not1 I008_422(w_008_422, w_007_136);
  nand2 I008_423(w_008_423, w_007_628, w_003_087);
  or2  I008_424(w_008_424, w_002_200, w_003_052);
  nand2 I008_425(w_008_425, w_006_097, w_001_040);
  not1 I008_426(w_008_426, w_001_1629);
  not1 I008_428(w_008_428, w_001_1416);
  nand2 I008_429(w_008_429, w_006_118, w_002_558);
  nand2 I008_431(w_008_431, w_003_117, w_002_312);
  and2 I008_433(w_008_433, w_007_021, w_005_131);
  or2  I008_434(w_008_434, w_007_1472, w_007_288);
  and2 I008_435(w_008_435, w_002_358, w_006_069);
  and2 I008_436(w_008_436, w_003_151, w_006_332);
  and2 I008_437(w_008_437, w_005_1368, w_006_287);
  and2 I008_438(w_008_438, w_003_312, w_001_121);
  not1 I008_442(w_008_442, w_005_528);
  and2 I008_443(w_008_443, w_002_014, w_000_1545);
  not1 I008_444(w_008_444, w_004_025);
  nand2 I008_445(w_008_445, w_004_943, w_006_044);
  nand2 I008_447(w_008_447, w_007_243, w_003_293);
  and2 I008_449(w_008_449, w_000_1378, w_002_519);
  nand2 I008_450(w_008_450, w_002_101, w_001_1238);
  not1 I008_453(w_008_453, w_004_1711);
  or2  I008_454(w_008_454, w_003_010, w_005_1656);
  or2  I008_455(w_008_455, w_007_080, w_001_519);
  nand2 I008_456(w_008_456, w_004_1038, w_002_004);
  not1 I008_457(w_008_457, w_004_1837);
  or2  I008_459(w_008_459, w_002_042, w_003_283);
  and2 I008_460(w_008_460, w_007_322, w_005_675);
  and2 I008_461(w_008_461, w_002_089, w_005_121);
  nand2 I008_463(w_008_463, w_001_665, w_001_725);
  not1 I008_464(w_008_464, w_007_1148);
  and2 I008_465(w_008_465, w_004_678, w_001_438);
  or2  I008_470(w_008_470, w_007_146, w_006_233);
  nand2 I008_472(w_008_472, w_007_798, w_004_1086);
  nand2 I008_473(w_008_473, w_000_1759, w_003_124);
  nand2 I008_474(w_008_474, w_001_026, w_003_202);
  and2 I008_475(w_008_475, w_000_1880, w_002_341);
  or2  I008_477(w_008_477, w_005_386, w_005_1392);
  and2 I008_479(w_008_479, w_005_1478, w_003_165);
  or2  I008_480(w_008_480, w_007_209, w_000_1344);
  and2 I008_481(w_008_481, w_003_186, w_000_756);
  nand2 I008_484(w_008_484, w_004_1594, w_000_581);
  and2 I008_485(w_008_485, w_000_973, w_005_1133);
  not1 I008_488(w_008_488, w_001_424);
  or2  I008_489(w_008_489, w_004_1873, w_006_174);
  nand2 I008_490(w_008_490, w_005_1103, w_002_454);
  or2  I008_491(w_008_491, w_002_575, w_006_210);
  or2  I008_495(w_008_495, w_006_237, w_007_1469);
  not1 I008_500(w_008_500, w_006_111);
  nand2 I008_501(w_008_501, w_004_920, w_001_1122);
  or2  I008_502(w_008_502, w_000_943, w_000_1182);
  not1 I008_504(w_008_504, w_007_360);
  or2  I008_506(w_008_506, w_006_289, w_000_1638);
  and2 I008_507(w_008_507, w_006_266, w_007_1284);
  nand2 I008_511(w_008_511, w_006_221, w_001_1047);
  nand2 I008_513(w_008_513, w_003_176, w_005_026);
  nand2 I008_515(w_008_515, w_006_169, w_003_319);
  nand2 I008_518(w_008_518, w_001_033, w_000_772);
  or2  I008_519(w_008_519, w_003_047, w_006_089);
  or2  I008_521(w_008_521, w_002_346, w_003_053);
  not1 I008_524(w_008_524, w_006_091);
  or2  I008_525(w_008_525, w_007_190, w_001_139);
  and2 I008_526(w_008_526, w_004_1466, w_002_345);
  and2 I008_527(w_008_527, w_005_708, w_006_157);
  nand2 I008_530(w_008_530, w_007_491, w_001_770);
  or2  I008_531(w_008_531, w_007_1214, w_002_196);
  and2 I008_533(w_008_533, w_002_155, w_000_1839);
  not1 I008_534(w_008_534, w_007_092);
  not1 I008_537(w_008_537, w_003_039);
  nand2 I008_538(w_008_538, w_002_385, w_006_153);
  nand2 I008_540(w_008_540, w_004_975, w_000_588);
  or2  I008_541(w_008_541, w_007_656, w_001_1454);
  not1 I008_543(w_008_543, w_002_431);
  and2 I008_544(w_008_544, w_005_303, w_007_1104);
  and2 I008_546(w_008_546, w_003_120, w_003_143);
  nand2 I008_547(w_008_547, w_003_123, w_000_1834);
  and2 I008_549(w_008_549, w_003_138, w_006_157);
  not1 I008_550(w_008_550, w_002_023);
  and2 I008_551(w_008_551, w_002_315, w_000_1647);
  and2 I008_552(w_008_552, w_001_204, w_000_1881);
  nand2 I008_553(w_008_553, w_003_083, w_006_095);
  nand2 I008_554(w_008_554, w_007_001, w_003_048);
  not1 I008_555(w_008_555, w_007_108);
  nand2 I008_556(w_008_556, w_002_292, w_005_1328);
  not1 I008_560(w_008_560, w_002_351);
  and2 I008_562(w_008_562, w_006_151, w_005_040);
  not1 I008_563(w_008_563, w_001_181);
  or2  I008_564(w_008_564, w_007_181, w_001_556);
  not1 I008_566(w_008_566, w_000_1044);
  and2 I008_567(w_008_567, w_000_1882, w_006_031);
  or2  I008_569(w_008_569, w_006_343, w_006_254);
  not1 I008_570(w_008_570, w_007_126);
  and2 I008_572(w_008_572, w_004_1788, w_007_438);
  not1 I008_573(w_008_573, w_007_1482);
  not1 I008_574(w_008_574, w_000_1728);
  and2 I008_577(w_008_577, w_000_1883, w_004_262);
  and2 I008_578(w_008_578, w_003_257, w_004_518);
  or2  I008_579(w_008_579, w_000_306, w_000_1550);
  and2 I008_580(w_008_580, w_007_1384, w_002_007);
  not1 I008_584(w_008_584, w_005_1445);
  not1 I008_589(w_008_589, w_001_899);
  and2 I008_591(w_008_591, w_003_201, w_005_152);
  and2 I008_593(w_008_593, w_001_278, w_001_537);
  or2  I008_594(w_008_594, w_004_025, w_004_661);
  nand2 I008_595(w_008_595, w_007_212, w_001_238);
  or2  I008_597(w_008_597, w_007_1474, w_006_301);
  not1 I008_599(w_008_599, w_007_299);
  nand2 I008_602(w_008_602, w_002_491, w_002_198);
  and2 I008_603(w_008_603, w_003_293, w_001_653);
  and2 I008_605(w_008_605, w_001_1140, w_007_628);
  and2 I008_608(w_008_608, w_005_1397, w_003_039);
  and2 I008_609(w_008_609, w_006_157, w_005_1449);
  nand2 I008_610(w_008_610, w_006_102, w_007_622);
  or2  I008_611(w_008_611, w_003_136, w_001_772);
  or2  I008_612(w_008_612, w_000_1753, w_007_847);
  not1 I008_615(w_008_615, w_006_043);
  and2 I008_616(w_008_616, w_003_204, w_007_114);
  nand2 I008_618(w_008_618, w_002_255, w_005_203);
  not1 I008_619(w_008_619, w_005_1631);
  or2  I008_620(w_008_620, w_004_664, w_006_283);
  or2  I008_621(w_008_621, w_007_1179, w_003_110);
  or2  I008_622(w_008_622, w_000_333, w_000_067);
  or2  I008_624(w_008_624, w_006_246, w_005_1088);
  not1 I008_626(w_008_626, w_002_490);
  not1 I008_627(w_008_627, w_000_407);
  and2 I008_628(w_008_628, w_000_1586, w_003_078);
  nand2 I008_632(w_008_632, w_003_122, w_005_610);
  nand2 I008_633(w_008_633, w_005_1561, w_001_1161);
  not1 I008_635(w_008_635, w_002_280);
  not1 I008_638(w_008_638, w_000_1477);
  nand2 I008_639(w_008_639, w_007_1328, w_002_094);
  not1 I008_644(w_008_644, w_005_585);
  or2  I008_645(w_008_645, w_005_1667, w_002_400);
  not1 I008_646(w_008_646, w_001_674);
  and2 I008_651(w_008_651, w_004_534, w_005_234);
  nand2 I008_652(w_008_652, w_002_147, w_001_243);
  nand2 I008_653(w_008_653, w_002_013, w_000_310);
  and2 I008_656(w_008_656, w_006_130, w_005_1525);
  or2  I008_657(w_008_657, w_002_409, w_001_292);
  and2 I008_659(w_008_659, w_004_1494, w_000_167);
  or2  I008_660(w_008_660, w_000_477, w_003_248);
  not1 I008_661(w_008_661, w_004_828);
  and2 I008_662(w_008_662, w_001_1680, w_001_919);
  nand2 I008_663(w_008_663, w_006_100, w_004_400);
  not1 I008_664(w_008_664, w_006_046);
  not1 I008_666(w_008_666, w_005_192);
  not1 I008_668(w_008_668, w_001_042);
  nand2 I008_670(w_008_670, w_000_889, w_003_249);
  or2  I008_673(w_008_673, w_006_045, w_003_276);
  not1 I008_674(w_008_674, w_006_242);
  not1 I008_675(w_008_675, w_007_064);
  not1 I008_677(w_008_677, w_006_317);
  or2  I008_678(w_008_678, w_007_230, w_004_1182);
  nand2 I008_679(w_008_679, w_007_253, w_002_230);
  not1 I008_680(w_008_680, w_006_261);
  or2  I008_681(w_008_681, w_003_168, w_005_074);
  nand2 I008_682(w_008_682, w_000_1795, w_006_272);
  not1 I008_683(w_008_683, w_002_173);
  or2  I008_684(w_008_684, w_006_113, w_007_235);
  nand2 I008_685(w_008_685, w_007_441, w_003_293);
  and2 I008_686(w_008_686, w_002_263, w_006_258);
  and2 I008_688(w_008_688, w_004_1638, w_007_996);
  or2  I008_689(w_008_689, w_005_1612, w_004_895);
  or2  I008_691(w_008_691, w_004_1899, w_002_055);
  or2  I008_692(w_008_692, w_007_1209, w_004_429);
  nand2 I008_694(w_008_694, w_003_020, w_001_1498);
  nand2 I008_696(w_008_696, w_000_499, w_004_262);
  not1 I008_698(w_008_698, w_004_959);
  nand2 I008_699(w_008_699, w_000_1740, w_007_1042);
  not1 I008_702(w_008_702, w_005_1166);
  not1 I008_703(w_008_703, w_004_1773);
  nand2 I008_704(w_008_704, w_007_170, w_001_407);
  nand2 I008_705(w_008_705, w_003_027, w_007_1229);
  nand2 I008_706(w_008_706, w_006_225, w_000_1235);
  and2 I008_707(w_008_707, w_002_022, w_002_216);
  and2 I008_709(w_008_709, w_004_804, w_002_580);
  not1 I008_712(w_008_712, w_003_247);
  not1 I008_713(w_008_713, w_001_1432);
  not1 I008_714(w_008_714, w_004_896);
  not1 I008_717(w_008_717, w_004_492);
  not1 I008_718(w_008_718, w_006_266);
  not1 I008_719(w_008_719, w_002_198);
  not1 I008_720(w_008_720, w_005_770);
  and2 I008_721(w_008_721, w_000_1885, w_002_472);
  not1 I008_727(w_008_727, w_000_1310);
  not1 I008_728(w_008_728, w_000_1288);
  or2  I008_729(w_008_729, w_002_214, w_001_1449);
  or2  I008_731(w_008_731, w_002_451, w_006_072);
  or2  I008_732(w_008_732, w_005_051, w_002_423);
  or2  I008_734(w_008_734, w_006_335, w_003_278);
  nand2 I008_735(w_008_735, w_000_985, w_001_946);
  nand2 I008_738(w_008_738, w_004_1388, w_005_073);
  nand2 I008_739(w_008_739, w_007_036, w_003_301);
  or2  I008_741(w_008_741, w_000_661, w_004_1832);
  not1 I008_742(w_008_742, w_005_1130);
  and2 I008_743(w_008_743, w_004_382, w_000_1702);
  or2  I008_744(w_008_744, w_006_274, w_000_1882);
  nand2 I008_745(w_008_745, w_005_307, w_006_221);
  and2 I008_747(w_008_747, w_000_1209, w_005_672);
  nand2 I008_748(w_008_748, w_001_504, w_005_438);
  nand2 I008_749(w_008_749, w_006_083, w_001_1622);
  or2  I008_750(w_008_750, w_006_108, w_004_1895);
  not1 I008_751(w_008_751, w_003_108);
  not1 I008_752(w_008_752, w_001_1633);
  not1 I008_753(w_008_753, w_003_211);
  and2 I008_755(w_008_755, w_005_1142, w_001_108);
  nand2 I008_756(w_008_756, w_000_1785, w_001_091);
  or2  I008_758(w_008_758, w_004_1744, w_000_1886);
  nand2 I008_759(w_008_759, w_004_011, w_005_1446);
  nand2 I008_760(w_008_760, w_000_1609, w_004_565);
  or2  I008_761(w_008_761, w_002_054, w_005_308);
  not1 I008_762(w_008_762, w_007_157);
  not1 I008_763(w_008_763, w_007_1566);
  nand2 I008_764(w_008_764, w_002_073, w_007_1134);
  not1 I008_765(w_008_765, w_004_879);
  not1 I008_766(w_008_766, w_007_490);
  not1 I008_767(w_008_767, w_004_799);
  or2  I008_769(w_008_769, w_003_017, w_001_038);
  or2  I008_770(w_008_770, w_004_1831, w_006_114);
  not1 I008_771(w_008_771, w_005_1609);
  and2 I008_772(w_008_772, w_006_089, w_007_1368);
  or2  I008_773(w_008_773, w_006_002, w_004_062);
  and2 I008_776(w_008_776, w_006_230, w_005_295);
  and2 I008_778(w_008_778, w_000_1421, w_005_406);
  not1 I008_779(w_008_779, w_004_126);
  not1 I008_783(w_008_783, w_007_137);
  or2  I008_785(w_008_785, w_002_244, w_002_352);
  not1 I008_787(w_008_787, w_003_183);
  or2  I008_788(w_008_788, w_005_133, w_001_1560);
  nand2 I008_790(w_008_790, w_000_984, w_006_113);
  or2  I008_791(w_008_791, w_004_039, w_003_183);
  and2 I008_793(w_008_793, w_003_188, w_005_1026);
  not1 I008_794(w_008_794, w_000_1162);
  and2 I008_795(w_008_795, w_006_290, w_001_044);
  or2  I008_796(w_008_796, w_004_1800, w_000_181);
  not1 I008_798(w_008_798, w_001_170);
  nand2 I008_799(w_008_799, w_007_458, w_002_181);
  and2 I008_801(w_008_801, w_000_744, w_004_1442);
  and2 I008_802(w_008_802, w_002_170, w_001_872);
  or2  I008_804(w_008_804, w_005_1329, w_006_088);
  nand2 I008_805(w_008_805, w_007_610, w_006_222);
  and2 I008_806(w_008_806, w_000_131, w_003_061);
  or2  I008_807(w_008_807, w_007_285, w_005_1123);
  nand2 I008_808(w_008_808, w_005_262, w_004_1478);
  not1 I008_809(w_008_809, w_001_947);
  nand2 I008_810(w_008_810, w_007_598, w_000_1828);
  nand2 I008_811(w_008_811, w_006_268, w_006_054);
  and2 I008_813(w_008_813, w_006_289, w_005_1637);
  nand2 I008_815(w_008_815, w_002_421, w_005_988);
  and2 I008_817(w_008_817, w_005_851, w_004_275);
  or2  I008_818(w_008_818, w_003_215, w_005_375);
  nand2 I008_819(w_008_819, w_005_178, w_005_338);
  nand2 I008_821(w_008_821, w_003_205, w_000_1192);
  or2  I008_823(w_008_823, w_004_1533, w_004_1329);
  nand2 I008_825(w_008_825, w_003_112, w_001_120);
  and2 I008_829(w_008_829, w_002_322, w_001_1406);
  nand2 I008_830(w_008_830, w_001_828, w_003_161);
  nand2 I008_831(w_008_831, w_007_101, w_007_712);
  and2 I008_833(w_008_833, w_001_741, w_007_725);
  nand2 I008_836(w_008_836, w_000_595, w_007_1460);
  nand2 I008_838(w_008_838, w_007_544, w_007_1473);
  or2  I008_841(w_008_841, w_005_228, w_005_1286);
  or2  I008_847(w_008_847, w_006_321, w_007_187);
  and2 I008_850(w_008_850, w_005_1267, w_002_014);
  nand2 I008_851(w_008_851, w_003_274, w_003_131);
  nand2 I008_853(w_008_853, w_001_061, w_005_1216);
  and2 I008_856(w_008_856, w_003_278, w_004_496);
  or2  I008_857(w_008_857, w_007_1456, w_000_1690);
  not1 I008_858(w_008_858, w_003_142);
  or2  I008_861(w_008_861, w_003_192, w_006_198);
  nand2 I008_862(w_008_862, w_004_1335, w_007_031);
  not1 I009_000(w_009_000, w_004_695);
  not1 I009_001(w_009_001, w_004_1863);
  not1 I009_002(w_009_002, w_008_180);
  nand2 I009_003(w_009_003, w_000_1871, w_006_053);
  not1 I009_004(w_009_004, w_003_009);
  or2  I009_005(w_009_005, w_007_360, w_008_480);
  nand2 I009_006(w_009_006, w_001_1531, w_003_136);
  and2 I009_007(w_009_007, w_000_218, w_005_612);
  not1 I009_008(w_009_008, w_002_204);
  or2  I009_009(w_009_009, w_003_285, w_007_855);
  and2 I009_010(w_009_010, w_005_1078, w_007_098);
  and2 I009_011(w_009_011, w_002_051, w_001_519);
  nand2 I009_012(w_009_012, w_000_1864, w_007_038);
  and2 I009_013(w_009_013, w_001_116, w_007_1524);
  and2 I009_014(w_009_014, w_004_137, w_004_435);
  nand2 I009_015(w_009_015, w_003_149, w_001_1226);
  and2 I009_016(w_009_016, w_002_573, w_004_136);
  not1 I009_017(w_009_017, w_005_170);
  or2  I009_018(w_009_018, w_006_001, w_003_190);
  not1 I009_019(w_009_019, w_001_181);
  not1 I009_020(w_009_020, w_000_1887);
  not1 I009_021(w_009_021, w_000_364);
  not1 I009_022(w_009_022, w_004_710);
  or2  I009_023(w_009_023, w_004_1114, w_000_1848);
  and2 I009_024(w_009_024, w_008_659, w_006_098);
  and2 I009_025(w_009_025, w_000_722, w_002_153);
  nand2 I009_026(w_009_026, w_007_804, w_007_154);
  and2 I009_027(w_009_027, w_000_432, w_007_370);
  not1 I009_028(w_009_028, w_005_734);
  or2  I009_029(w_009_029, w_000_1797, w_008_692);
  nand2 I009_030(w_009_030, w_008_027, w_006_077);
  or2  I009_031(w_009_031, w_001_1551, w_002_080);
  or2  I009_032(w_009_032, w_004_015, w_008_266);
  nand2 I009_033(w_009_033, w_004_1774, w_000_918);
  not1 I009_034(w_009_034, w_005_1288);
  or2  I009_035(w_009_035, w_000_023, w_007_800);
  and2 I009_036(w_009_036, w_006_021, w_006_086);
  not1 I009_037(w_009_037, w_001_915);
  and2 I009_038(w_009_038, w_000_818, w_005_472);
  and2 I009_039(w_009_039, w_000_839, w_000_867);
  not1 I009_040(w_009_040, w_004_993);
  or2  I009_041(w_009_041, w_006_176, w_007_518);
  or2  I009_042(w_009_042, w_005_893, w_007_1570);
  or2  I009_043(w_009_043, w_002_280, w_001_1581);
  not1 I009_044(w_009_044, w_000_848);
  not1 I009_045(w_009_045, w_001_1667);
  and2 I009_046(w_009_046, w_008_246, w_003_087);
  and2 I009_047(w_009_047, w_004_769, w_006_299);
  nand2 I009_048(w_009_048, w_001_1579, w_004_1652);
  and2 I009_049(w_009_049, w_000_898, w_000_1888);
  nand2 I009_050(w_009_050, w_003_274, w_002_558);
  or2  I009_051(w_009_051, w_002_353, w_007_1097);
  and2 I009_052(w_009_052, w_001_665, w_007_1299);
  and2 I009_053(w_009_053, w_000_1629, w_006_275);
  and2 I009_054(w_009_054, w_005_1409, w_006_038);
  or2  I009_055(w_009_055, w_008_078, w_008_028);
  or2  I009_056(w_009_056, w_000_1599, w_000_1091);
  nand2 I009_057(w_009_057, w_006_061, w_008_276);
  nand2 I009_058(w_009_058, w_002_112, w_005_1663);
  nand2 I009_059(w_009_059, w_005_738, w_005_1529);
  or2  I009_060(w_009_060, w_006_226, w_005_636);
  and2 I009_061(w_009_061, w_007_1565, w_003_243);
  or2  I009_062(w_009_062, w_008_100, w_000_147);
  or2  I009_063(w_009_063, w_004_1532, w_000_456);
  and2 I009_064(w_009_064, w_004_636, w_002_470);
  and2 I009_065(w_009_065, w_008_589, w_006_043);
  nand2 I009_066(w_009_066, w_007_475, w_002_100);
  and2 I009_067(w_009_067, w_007_774, w_000_385);
  not1 I009_068(w_009_068, w_008_680);
  and2 I009_069(w_009_069, w_006_044, w_002_087);
  and2 I009_070(w_009_070, w_000_677, w_004_1415);
  not1 I009_071(w_009_071, w_004_1885);
  not1 I009_072(w_009_072, w_003_091);
  and2 I009_073(w_009_073, w_005_1026, w_004_1594);
  and2 I009_074(w_009_074, w_006_018, w_001_1121);
  nand2 I009_075(w_009_075, w_007_1451, w_003_272);
  and2 I009_076(w_009_076, w_000_1308, w_005_125);
  or2  I009_077(w_009_077, w_005_478, w_000_966);
  and2 I009_078(w_009_078, w_003_243, w_000_1025);
  not1 I009_079(w_009_079, w_006_152);
  and2 I009_080(w_009_080, w_000_090, w_000_982);
  and2 I009_081(w_009_081, w_001_103, w_007_009);
  nand2 I009_082(w_009_082, w_001_897, w_000_227);
  not1 I009_083(w_009_083, w_005_379);
  nand2 I009_084(w_009_084, w_008_344, w_004_490);
  or2  I009_085(w_009_085, w_007_069, w_003_200);
  nand2 I009_086(w_009_086, w_008_246, w_006_277);
  not1 I009_087(w_009_087, w_007_1603);
  not1 I009_088(w_009_088, w_008_841);
  or2  I009_089(w_009_089, w_006_237, w_006_021);
  and2 I009_090(w_009_090, w_005_1259, w_001_1351);
  not1 I009_091(w_009_091, w_000_913);
  nand2 I009_092(w_009_092, w_004_618, w_005_812);
  not1 I009_093(w_009_093, w_008_455);
  and2 I009_094(w_009_094, w_001_723, w_002_503);
  nand2 I009_095(w_009_095, w_003_069, w_004_1054);
  not1 I009_096(w_009_096, w_001_1020);
  nand2 I009_097(w_009_097, w_001_856, w_007_1618);
  not1 I009_098(w_009_098, w_000_1025);
  nand2 I009_099(w_009_099, w_001_848, w_000_174);
  or2  I009_100(w_009_100, w_002_366, w_005_979);
  and2 I009_101(w_009_101, w_006_326, w_007_176);
  or2  I009_102(w_009_102, w_001_597, w_005_205);
  and2 I009_103(w_009_103, w_007_900, w_004_1495);
  and2 I009_104(w_009_104, w_003_185, w_000_314);
  not1 I009_105(w_009_105, w_005_195);
  not1 I009_106(w_009_106, w_003_044);
  and2 I009_107(w_009_107, w_005_1357, w_006_155);
  or2  I009_108(w_009_108, w_003_297, w_005_955);
  not1 I009_109(w_009_109, w_004_1905);
  or2  I009_110(w_009_110, w_006_341, w_008_524);
  and2 I009_111(w_009_111, w_005_633, w_001_185);
  or2  I009_112(w_009_114, w_008_460, w_009_113);
  or2  I009_113(w_009_115, w_009_114, w_004_462);
  nand2 I009_114(w_009_116, w_009_115, w_008_176);
  nand2 I009_115(w_009_117, w_009_116, w_003_077);
  and2 I009_116(w_009_118, w_009_131, w_009_117);
  nand2 I009_117(w_009_119, w_008_703, w_009_118);
  nand2 I009_118(w_009_120, w_009_119, w_008_611);
  and2 I009_119(w_009_113, w_009_120, w_001_722);
  and2 I009_120(w_009_125, w_009_124, w_007_166);
  or2  I009_121(w_009_126, w_009_125, w_002_270);
  nand2 I009_122(w_009_127, w_002_368, w_009_126);
  not1 I009_123(w_009_128, w_009_127);
  not1 I009_124(w_009_129, w_009_128);
  not1 I009_125(w_009_124, w_009_118);
  and2 I009_126(w_009_131, w_002_481, w_009_129);
  not1 I010_001(w_010_001, w_004_1534);
  nand2 I010_002(w_010_002, w_001_641, w_002_210);
  or2  I010_003(w_010_003, w_002_183, w_008_185);
  not1 I010_004(w_010_004, w_003_211);
  not1 I010_005(w_010_005, w_006_028);
  nand2 I010_006(w_010_006, w_005_1436, w_004_1294);
  not1 I010_007(w_010_007, w_009_008);
  not1 I010_008(w_010_008, w_009_047);
  and2 I010_009(w_010_009, w_001_233, w_005_183);
  and2 I010_010(w_010_010, w_006_041, w_005_1669);
  or2  I010_011(w_010_011, w_004_398, w_007_1258);
  nand2 I010_012(w_010_012, w_001_1053, w_000_1827);
  and2 I010_013(w_010_013, w_007_1264, w_000_1851);
  not1 I010_014(w_010_014, w_001_643);
  and2 I010_015(w_010_015, w_000_1155, w_000_1744);
  nand2 I010_017(w_010_017, w_004_1379, w_000_1133);
  and2 I010_018(w_010_018, w_006_155, w_006_005);
  nand2 I010_019(w_010_019, w_007_1130, w_007_154);
  not1 I010_020(w_010_020, w_004_1770);
  not1 I010_021(w_010_021, w_007_1360);
  or2  I010_022(w_010_022, w_001_262, w_002_380);
  or2  I010_023(w_010_023, w_008_646, w_008_222);
  or2  I010_024(w_010_024, w_002_144, w_001_036);
  and2 I010_025(w_010_025, w_000_1609, w_004_1747);
  and2 I010_026(w_010_026, w_001_877, w_001_978);
  nand2 I010_027(w_010_027, w_005_748, w_003_213);
  or2  I010_028(w_010_028, w_004_226, w_003_048);
  not1 I010_029(w_010_029, w_006_318);
  and2 I010_030(w_010_030, w_005_959, w_004_399);
  nand2 I010_031(w_010_031, w_007_477, w_001_787);
  nand2 I010_032(w_010_032, w_006_198, w_003_219);
  nand2 I010_033(w_010_033, w_005_194, w_000_892);
  not1 I010_034(w_010_034, w_003_097);
  nand2 I010_035(w_010_035, w_000_1635, w_002_038);
  or2  I010_036(w_010_036, w_001_1045, w_004_1626);
  and2 I010_037(w_010_037, w_000_377, w_009_085);
  nand2 I010_038(w_010_038, w_000_1097, w_004_638);
  nand2 I010_039(w_010_039, w_007_1178, w_009_082);
  nand2 I010_040(w_010_040, w_009_095, w_007_925);
  and2 I010_041(w_010_041, w_008_225, w_004_1293);
  or2  I010_042(w_010_042, w_005_1464, w_002_563);
  not1 I010_043(w_010_043, w_008_078);
  nand2 I010_044(w_010_044, w_009_021, w_006_020);
  not1 I010_045(w_010_045, w_000_658);
  or2  I010_046(w_010_046, w_000_188, w_008_819);
  and2 I010_047(w_010_047, w_000_1683, w_007_1415);
  and2 I010_048(w_010_048, w_006_002, w_006_011);
  nand2 I010_049(w_010_049, w_003_195, w_002_471);
  or2  I010_050(w_010_050, w_002_360, w_008_062);
  or2  I010_051(w_010_051, w_007_434, w_005_152);
  or2  I010_054(w_010_054, w_000_1098, w_001_1288);
  and2 I010_055(w_010_055, w_009_003, w_002_535);
  not1 I010_056(w_010_056, w_004_1140);
  nand2 I010_057(w_010_057, w_008_635, w_004_780);
  not1 I010_058(w_010_058, w_001_1566);
  or2  I010_059(w_010_059, w_000_1011, w_006_096);
  and2 I010_060(w_010_060, w_000_1586, w_001_363);
  nand2 I010_061(w_010_061, w_003_214, w_009_092);
  not1 I010_062(w_010_062, w_008_783);
  not1 I010_063(w_010_063, w_001_300);
  and2 I010_064(w_010_064, w_001_1505, w_005_139);
  or2  I010_065(w_010_065, w_007_928, w_002_454);
  or2  I010_066(w_010_066, w_005_142, w_008_262);
  or2  I010_067(w_010_067, w_000_713, w_006_295);
  and2 I010_068(w_010_068, w_009_109, w_009_101);
  and2 I010_069(w_010_069, w_000_469, w_000_441);
  nand2 I010_070(w_010_070, w_007_755, w_006_154);
  or2  I010_071(w_010_071, w_008_761, w_009_038);
  and2 I010_073(w_010_073, w_001_052, w_001_987);
  not1 I010_074(w_010_074, w_002_229);
  nand2 I010_076(w_010_076, w_008_117, w_002_203);
  and2 I010_077(w_010_077, w_001_671, w_003_049);
  and2 I010_078(w_010_078, w_002_503, w_004_904);
  or2  I010_079(w_010_079, w_000_1067, w_009_006);
  or2  I010_080(w_010_080, w_001_1681, w_007_261);
  not1 I010_081(w_010_081, w_007_1588);
  or2  I010_082(w_010_082, w_004_1264, w_008_324);
  or2  I010_083(w_010_083, w_003_193, w_005_914);
  and2 I010_084(w_010_084, w_008_595, w_001_392);
  not1 I010_085(w_010_085, w_005_1296);
  nand2 I010_086(w_010_086, w_005_363, w_003_119);
  or2  I010_087(w_010_087, w_006_081, w_002_107);
  nand2 I010_088(w_010_088, w_009_081, w_008_501);
  or2  I010_089(w_010_089, w_009_042, w_000_1852);
  and2 I010_090(w_010_090, w_005_1118, w_002_157);
  or2  I010_091(w_010_091, w_003_137, w_005_278);
  not1 I010_092(w_010_092, w_009_056);
  or2  I010_093(w_010_093, w_004_175, w_004_260);
  and2 I010_094(w_010_094, w_007_1313, w_000_1366);
  not1 I010_095(w_010_095, w_000_1084);
  and2 I010_096(w_010_096, w_009_007, w_006_237);
  nand2 I010_097(w_010_097, w_004_051, w_005_1199);
  and2 I010_098(w_010_098, w_001_1289, w_002_149);
  nand2 I010_099(w_010_099, w_003_067, w_006_063);
  and2 I010_101(w_010_101, w_003_168, w_000_1516);
  or2  I010_102(w_010_102, w_006_245, w_002_571);
  nand2 I010_103(w_010_103, w_005_1019, w_002_200);
  not1 I010_104(w_010_104, w_009_067);
  nand2 I010_105(w_010_105, w_003_287, w_006_302);
  not1 I010_106(w_010_106, w_003_125);
  and2 I010_108(w_010_108, w_000_236, w_000_016);
  or2  I010_109(w_010_109, w_009_054, w_003_274);
  or2  I010_110(w_010_110, w_000_893, w_007_1083);
  nand2 I010_111(w_010_111, w_006_038, w_005_1461);
  or2  I010_112(w_010_112, w_001_107, w_004_576);
  and2 I010_113(w_010_113, w_005_994, w_000_230);
  not1 I010_114(w_010_114, w_000_731);
  nand2 I010_115(w_010_115, w_001_1099, w_002_424);
  or2  I010_116(w_010_116, w_008_621, w_008_718);
  nand2 I010_117(w_010_117, w_006_153, w_006_324);
  and2 I010_118(w_010_118, w_003_186, w_003_207);
  or2  I010_119(w_010_119, w_007_063, w_000_075);
  and2 I010_121(w_010_121, w_001_1388, w_005_794);
  and2 I010_122(w_010_122, w_000_406, w_003_098);
  and2 I010_123(w_010_123, w_002_026, w_005_323);
  not1 I010_124(w_010_124, w_003_082);
  not1 I010_125(w_010_125, w_007_188);
  nand2 I010_126(w_010_126, w_004_1474, w_001_307);
  and2 I010_127(w_010_127, w_006_039, w_006_217);
  and2 I010_128(w_010_128, w_007_1334, w_009_107);
  not1 I010_129(w_010_129, w_009_097);
  and2 I010_131(w_010_131, w_009_016, w_004_1204);
  not1 I010_132(w_010_132, w_001_1392);
  or2  I010_133(w_010_133, w_005_1218, w_002_384);
  not1 I010_134(w_010_134, w_008_144);
  or2  I010_135(w_010_135, w_004_1128, w_000_1310);
  nand2 I010_136(w_010_136, w_004_1484, w_007_359);
  or2  I010_138(w_010_138, w_006_034, w_001_1452);
  and2 I010_139(w_010_139, w_004_1197, w_004_359);
  nand2 I010_140(w_010_140, w_008_744, w_002_187);
  and2 I010_141(w_010_141, w_003_163, w_008_163);
  or2  I010_146(w_010_146, w_007_267, w_007_1259);
  not1 I010_147(w_010_147, w_007_1182);
  nand2 I010_149(w_010_149, w_009_003, w_002_303);
  not1 I010_150(w_010_150, w_006_247);
  nand2 I010_151(w_010_151, w_009_055, w_005_244);
  nand2 I010_153(w_010_153, w_006_081, w_006_217);
  nand2 I010_154(w_010_154, w_005_1119, w_000_534);
  not1 I010_155(w_010_155, w_000_318);
  or2  I010_156(w_010_156, w_009_001, w_001_1305);
  nand2 I010_157(w_010_157, w_007_592, w_009_009);
  nand2 I010_158(w_010_158, w_004_1053, w_008_268);
  nand2 I010_159(w_010_159, w_009_085, w_000_317);
  not1 I010_160(w_010_160, w_008_254);
  not1 I010_161(w_010_161, w_003_125);
  not1 I010_162(w_010_162, w_007_624);
  or2  I010_163(w_010_163, w_008_808, w_002_329);
  or2  I010_164(w_010_164, w_007_213, w_002_139);
  and2 I010_165(w_010_165, w_001_898, w_002_537);
  or2  I010_166(w_010_166, w_001_448, w_008_526);
  nand2 I010_167(w_010_167, w_008_188, w_009_064);
  not1 I010_168(w_010_168, w_005_1150);
  or2  I010_169(w_010_169, w_002_126, w_002_120);
  nand2 I010_170(w_010_170, w_004_232, w_006_080);
  or2  I010_171(w_010_171, w_001_1251, w_007_482);
  not1 I010_172(w_010_172, w_001_1371);
  nand2 I010_173(w_010_173, w_002_038, w_009_050);
  nand2 I010_174(w_010_174, w_007_295, w_002_214);
  or2  I010_175(w_010_175, w_007_904, w_008_807);
  not1 I010_176(w_010_176, w_000_1574);
  or2  I010_177(w_010_177, w_005_158, w_008_192);
  nand2 I010_178(w_010_178, w_009_100, w_006_043);
  or2  I010_180(w_010_180, w_002_157, w_005_268);
  not1 I010_181(w_010_181, w_004_214);
  not1 I010_184(w_010_184, w_002_048);
  nand2 I010_185(w_010_185, w_001_1446, w_006_212);
  nand2 I010_186(w_010_186, w_007_1049, w_002_511);
  not1 I010_188(w_010_188, w_004_1410);
  and2 I010_189(w_010_189, w_000_1557, w_005_322);
  or2  I010_190(w_010_190, w_007_924, w_001_1232);
  not1 I010_191(w_010_191, w_003_180);
  not1 I010_192(w_010_192, w_006_266);
  not1 I010_193(w_010_193, w_007_001);
  nand2 I010_194(w_010_194, w_008_162, w_003_255);
  or2  I010_196(w_010_196, w_008_148, w_005_977);
  nand2 I010_197(w_010_197, w_007_1450, w_003_233);
  nand2 I010_198(w_010_198, w_005_780, w_006_317);
  not1 I010_199(w_010_199, w_003_263);
  and2 I010_200(w_010_200, w_002_560, w_004_1330);
  nand2 I010_201(w_010_201, w_009_033, w_006_187);
  or2  I010_202(w_010_202, w_004_713, w_002_026);
  nand2 I010_203(w_010_203, w_008_543, w_007_887);
  or2  I010_204(w_010_204, w_000_1761, w_006_049);
  or2  I010_205(w_010_205, w_004_1054, w_001_1629);
  or2  I010_206(w_010_206, w_003_121, w_001_467);
  nand2 I010_207(w_010_207, w_008_401, w_002_383);
  or2  I010_208(w_010_208, w_000_1123, w_000_1889);
  not1 I010_210(w_010_210, w_007_141);
  nand2 I010_211(w_010_211, w_003_182, w_004_079);
  and2 I010_212(w_010_212, w_007_085, w_009_030);
  not1 I010_213(w_010_213, w_000_178);
  not1 I010_214(w_010_214, w_000_1796);
  not1 I010_215(w_010_215, w_007_634);
  and2 I010_216(w_010_216, w_000_536, w_007_779);
  not1 I010_217(w_010_217, w_009_011);
  or2  I010_219(w_010_219, w_004_1456, w_003_114);
  nand2 I010_220(w_010_220, w_002_441, w_004_984);
  or2  I010_221(w_010_221, w_004_602, w_006_080);
  or2  I010_222(w_010_222, w_005_786, w_007_314);
  nand2 I010_223(w_010_223, w_004_717, w_007_270);
  or2  I010_224(w_010_224, w_003_083, w_001_285);
  and2 I010_225(w_010_225, w_005_812, w_002_200);
  not1 I010_226(w_010_226, w_006_018);
  not1 I010_227(w_010_227, w_002_510);
  nand2 I010_228(w_010_228, w_008_653, w_007_318);
  not1 I010_229(w_010_229, w_003_177);
  nand2 I010_230(w_010_230, w_003_172, w_004_1850);
  or2  I010_231(w_010_231, w_008_066, w_002_449);
  and2 I010_233(w_010_233, w_000_1850, w_000_614);
  and2 I010_234(w_010_234, w_004_664, w_004_452);
  or2  I010_235(w_010_235, w_001_1122, w_009_054);
  nand2 I010_236(w_010_236, w_007_979, w_001_941);
  not1 I010_237(w_010_237, w_001_1581);
  or2  I010_238(w_010_238, w_005_624, w_000_495);
  and2 I010_239(w_010_239, w_002_505, w_000_722);
  not1 I010_241(w_010_241, w_004_705);
  not1 I010_242(w_010_242, w_008_374);
  and2 I010_244(w_010_244, w_000_1253, w_000_1791);
  not1 I010_245(w_010_245, w_004_044);
  nand2 I010_246(w_010_246, w_009_108, w_005_015);
  nand2 I010_247(w_010_247, w_001_512, w_007_811);
  nand2 I010_248(w_010_248, w_009_019, w_007_159);
  and2 I010_250(w_010_250, w_000_117, w_006_008);
  not1 I010_251(w_010_251, w_008_318);
  and2 I010_252(w_010_252, w_002_392, w_009_082);
  and2 I010_253(w_010_253, w_004_1244, w_009_042);
  and2 I010_254(w_010_254, w_008_661, w_005_1079);
  or2  I010_256(w_010_256, w_006_122, w_005_966);
  not1 I010_259(w_010_259, w_003_299);
  not1 I010_260(w_010_260, w_005_789);
  nand2 I010_261(w_010_261, w_005_1450, w_000_1647);
  nand2 I010_262(w_010_262, w_007_862, w_004_1769);
  nand2 I010_263(w_010_263, w_002_109, w_008_273);
  nand2 I010_264(w_010_264, w_001_1144, w_004_1415);
  or2  I010_265(w_010_265, w_008_114, w_009_082);
  not1 I010_266(w_010_266, w_004_1053);
  or2  I010_267(w_010_267, w_001_152, w_004_1069);
  or2  I010_268(w_010_268, w_006_028, w_004_476);
  not1 I010_269(w_010_269, w_008_245);
  or2  I010_270(w_010_270, w_000_136, w_007_740);
  nand2 I010_271(w_010_271, w_000_236, w_004_278);
  not1 I010_272(w_010_272, w_004_122);
  or2  I010_273(w_010_273, w_008_731, w_009_090);
  or2  I010_274(w_010_274, w_003_188, w_003_052);
  or2  I010_275(w_010_275, w_002_494, w_008_228);
  not1 I010_276(w_010_276, w_008_825);
  nand2 I010_277(w_010_277, w_001_961, w_006_159);
  or2  I010_278(w_010_278, w_006_052, w_009_104);
  not1 I010_279(w_010_279, w_005_1346);
  nand2 I010_280(w_010_280, w_003_015, w_000_1717);
  and2 I010_281(w_010_281, w_003_258, w_008_802);
  nand2 I010_282(w_010_282, w_002_161, w_001_610);
  or2  I010_283(w_010_283, w_002_005, w_000_153);
  and2 I010_284(w_010_284, w_008_831, w_003_095);
  and2 I010_285(w_010_285, w_002_037, w_000_877);
  not1 I010_286(w_010_286, w_009_073);
  or2  I010_287(w_010_287, w_002_108, w_009_081);
  and2 I010_288(w_010_288, w_009_069, w_004_581);
  not1 I010_290(w_010_290, w_006_048);
  nand2 I010_291(w_010_291, w_005_1473, w_004_042);
  or2  I010_292(w_010_292, w_009_001, w_000_1076);
  nand2 I010_293(w_010_293, w_001_019, w_000_563);
  and2 I010_294(w_010_294, w_002_033, w_004_1453);
  not1 I010_295(w_010_295, w_008_035);
  and2 I010_297(w_010_297, w_007_1261, w_009_098);
  and2 I010_298(w_010_298, w_006_075, w_000_1740);
  and2 I010_299(w_010_299, w_009_077, w_006_104);
  or2  I010_300(w_010_300, w_000_1197, w_001_1045);
  and2 I010_302(w_010_302, w_006_124, w_009_072);
  not1 I010_303(w_010_303, w_001_1642);
  nand2 I010_304(w_010_304, w_002_316, w_003_040);
  nand2 I010_305(w_010_305, w_004_420, w_009_023);
  not1 I010_306(w_010_306, w_008_326);
  nand2 I010_307(w_010_307, w_000_741, w_008_015);
  not1 I010_308(w_010_308, w_006_282);
  and2 I010_309(w_010_309, w_005_446, w_009_001);
  or2  I010_310(w_010_310, w_003_287, w_009_021);
  nand2 I010_311(w_010_311, w_003_273, w_000_1524);
  and2 I010_312(w_010_312, w_004_296, w_008_470);
  or2  I010_315(w_010_315, w_006_067, w_009_039);
  not1 I010_316(w_010_316, w_008_199);
  nand2 I010_317(w_010_317, w_004_663, w_002_053);
  not1 I010_318(w_010_318, w_006_139);
  nand2 I010_320(w_010_320, w_009_015, w_005_023);
  and2 I010_321(w_010_321, w_005_777, w_004_839);
  not1 I010_322(w_010_322, w_002_070);
  and2 I010_323(w_010_323, w_005_097, w_004_1179);
  and2 I010_324(w_010_324, w_008_195, w_008_422);
  or2  I010_325(w_010_325, w_004_1601, w_008_628);
  and2 I010_326(w_010_326, w_000_1609, w_006_175);
  and2 I010_327(w_010_327, w_003_222, w_008_544);
  and2 I010_328(w_010_328, w_003_280, w_006_323);
  not1 I010_329(w_010_329, w_002_041);
  nand2 I010_330(w_010_330, w_007_1002, w_007_1047);
  or2  I010_331(w_010_331, w_005_146, w_005_1292);
  not1 I010_332(w_010_332, w_005_272);
  nand2 I010_333(w_010_333, w_005_206, w_001_057);
  or2  I010_334(w_010_334, w_004_641, w_006_047);
  not1 I010_336(w_010_336, w_004_1399);
  or2  I010_337(w_010_337, w_003_114, w_004_1553);
  nand2 I010_338(w_010_338, w_001_1374, w_000_1323);
  or2  I010_339(w_010_339, w_008_218, w_004_1643);
  and2 I010_342(w_010_342, w_009_090, w_008_691);
  not1 I010_343(w_010_343, w_005_034);
  and2 I010_344(w_010_344, w_001_1262, w_005_263);
  or2  I010_345(w_010_345, w_006_210, w_000_1654);
  not1 I010_346(w_010_346, w_004_1649);
  and2 I010_347(w_010_347, w_001_1392, w_007_774);
  and2 I010_348(w_010_348, w_002_263, w_005_178);
  not1 I010_350(w_010_350, w_006_064);
  not1 I010_351(w_010_351, w_007_055);
  not1 I010_352(w_010_352, w_000_1020);
  and2 I010_353(w_010_353, w_009_054, w_008_460);
  and2 I010_354(w_010_354, w_007_1393, w_007_931);
  and2 I010_355(w_010_355, w_001_707, w_002_085);
  or2  I010_356(w_010_356, w_002_361, w_002_521);
  or2  I010_357(w_010_357, w_007_393, w_001_751);
  and2 I010_358(w_010_358, w_009_110, w_008_861);
  not1 I010_359(w_010_359, w_000_300);
  and2 I010_360(w_010_360, w_008_248, w_008_755);
  nand2 I010_363(w_010_363, w_001_1023, w_007_1486);
  nand2 I010_365(w_010_365, w_003_240, w_001_134);
  nand2 I010_366(w_010_366, w_003_147, w_007_531);
  or2  I010_367(w_010_367, w_006_263, w_008_073);
  and2 I010_369(w_010_369, w_001_300, w_000_1890);
  or2  I010_370(w_010_370, w_007_206, w_004_134);
  or2  I010_371(w_010_371, w_008_727, w_007_691);
  and2 I010_372(w_010_372, w_000_1177, w_007_746);
  and2 I010_373(w_010_373, w_007_005, w_001_073);
  and2 I010_374(w_010_374, w_000_188, w_008_082);
  nand2 I010_375(w_010_375, w_007_079, w_001_539);
  nand2 I010_376(w_010_376, w_007_318, w_009_077);
  and2 I010_377(w_010_377, w_003_071, w_006_116);
  not1 I010_378(w_010_378, w_001_1274);
  nand2 I010_379(w_010_379, w_008_020, w_006_071);
  not1 I010_380(w_010_380, w_007_1562);
  not1 I010_381(w_010_381, w_007_127);
  or2  I010_382(w_010_382, w_002_214, w_008_500);
  not1 I010_384(w_010_384, w_007_1010);
  or2  I010_385(w_010_385, w_008_541, w_001_932);
  nand2 I010_386(w_010_386, w_006_168, w_008_046);
  and2 I010_387(w_010_387, w_005_103, w_009_046);
  or2  I010_388(w_010_388, w_009_005, w_002_183);
  and2 I010_391(w_010_391, w_009_011, w_005_671);
  nand2 I010_392(w_010_392, w_002_427, w_001_722);
  and2 I010_394(w_010_394, w_007_1374, w_009_089);
  and2 I010_397(w_010_397, w_009_108, w_005_574);
  nand2 I010_398(w_010_398, w_004_148, w_000_186);
  nand2 I010_399(w_010_399, w_008_856, w_001_176);
  not1 I010_400(w_010_400, w_009_055);
  and2 I010_401(w_010_401, w_008_511, w_007_1022);
  nand2 I010_402(w_010_402, w_003_088, w_003_154);
  and2 I010_403(w_010_403, w_005_025, w_004_756);
  nand2 I010_405(w_010_405, w_003_151, w_004_1033);
  or2  I010_406(w_010_406, w_005_1561, w_001_274);
  and2 I010_408(w_010_408, w_003_256, w_008_753);
  nand2 I010_411(w_010_411, w_000_381, w_006_065);
  and2 I010_413(w_010_413, w_001_271, w_007_221);
  or2  I010_414(w_010_414, w_001_026, w_005_197);
  nand2 I010_415(w_010_415, w_003_215, w_007_066);
  nand2 I010_416(w_010_416, w_007_1142, w_006_306);
  not1 I010_417(w_010_417, w_001_1516);
  and2 I010_419(w_010_419, w_005_796, w_003_078);
  nand2 I010_420(w_010_420, w_002_015, w_006_135);
  and2 I010_421(w_009_122, w_007_808, w_009_113);
  or2  I011_000(w_011_000, w_009_088, w_010_277);
  not1 I011_001(w_011_001, w_009_071);
  nand2 I011_002(w_011_002, w_000_1739, w_003_109);
  not1 I011_003(w_011_003, w_005_752);
  nand2 I011_004(w_011_004, w_007_279, w_010_102);
  and2 I011_005(w_011_005, w_007_064, w_005_1043);
  not1 I011_006(w_011_006, w_002_077);
  or2  I011_007(w_011_007, w_002_220, w_001_1147);
  and2 I011_009(w_011_009, w_005_1653, w_009_063);
  nand2 I011_010(w_011_010, w_003_223, w_000_1089);
  nand2 I011_011(w_011_011, w_010_280, w_004_1008);
  not1 I011_014(w_011_014, w_001_101);
  nand2 I011_015(w_011_015, w_007_057, w_004_1868);
  not1 I011_016(w_011_016, w_002_346);
  not1 I011_018(w_011_018, w_006_145);
  not1 I011_019(w_011_019, w_000_837);
  and2 I011_020(w_011_020, w_008_193, w_003_226);
  not1 I011_021(w_011_021, w_001_022);
  and2 I011_022(w_011_022, w_004_916, w_002_545);
  and2 I011_026(w_011_026, w_008_819, w_002_528);
  or2  I011_028(w_011_028, w_007_1184, w_004_396);
  and2 I011_031(w_011_031, w_005_856, w_003_219);
  not1 I011_033(w_011_033, w_000_1257);
  or2  I011_034(w_011_034, w_006_068, w_005_1298);
  and2 I011_035(w_011_035, w_009_046, w_001_785);
  not1 I011_036(w_011_036, w_007_755);
  not1 I011_037(w_011_037, w_007_875);
  not1 I011_038(w_011_038, w_010_091);
  and2 I011_039(w_011_039, w_005_260, w_007_294);
  and2 I011_040(w_011_040, w_005_294, w_010_117);
  or2  I011_041(w_011_041, w_007_1530, w_009_083);
  or2  I011_042(w_011_042, w_008_136, w_000_1893);
  or2  I011_043(w_011_043, w_004_1841, w_001_086);
  nand2 I011_044(w_011_044, w_009_081, w_010_358);
  not1 I011_046(w_011_046, w_002_211);
  or2  I011_051(w_011_051, w_009_000, w_001_038);
  not1 I011_052(w_011_052, w_005_1478);
  and2 I011_056(w_011_056, w_008_633, w_008_734);
  not1 I011_057(w_011_057, w_004_374);
  not1 I011_058(w_011_058, w_009_027);
  and2 I011_060(w_011_060, w_006_054, w_007_1598);
  and2 I011_062(w_011_062, w_005_559, w_007_104);
  nand2 I011_063(w_011_063, w_004_1602, w_000_1844);
  or2  I011_064(w_011_064, w_002_570, w_007_307);
  or2  I011_065(w_011_065, w_009_099, w_001_306);
  nand2 I011_067(w_011_067, w_003_111, w_007_703);
  or2  I011_068(w_011_068, w_004_425, w_007_1026);
  nand2 I011_070(w_011_070, w_004_587, w_008_156);
  not1 I011_071(w_011_071, w_010_327);
  not1 I011_072(w_011_072, w_009_035);
  nand2 I011_073(w_011_073, w_010_328, w_010_124);
  nand2 I011_074(w_011_074, w_002_256, w_008_404);
  and2 I011_076(w_011_076, w_008_696, w_008_236);
  and2 I011_077(w_011_077, w_010_333, w_000_1869);
  not1 I011_079(w_011_079, w_004_1832);
  not1 I011_080(w_011_080, w_001_377);
  not1 I011_081(w_011_081, w_003_025);
  nand2 I011_085(w_011_085, w_000_1894, w_007_1153);
  and2 I011_086(w_011_086, w_009_008, w_009_052);
  and2 I011_088(w_011_088, w_000_1895, w_005_251);
  not1 I011_091(w_011_091, w_002_483);
  nand2 I011_092(w_011_092, w_003_194, w_009_020);
  or2  I011_093(w_011_093, w_001_340, w_005_087);
  nand2 I011_094(w_011_094, w_005_1421, w_010_031);
  and2 I011_097(w_011_097, w_009_053, w_000_1328);
  nand2 I011_098(w_011_098, w_000_999, w_004_1430);
  nand2 I011_100(w_011_100, w_002_070, w_009_105);
  and2 I011_101(w_011_101, w_009_055, w_010_324);
  or2  I011_102(w_011_102, w_003_184, w_010_085);
  nand2 I011_103(w_011_103, w_009_016, w_003_073);
  and2 I011_104(w_011_104, w_006_315, w_002_086);
  or2  I011_105(w_011_105, w_006_075, w_010_077);
  or2  I011_107(w_011_107, w_003_125, w_006_196);
  and2 I011_108(w_011_108, w_005_229, w_000_1033);
  or2  I011_109(w_011_109, w_010_276, w_002_253);
  or2  I011_111(w_011_111, w_008_638, w_010_366);
  or2  I011_112(w_011_112, w_008_035, w_004_1096);
  or2  I011_114(w_011_114, w_008_544, w_000_1147);
  or2  I011_115(w_011_115, w_003_208, w_000_347);
  and2 I011_117(w_011_117, w_001_570, w_005_653);
  and2 I011_118(w_011_118, w_002_079, w_007_742);
  or2  I011_119(w_011_119, w_010_191, w_000_1241);
  and2 I011_120(w_011_120, w_000_1763, w_009_096);
  nand2 I011_122(w_011_122, w_010_234, w_005_1308);
  or2  I011_123(w_011_123, w_010_046, w_003_156);
  nand2 I011_125(w_011_125, w_004_222, w_003_144);
  and2 I011_126(w_011_126, w_006_303, w_009_004);
  nand2 I011_127(w_011_127, w_006_252, w_009_043);
  nand2 I011_128(w_011_128, w_003_144, w_008_181);
  and2 I011_129(w_011_129, w_005_341, w_010_042);
  and2 I011_132(w_011_132, w_005_257, w_004_1149);
  or2  I011_133(w_011_133, w_001_1387, w_010_228);
  and2 I011_135(w_011_135, w_002_349, w_006_323);
  nand2 I011_136(w_011_136, w_001_1602, w_002_154);
  not1 I011_137(w_011_137, w_001_274);
  or2  I011_140(w_011_140, w_003_117, w_004_029);
  nand2 I011_141(w_011_141, w_001_596, w_000_160);
  and2 I011_142(w_011_142, w_003_201, w_008_200);
  not1 I011_143(w_011_143, w_007_997);
  or2  I011_144(w_011_144, w_005_930, w_007_891);
  not1 I011_147(w_011_147, w_001_1427);
  or2  I011_148(w_011_148, w_002_023, w_002_323);
  not1 I011_150(w_011_150, w_005_729);
  nand2 I011_151(w_011_151, w_008_794, w_006_311);
  nand2 I011_152(w_011_152, w_001_226, w_000_198);
  or2  I011_154(w_011_154, w_002_413, w_006_218);
  or2  I011_155(w_011_155, w_009_081, w_006_059);
  and2 I011_157(w_011_157, w_001_1314, w_000_192);
  and2 I011_159(w_011_159, w_001_081, w_006_090);
  and2 I011_160(w_011_160, w_008_501, w_008_013);
  and2 I011_161(w_011_161, w_000_1832, w_009_087);
  or2  I011_163(w_011_163, w_009_063, w_006_111);
  nand2 I011_164(w_011_164, w_005_1394, w_004_206);
  or2  I011_166(w_011_166, w_003_229, w_005_654);
  or2  I011_169(w_011_169, w_004_046, w_006_275);
  not1 I011_170(w_011_170, w_005_1548);
  and2 I011_171(w_011_171, w_009_106, w_001_1517);
  or2  I011_172(w_011_172, w_009_010, w_006_188);
  and2 I011_173(w_011_173, w_000_1186, w_007_186);
  nand2 I011_176(w_011_176, w_008_144, w_004_1656);
  and2 I011_177(w_011_177, w_007_1204, w_006_146);
  not1 I011_181(w_011_181, w_005_1542);
  nand2 I011_182(w_011_182, w_010_268, w_003_090);
  nand2 I011_184(w_011_184, w_006_100, w_000_239);
  not1 I011_185(w_011_185, w_005_1584);
  nand2 I011_188(w_011_188, w_010_300, w_001_1308);
  not1 I011_189(w_011_189, w_009_093);
  not1 I011_190(w_011_190, w_003_079);
  not1 I011_193(w_011_193, w_003_059);
  and2 I011_194(w_011_194, w_000_1583, w_005_952);
  or2  I011_196(w_011_196, w_001_630, w_000_1505);
  not1 I011_197(w_011_197, w_000_1584);
  or2  I011_199(w_011_199, w_001_367, w_004_770);
  and2 I011_201(w_011_201, w_005_1672, w_000_729);
  nand2 I011_203(w_011_203, w_006_307, w_003_300);
  nand2 I011_204(w_011_204, w_004_303, w_001_1196);
  and2 I011_205(w_011_205, w_007_304, w_007_441);
  not1 I011_206(w_011_206, w_010_344);
  or2  I011_208(w_011_208, w_010_112, w_000_1882);
  nand2 I011_209(w_011_209, w_006_339, w_006_322);
  not1 I011_210(w_011_210, w_007_318);
  nand2 I011_213(w_011_213, w_003_006, w_005_114);
  nand2 I011_215(w_011_215, w_009_079, w_007_366);
  not1 I011_216(w_011_216, w_003_096);
  or2  I011_217(w_011_217, w_010_244, w_000_1741);
  nand2 I011_219(w_011_219, w_002_084, w_003_186);
  not1 I011_221(w_011_221, w_008_195);
  nand2 I011_224(w_011_224, w_007_084, w_009_057);
  nand2 I011_225(w_011_225, w_007_149, w_002_434);
  and2 I011_227(w_011_227, w_002_459, w_002_064);
  nand2 I011_228(w_011_228, w_006_026, w_010_252);
  or2  I011_229(w_011_229, w_006_099, w_000_019);
  or2  I011_230(w_011_230, w_002_471, w_004_1027);
  or2  I011_232(w_011_232, w_007_1583, w_007_1233);
  and2 I011_233(w_011_233, w_006_175, w_000_091);
  not1 I011_235(w_011_235, w_006_134);
  and2 I011_242(w_011_242, w_001_143, w_004_1186);
  nand2 I011_243(w_011_243, w_009_012, w_009_015);
  or2  I011_244(w_011_244, w_004_1248, w_008_563);
  nand2 I011_246(w_011_246, w_002_482, w_000_1506);
  or2  I011_247(w_011_247, w_006_094, w_002_200);
  not1 I011_250(w_011_250, w_003_184);
  and2 I011_256(w_011_256, w_000_1640, w_005_1125);
  and2 I011_257(w_011_257, w_000_1196, w_008_279);
  not1 I011_258(w_011_258, w_007_916);
  and2 I011_260(w_011_260, w_006_069, w_002_433);
  not1 I011_262(w_011_262, w_004_375);
  and2 I011_263(w_011_263, w_009_079, w_010_018);
  nand2 I011_265(w_011_265, w_002_525, w_003_225);
  nand2 I011_267(w_011_267, w_008_540, w_006_145);
  and2 I011_272(w_011_272, w_009_064, w_010_132);
  and2 I011_273(w_011_273, w_000_1072, w_002_213);
  or2  I011_283(w_011_283, w_003_123, w_006_234);
  and2 I011_286(w_011_286, w_000_1896, w_010_173);
  and2 I011_290(w_011_290, w_006_249, w_002_376);
  not1 I011_293(w_011_293, w_008_018);
  and2 I011_295(w_011_295, w_009_000, w_005_580);
  nand2 I011_297(w_011_297, w_006_001, w_004_301);
  or2  I011_298(w_011_298, w_008_437, w_002_565);
  not1 I011_303(w_011_303, w_002_579);
  not1 I011_304(w_011_304, w_006_245);
  and2 I011_307(w_011_307, w_004_1855, w_003_060);
  or2  I011_309(w_011_309, w_002_447, w_003_200);
  nand2 I011_313(w_011_313, w_002_564, w_007_1263);
  and2 I011_314(w_011_314, w_010_315, w_000_1474);
  not1 I011_315(w_011_315, w_000_1635);
  nand2 I011_316(w_011_316, w_000_1028, w_005_097);
  and2 I011_318(w_011_318, w_003_140, w_000_1655);
  or2  I011_320(w_011_320, w_007_222, w_002_585);
  not1 I011_323(w_011_323, w_005_1224);
  not1 I011_324(w_011_324, w_003_084);
  not1 I011_325(w_011_325, w_004_590);
  not1 I011_327(w_011_327, w_001_281);
  or2  I011_328(w_011_328, w_006_252, w_007_1219);
  not1 I011_332(w_011_332, w_002_130);
  not1 I011_333(w_011_333, w_001_1142);
  and2 I011_334(w_011_334, w_002_231, w_010_266);
  nand2 I011_338(w_011_338, w_004_1619, w_002_081);
  not1 I011_339(w_011_339, w_008_217);
  and2 I011_344(w_011_344, w_007_1197, w_000_1889);
  and2 I011_345(w_011_345, w_000_565, w_003_223);
  nand2 I011_347(w_011_347, w_005_1447, w_007_214);
  and2 I011_350(w_011_350, w_007_307, w_005_159);
  or2  I011_353(w_011_353, w_008_489, w_004_1390);
  or2  I011_354(w_011_354, w_000_1228, w_001_337);
  and2 I011_357(w_011_357, w_003_267, w_008_381);
  and2 I011_360(w_011_360, w_006_057, w_004_181);
  not1 I011_361(w_011_361, w_003_153);
  nand2 I011_363(w_011_363, w_001_615, w_008_006);
  not1 I011_365(w_011_365, w_009_098);
  not1 I011_368(w_011_368, w_000_539);
  and2 I011_369(w_011_369, w_009_023, w_004_1861);
  not1 I011_371(w_011_371, w_002_506);
  or2  I011_372(w_011_372, w_008_241, w_006_336);
  nand2 I011_374(w_011_374, w_006_092, w_008_122);
  nand2 I011_378(w_011_378, w_009_026, w_002_340);
  and2 I011_381(w_011_381, w_005_209, w_008_197);
  not1 I011_383(w_011_383, w_005_605);
  nand2 I011_384(w_011_384, w_004_220, w_003_126);
  nand2 I011_386(w_011_386, w_008_743, w_004_1200);
  and2 I011_388(w_011_388, w_008_103, w_009_080);
  or2  I011_389(w_011_389, w_003_185, w_002_045);
  nand2 I011_390(w_011_390, w_007_790, w_000_1672);
  or2  I011_391(w_011_391, w_008_798, w_005_047);
  not1 I011_394(w_011_394, w_000_1111);
  not1 I011_395(w_011_395, w_006_256);
  nand2 I011_398(w_011_398, w_007_951, w_010_367);
  nand2 I011_401(w_011_401, w_007_1360, w_003_163);
  and2 I011_402(w_011_402, w_006_182, w_001_1125);
  and2 I011_403(w_011_403, w_000_398, w_008_765);
  nand2 I011_404(w_011_404, w_004_929, w_004_1888);
  and2 I011_405(w_011_405, w_001_1449, w_009_096);
  and2 I011_406(w_011_406, w_010_305, w_002_093);
  not1 I011_407(w_011_407, w_000_1713);
  and2 I011_411(w_011_411, w_009_062, w_009_014);
  and2 I011_412(w_011_412, w_008_806, w_005_046);
  not1 I011_414(w_011_414, w_010_157);
  nand2 I011_417(w_011_417, w_002_001, w_006_085);
  not1 I011_419(w_011_419, w_010_202);
  and2 I011_420(w_011_420, w_006_066, w_001_895);
  nand2 I011_424(w_011_424, w_001_593, w_009_035);
  nand2 I011_425(w_011_425, w_000_502, w_001_475);
  and2 I011_426(w_011_426, w_000_577, w_007_568);
  or2  I011_428(w_011_428, w_009_035, w_005_1239);
  nand2 I011_429(w_011_429, w_008_164, w_010_388);
  nand2 I011_432(w_011_432, w_000_441, w_010_018);
  not1 I011_433(w_011_433, w_004_938);
  and2 I011_435(w_011_435, w_000_1413, w_003_049);
  or2  I011_436(w_011_436, w_010_324, w_003_274);
  or2  I011_439(w_011_439, w_000_006, w_007_636);
  and2 I011_440(w_011_440, w_009_023, w_003_089);
  not1 I011_441(w_011_441, w_000_1046);
  and2 I011_444(w_011_444, w_006_093, w_010_227);
  nand2 I011_445(w_011_445, w_010_108, w_007_293);
  not1 I011_449(w_011_449, w_007_272);
  not1 I011_453(w_011_453, w_009_036);
  not1 I011_454(w_011_454, w_003_273);
  or2  I011_455(w_011_455, w_004_778, w_009_107);
  and2 I011_459(w_011_459, w_010_229, w_010_299);
  not1 I011_460(w_011_460, w_008_209);
  or2  I011_461(w_011_461, w_000_1812, w_002_011);
  nand2 I011_463(w_011_463, w_006_290, w_009_048);
  nand2 I011_464(w_011_464, w_000_740, w_009_093);
  nand2 I011_465(w_011_465, w_007_639, w_001_233);
  nand2 I011_466(w_011_466, w_001_568, w_006_196);
  and2 I011_469(w_011_469, w_002_199, w_005_039);
  not1 I011_470(w_011_470, w_001_609);
  not1 I011_471(w_011_471, w_000_622);
  or2  I011_474(w_011_474, w_009_012, w_008_282);
  not1 I011_475(w_011_475, w_008_360);
  or2  I011_479(w_011_479, w_002_467, w_009_075);
  not1 I011_480(w_011_480, w_006_260);
  not1 I011_482(w_011_482, w_008_685);
  nand2 I011_483(w_011_483, w_010_199, w_000_1659);
  not1 I011_485(w_011_485, w_004_373);
  and2 I011_489(w_011_489, w_000_203, w_000_633);
  not1 I011_490(w_011_490, w_009_068);
  nand2 I011_491(w_011_491, w_010_245, w_004_1054);
  not1 I011_492(w_011_492, w_006_161);
  or2  I011_493(w_011_493, w_001_818, w_002_463);
  not1 I011_496(w_011_496, w_003_073);
  not1 I011_498(w_011_498, w_002_148);
  nand2 I011_501(w_011_501, w_001_1074, w_004_585);
  not1 I011_503(w_011_503, w_009_008);
  or2  I011_504(w_011_504, w_004_1597, w_003_070);
  or2  I011_508(w_011_508, w_005_1560, w_004_714);
  or2  I011_509(w_011_509, w_005_530, w_006_148);
  and2 I011_510(w_011_510, w_004_501, w_009_068);
  not1 I011_512(w_011_512, w_003_293);
  and2 I011_515(w_011_515, w_009_061, w_005_1137);
  or2  I011_517(w_011_517, w_000_393, w_009_107);
  not1 I011_522(w_011_522, w_007_740);
  and2 I011_523(w_011_523, w_007_189, w_002_155);
  or2  I011_525(w_011_525, w_000_1782, w_004_1206);
  nand2 I011_527(w_011_527, w_009_094, w_003_027);
  not1 I011_532(w_011_532, w_007_144);
  and2 I011_533(w_011_533, w_009_019, w_007_000);
  not1 I011_534(w_011_534, w_008_612);
  nand2 I011_536(w_011_536, w_010_031, w_005_494);
  not1 I011_538(w_011_538, w_005_228);
  and2 I011_539(w_011_539, w_004_1911, w_010_392);
  or2  I011_541(w_011_541, w_002_559, w_004_597);
  or2  I011_542(w_011_542, w_002_163, w_004_909);
  or2  I011_543(w_011_543, w_007_131, w_000_447);
  or2  I011_546(w_011_546, w_004_064, w_010_190);
  not1 I011_547(w_011_547, w_007_1377);
  nand2 I011_548(w_011_548, w_008_206, w_002_471);
  nand2 I011_550(w_011_550, w_004_112, w_009_081);
  or2  I011_551(w_011_551, w_005_095, w_003_097);
  or2  I011_552(w_011_552, w_000_1107, w_001_1384);
  and2 I011_553(w_011_553, w_005_1449, w_008_100);
  and2 I011_557(w_011_557, w_003_009, w_003_293);
  or2  I011_559(w_011_559, w_002_574, w_002_089);
  nand2 I011_560(w_011_560, w_000_865, w_005_1159);
  and2 I011_565(w_011_565, w_004_123, w_000_392);
  or2  I011_568(w_011_568, w_009_059, w_001_678);
  nand2 I011_572(w_011_572, w_000_1149, w_005_038);
  and2 I011_573(w_011_573, w_010_201, w_009_034);
  and2 I011_574(w_011_574, w_010_354, w_010_318);
  nand2 I011_575(w_011_575, w_009_005, w_004_082);
  or2  I011_576(w_011_576, w_007_613, w_003_052);
  or2  I011_578(w_011_578, w_003_108, w_006_246);
  not1 I011_579(w_011_579, w_004_331);
  and2 I011_580(w_011_580, w_002_555, w_007_136);
  nand2 I011_582(w_011_582, w_002_577, w_000_1504);
  and2 I011_583(w_011_583, w_001_1188, w_005_053);
  and2 I011_584(w_011_584, w_001_106, w_003_006);
  and2 I011_586(w_011_586, w_002_181, w_009_079);
  nand2 I011_587(w_011_587, w_003_056, w_007_223);
  or2  I011_588(w_011_588, w_007_1551, w_001_1098);
  nand2 I011_589(w_011_589, w_000_895, w_005_1190);
  not1 I011_592(w_011_592, w_001_973);
  and2 I011_594(w_011_594, w_010_284, w_003_166);
  nand2 I011_596(w_011_596, w_004_588, w_010_311);
  and2 I011_597(w_011_597, w_006_029, w_009_073);
  or2  I011_598(w_011_598, w_003_129, w_009_004);
  or2  I011_610(w_011_610, w_007_1137, w_006_065);
  or2  I011_611(w_011_611, w_009_011, w_006_022);
  not1 I011_613(w_011_613, w_002_293);
  nand2 I011_617(w_011_617, w_010_167, w_004_836);
  and2 I011_619(w_011_619, w_004_912, w_005_1112);
  not1 I011_620(w_011_620, w_008_351);
  and2 I011_622(w_011_622, w_005_1116, w_000_730);
  and2 I011_623(w_011_623, w_010_099, w_009_031);
  not1 I011_624(w_011_624, w_008_346);
  or2  I011_626(w_011_626, w_003_226, w_007_781);
  or2  I011_628(w_011_628, w_005_333, w_007_1089);
  or2  I011_631(w_011_631, w_009_028, w_002_286);
  and2 I011_633(w_011_633, w_001_248, w_009_031);
  not1 I011_635(w_011_635, w_008_393);
  and2 I011_638(w_011_638, w_000_1877, w_007_251);
  nand2 I011_639(w_011_639, w_003_063, w_000_1789);
  nand2 I011_640(w_011_640, w_009_028, w_003_125);
  or2  I011_642(w_011_642, w_008_473, w_000_1156);
  nand2 I011_643(w_011_643, w_010_262, w_003_048);
  and2 I011_645(w_011_645, w_002_372, w_010_398);
  not1 I011_648(w_011_648, w_002_182);
  and2 I011_650(w_011_650, w_001_626, w_003_029);
  not1 I011_652(w_011_652, w_010_168);
  and2 I011_653(w_011_653, w_003_120, w_000_169);
  nand2 I011_654(w_011_654, w_009_000, w_008_720);
  nand2 I011_659(w_011_659, w_008_034, w_005_578);
  not1 I011_660(w_011_660, w_008_793);
  and2 I011_665(w_011_665, w_001_1514, w_004_604);
  not1 I011_666(w_011_666, w_001_990);
  and2 I011_667(w_011_667, w_007_200, w_004_1259);
  and2 I011_669(w_011_669, w_007_289, w_010_408);
  nand2 I011_670(w_011_670, w_010_151, w_010_005);
  not1 I011_674(w_011_674, w_010_227);
  and2 I011_676(w_011_676, w_010_027, w_008_732);
  not1 I011_677(w_011_677, w_005_1011);
  and2 I011_678(w_011_678, w_009_104, w_005_1447);
  not1 I011_679(w_011_679, w_007_1129);
  not1 I011_680(w_011_680, w_003_286);
  not1 I011_685(w_011_685, w_007_935);
  or2  I011_687(w_011_687, w_004_584, w_007_411);
  not1 I011_688(w_011_688, w_001_202);
  nand2 I011_691(w_011_691, w_005_1237, w_002_344);
  nand2 I011_692(w_011_692, w_009_035, w_000_1251);
  nand2 I011_694(w_011_694, w_008_128, w_005_096);
  nand2 I011_695(w_011_695, w_006_262, w_005_253);
  nand2 I011_696(w_011_696, w_004_545, w_001_1665);
  not1 I011_698(w_011_698, w_005_1330);
  not1 I011_699(w_011_699, w_003_262);
  not1 I011_700(w_011_700, w_008_680);
  or2  I011_702(w_011_702, w_002_085, w_003_100);
  and2 I011_703(w_011_703, w_007_1551, w_006_015);
  not1 I011_704(w_011_704, w_010_347);
  and2 I011_705(w_011_705, w_006_196, w_004_625);
  and2 I011_706(w_011_706, w_004_1655, w_001_1143);
  not1 I011_707(w_011_707, w_009_032);
  not1 I011_708(w_011_708, w_010_063);
  or2  I011_711(w_011_711, w_001_1096, w_003_097);
  nand2 I011_715(w_011_715, w_010_009, w_005_1239);
  nand2 I011_716(w_011_716, w_005_1669, w_002_252);
  or2  I011_718(w_011_718, w_005_1569, w_010_272);
  not1 I011_721(w_011_721, w_006_203);
  not1 I011_725(w_011_725, w_006_216);
  not1 I011_727(w_011_727, w_006_089);
  or2  I011_731(w_011_731, w_010_122, w_000_1535);
  nand2 I011_733(w_011_733, w_007_732, w_009_060);
  nand2 I011_734(w_011_734, w_005_170, w_002_064);
  not1 I011_735(w_011_735, w_009_122);
  not1 I011_738(w_011_738, w_010_086);
  or2  I011_739(w_011_739, w_009_018, w_007_088);
  and2 I011_741(w_011_741, w_007_322, w_009_056);
  and2 I011_742(w_011_742, w_004_001, w_009_003);
  or2  I011_743(w_011_743, w_009_047, w_000_671);
  not1 I011_749(w_011_749, w_001_017);
  or2  I011_751(w_011_751, w_007_443, w_002_126);
  nand2 I011_752(w_011_752, w_000_781, w_006_099);
  not1 I011_753(w_011_753, w_005_1211);
  nand2 I011_755(w_011_755, w_000_380, w_007_1599);
  or2  I011_757(w_011_757, w_008_538, w_009_012);
  or2  I011_758(w_011_758, w_006_207, w_002_398);
  not1 I011_762(w_011_762, w_008_454);
  and2 I011_763(w_011_763, w_003_069, w_010_103);
  not1 I011_764(w_011_764, w_007_701);
  or2  I011_765(w_011_765, w_003_018, w_004_1394);
  and2 I011_770(w_011_770, w_009_043, w_003_034);
  or2  I011_771(w_011_771, w_000_953, w_003_319);
  nand2 I011_773(w_011_773, w_001_1267, w_010_180);
  nand2 I011_775(w_011_775, w_010_076, w_005_1213);
  not1 I011_779(w_011_779, w_005_535);
  not1 I011_780(w_011_780, w_002_300);
  and2 I011_782(w_011_782, w_003_095, w_001_021);
  not1 I011_783(w_011_783, w_007_1616);
  nand2 I011_785(w_011_785, w_010_193, w_009_082);
  or2  I011_787(w_011_787, w_004_1023, w_009_072);
  and2 I011_790(w_011_790, w_001_422, w_003_040);
  not1 I011_791(w_011_791, w_003_066);
  nand2 I011_794(w_011_794, w_009_100, w_010_038);
  not1 I011_795(w_011_795, w_005_173);
  nand2 I011_796(w_011_796, w_002_319, w_005_127);
  nand2 I011_798(w_011_798, w_006_004, w_005_644);
  not1 I011_800(w_011_800, w_007_814);
  and2 I011_802(w_011_802, w_002_488, w_002_346);
  and2 I011_803(w_011_803, w_003_205, w_010_068);
  or2  I011_804(w_011_804, w_003_010, w_007_772);
  or2  I011_805(w_011_805, w_003_176, w_004_1276);
  and2 I011_809(w_011_809, w_010_284, w_006_174);
  and2 I011_810(w_011_810, w_006_225, w_008_526);
  or2  I011_811(w_011_811, w_008_645, w_001_1496);
  or2  I011_813(w_011_813, w_004_1135, w_006_186);
  not1 I011_814(w_011_814, w_005_1167);
  nand2 I011_815(w_011_815, w_010_141, w_000_247);
  or2  I011_816(w_011_816, w_009_083, w_006_228);
  and2 I011_817(w_011_817, w_010_181, w_000_461);
  nand2 I011_819(w_011_819, w_006_078, w_005_1622);
  or2  I011_822(w_011_822, w_009_078, w_008_228);
  nand2 I011_826(w_011_826, w_008_609, w_009_003);
  nand2 I011_829(w_011_829, w_001_1014, w_009_053);
  nand2 I011_830(w_011_830, w_010_223, w_004_529);
  and2 I011_832(w_011_832, w_001_1665, w_004_1549);
  and2 I011_833(w_011_833, w_008_056, w_005_860);
  or2  I011_835(w_011_835, w_007_1323, w_006_302);
  and2 I011_836(w_011_836, w_009_006, w_001_1321);
  nand2 I011_837(w_011_837, w_006_204, w_003_138);
  not1 I011_838(w_011_838, w_002_312);
  nand2 I011_839(w_011_839, w_006_120, w_009_052);
  not1 I011_840(w_011_840, w_001_1585);
  nand2 I011_845(w_011_845, w_009_091, w_007_869);
  nand2 I011_846(w_011_846, w_003_314, w_008_127);
  and2 I011_848(w_011_848, w_007_054, w_003_053);
  and2 I011_849(w_011_849, w_009_005, w_010_049);
  or2  I011_850(w_011_850, w_002_034, w_006_185);
  and2 I011_852(w_011_852, w_009_006, w_000_875);
  not1 I011_853(w_011_853, w_005_228);
  nand2 I011_854(w_011_854, w_010_229, w_002_336);
  nand2 I011_856(w_011_856, w_008_365, w_006_305);
  or2  I011_857(w_011_857, w_001_554, w_006_207);
  or2  I011_858(w_011_858, w_002_183, w_010_019);
  and2 I011_861(w_011_861, w_007_941, w_001_1281);
  nand2 I011_862(w_011_862, w_010_334, w_001_316);
  not1 I011_865(w_011_865, w_006_284);
  and2 I011_866(w_011_866, w_005_1381, w_006_088);
  and2 I011_867(w_011_867, w_005_1274, w_004_1611);
  not1 I011_869(w_011_869, w_008_096);
  or2  I011_870(w_011_870, w_009_007, w_009_041);
  not1 I011_871(w_011_871, w_003_056);
  nand2 I011_872(w_011_872, w_001_453, w_000_1022);
  or2  I011_875(w_011_875, w_006_009, w_003_256);
  not1 I011_876(w_011_876, w_007_354);
  and2 I011_877(w_011_877, w_006_048, w_006_189);
  not1 I011_878(w_011_878, w_006_271);
  not1 I011_879(w_011_879, w_007_091);
  or2  I011_881(w_011_881, w_008_327, w_000_101);
  not1 I011_883(w_011_883, w_000_1769);
  not1 I012_000(w_012_000, w_003_017);
  nand2 I012_002(w_012_002, w_000_1690, w_001_212);
  or2  I012_003(w_012_003, w_000_1033, w_009_057);
  not1 I012_006(w_012_006, w_008_076);
  or2  I012_007(w_012_007, w_003_175, w_000_488);
  or2  I012_008(w_012_008, w_003_251, w_000_655);
  not1 I012_011(w_012_011, w_009_095);
  or2  I012_016(w_012_016, w_004_1594, w_007_042);
  not1 I012_017(w_012_017, w_005_310);
  not1 I012_018(w_012_018, w_000_000);
  or2  I012_020(w_012_020, w_010_348, w_007_330);
  or2  I012_021(w_012_021, w_011_100, w_001_143);
  or2  I012_022(w_012_022, w_002_035, w_006_335);
  and2 I012_023(w_012_023, w_002_367, w_011_204);
  or2  I012_025(w_012_025, w_002_372, w_004_590);
  not1 I012_026(w_012_026, w_005_652);
  or2  I012_027(w_012_027, w_001_958, w_006_268);
  and2 I012_029(w_012_029, w_002_081, w_006_061);
  not1 I012_031(w_012_031, w_003_141);
  nand2 I012_033(w_012_033, w_000_1114, w_008_216);
  nand2 I012_034(w_012_034, w_009_055, w_010_256);
  or2  I012_035(w_012_035, w_010_128, w_001_1616);
  and2 I012_036(w_012_036, w_007_1054, w_004_1563);
  not1 I012_039(w_012_039, w_007_043);
  and2 I012_040(w_012_040, w_003_259, w_004_157);
  not1 I012_041(w_012_041, w_006_223);
  and2 I012_042(w_012_042, w_004_156, w_009_052);
  or2  I012_043(w_012_043, w_009_002, w_009_044);
  nand2 I012_044(w_012_044, w_000_1008, w_007_722);
  or2  I012_045(w_012_045, w_011_665, w_005_278);
  not1 I012_049(w_012_049, w_005_182);
  or2  I012_050(w_012_050, w_002_023, w_008_069);
  or2  I012_051(w_012_051, w_003_056, w_002_482);
  or2  I012_052(w_012_052, w_011_436, w_001_575);
  and2 I012_053(w_012_053, w_001_331, w_000_1565);
  nand2 I012_054(w_012_054, w_007_543, w_011_733);
  not1 I012_056(w_012_056, w_004_1422);
  and2 I012_058(w_012_058, w_008_810, w_002_011);
  nand2 I012_059(w_012_059, w_007_151, w_003_056);
  or2  I012_061(w_012_061, w_003_164, w_008_396);
  or2  I012_065(w_012_065, w_004_1481, w_000_323);
  and2 I012_066(w_012_066, w_008_699, w_010_251);
  and2 I012_067(w_012_067, w_008_234, w_004_528);
  nand2 I012_068(w_012_068, w_001_432, w_009_053);
  not1 I012_071(w_012_071, w_004_1228);
  not1 I012_073(w_012_073, w_003_193);
  not1 I012_075(w_012_075, w_003_131);
  nand2 I012_076(w_012_076, w_003_137, w_001_851);
  nand2 I012_077(w_012_077, w_003_048, w_005_532);
  not1 I012_078(w_012_078, w_002_383);
  nand2 I012_079(w_012_079, w_004_579, w_003_240);
  not1 I012_083(w_012_083, w_002_399);
  nand2 I012_085(w_012_085, w_006_199, w_005_953);
  not1 I012_087(w_012_087, w_006_169);
  or2  I012_090(w_012_090, w_010_227, w_007_1477);
  not1 I012_091(w_012_091, w_008_531);
  and2 I012_093(w_012_093, w_000_007, w_006_309);
  or2  I012_094(w_012_094, w_004_543, w_002_116);
  not1 I012_095(w_012_095, w_008_850);
  nand2 I012_096(w_012_096, w_003_070, w_007_1140);
  nand2 I012_097(w_012_097, w_009_043, w_002_526);
  and2 I012_099(w_012_099, w_008_402, w_004_513);
  not1 I012_100(w_012_100, w_002_072);
  nand2 I012_101(w_012_101, w_006_061, w_001_1342);
  nand2 I012_102(w_012_102, w_010_216, w_011_753);
  and2 I012_104(w_012_104, w_005_402, w_009_003);
  and2 I012_105(w_012_105, w_010_027, w_004_167);
  or2  I012_106(w_012_106, w_000_680, w_000_270);
  not1 I012_107(w_012_107, w_003_308);
  or2  I012_109(w_012_109, w_002_098, w_001_1657);
  or2  I012_110(w_012_110, w_004_1533, w_001_295);
  nand2 I012_111(w_012_111, w_010_112, w_011_676);
  not1 I012_112(w_012_112, w_007_103);
  or2  I012_116(w_012_116, w_007_1522, w_008_811);
  or2  I012_119(w_012_119, w_011_002, w_000_1451);
  and2 I012_122(w_012_122, w_008_683, w_010_287);
  not1 I012_123(w_012_123, w_001_1509);
  nand2 I012_125(w_012_125, w_008_303, w_010_156);
  nand2 I012_129(w_012_129, w_010_021, w_006_330);
  not1 I012_130(w_012_130, w_007_1223);
  not1 I012_132(w_012_132, w_009_033);
  and2 I012_133(w_012_133, w_010_401, w_002_159);
  and2 I012_137(w_012_137, w_003_268, w_003_266);
  nand2 I012_139(w_012_139, w_008_681, w_011_171);
  and2 I012_141(w_012_141, w_000_320, w_009_106);
  nand2 I012_142(w_012_142, w_005_056, w_001_1070);
  nand2 I012_143(w_012_143, w_005_402, w_007_680);
  and2 I012_144(w_012_144, w_008_479, w_009_007);
  and2 I012_145(w_012_145, w_004_1428, w_001_859);
  nand2 I012_146(w_012_146, w_001_404, w_005_1653);
  or2  I012_147(w_012_147, w_009_090, w_001_068);
  or2  I012_153(w_012_153, w_005_008, w_010_267);
  or2  I012_154(w_012_154, w_011_193, w_007_162);
  or2  I012_155(w_012_155, w_011_489, w_001_173);
  nand2 I012_156(w_012_156, w_009_015, w_003_240);
  not1 I012_157(w_012_157, w_008_047);
  and2 I012_159(w_012_159, w_004_1827, w_005_758);
  not1 I012_161(w_012_161, w_008_453);
  nand2 I012_162(w_012_162, w_000_1827, w_008_065);
  not1 I012_163(w_012_163, w_005_880);
  not1 I012_164(w_012_164, w_001_1019);
  not1 I012_165(w_012_165, w_008_094);
  nand2 I012_166(w_012_166, w_010_324, w_006_322);
  nand2 I012_168(w_012_168, w_004_487, w_003_110);
  and2 I012_169(w_012_169, w_000_297, w_000_1900);
  not1 I012_170(w_012_170, w_009_050);
  nand2 I012_171(w_012_171, w_005_069, w_005_756);
  not1 I012_172(w_012_172, w_005_933);
  or2  I012_173(w_012_173, w_003_030, w_004_561);
  nand2 I012_174(w_012_174, w_010_041, w_011_056);
  and2 I012_175(w_012_175, w_003_255, w_011_022);
  nand2 I012_176(w_012_176, w_004_087, w_007_947);
  or2  I012_177(w_012_177, w_008_244, w_001_1534);
  and2 I012_180(w_012_180, w_009_107, w_009_072);
  nand2 I012_181(w_012_181, w_006_175, w_006_053);
  or2  I012_183(w_012_183, w_006_022, w_010_331);
  and2 I012_184(w_012_184, w_004_701, w_010_283);
  or2  I012_186(w_012_186, w_004_1708, w_004_1250);
  and2 I012_187(w_012_187, w_003_160, w_004_922);
  or2  I012_188(w_012_188, w_005_261, w_003_046);
  or2  I012_189(w_012_189, w_008_016, w_007_966);
  not1 I012_191(w_012_191, w_011_764);
  and2 I012_193(w_012_193, w_007_1520, w_000_745);
  and2 I012_194(w_012_194, w_008_712, w_000_1838);
  nand2 I012_195(w_012_195, w_010_090, w_002_128);
  nand2 I012_196(w_012_196, w_010_098, w_003_264);
  and2 I012_198(w_012_198, w_004_1109, w_011_080);
  nand2 I012_199(w_012_199, w_010_003, w_007_1313);
  and2 I012_201(w_012_201, w_001_234, w_007_215);
  and2 I012_202(w_012_202, w_009_063, w_007_1435);
  nand2 I012_204(w_012_204, w_007_053, w_000_1270);
  not1 I012_205(w_012_205, w_011_204);
  not1 I012_206(w_012_206, w_007_401);
  nand2 I012_209(w_012_209, w_009_036, w_006_109);
  not1 I012_210(w_012_210, w_010_096);
  or2  I012_211(w_012_211, w_007_051, w_005_658);
  and2 I012_212(w_012_212, w_004_809, w_001_1432);
  nand2 I012_213(w_012_213, w_007_1044, w_007_1061);
  nand2 I012_214(w_012_214, w_000_1503, w_006_053);
  not1 I012_215(w_012_215, w_009_094);
  or2  I012_216(w_012_216, w_006_122, w_000_1527);
  and2 I012_217(w_012_217, w_002_471, w_006_321);
  not1 I012_218(w_012_218, w_003_067);
  not1 I012_219(w_012_219, w_000_828);
  not1 I012_221(w_012_221, w_001_1119);
  not1 I012_222(w_012_222, w_008_569);
  nand2 I012_223(w_012_223, w_010_202, w_001_852);
  and2 I012_224(w_012_224, w_004_1792, w_011_128);
  not1 I012_227(w_012_227, w_006_280);
  not1 I012_228(w_012_228, w_009_007);
  nand2 I012_229(w_012_229, w_011_052, w_010_259);
  not1 I012_231(w_012_231, w_003_087);
  not1 I012_232(w_012_232, w_007_1590);
  nand2 I012_233(w_012_233, w_005_785, w_005_1628);
  and2 I012_235(w_012_235, w_011_044, w_001_1270);
  nand2 I012_236(w_012_236, w_000_1091, w_005_059);
  and2 I012_237(w_012_237, w_001_1675, w_007_1480);
  or2  I012_238(w_012_238, w_011_119, w_000_1118);
  or2  I012_239(w_012_239, w_003_028, w_003_192);
  and2 I012_240(w_012_240, w_006_168, w_007_001);
  or2  I012_241(w_012_241, w_011_856, w_005_025);
  not1 I012_242(w_012_242, w_008_657);
  or2  I012_243(w_012_243, w_002_391, w_005_1331);
  and2 I012_246(w_012_246, w_011_654, w_011_419);
  and2 I012_249(w_012_249, w_007_828, w_006_085);
  nand2 I012_250(w_012_250, w_011_000, w_010_197);
  nand2 I012_252(w_012_252, w_006_137, w_009_053);
  and2 I012_254(w_012_254, w_005_800, w_002_147);
  not1 I012_255(w_012_255, w_007_466);
  not1 I012_257(w_012_257, w_004_672);
  and2 I012_258(w_012_258, w_009_036, w_002_119);
  not1 I012_259(w_012_259, w_004_036);
  or2  I012_260(w_012_260, w_001_366, w_006_209);
  not1 I012_261(w_012_261, w_005_465);
  or2  I012_262(w_012_262, w_009_030, w_005_016);
  and2 I012_264(w_012_264, w_010_092, w_004_1080);
  and2 I012_265(w_012_265, w_004_1848, w_001_852);
  not1 I012_266(w_012_266, w_007_790);
  nand2 I012_268(w_012_268, w_009_078, w_000_216);
  nand2 I012_269(w_012_269, w_002_111, w_004_816);
  not1 I012_270(w_012_270, w_008_805);
  or2  I012_271(w_012_271, w_011_107, w_003_155);
  nand2 I012_272(w_012_272, w_003_184, w_007_1159);
  or2  I012_273(w_012_273, w_007_309, w_000_457);
  nand2 I012_274(w_012_274, w_004_753, w_002_173);
  not1 I012_276(w_012_276, w_006_121);
  and2 I012_277(w_012_277, w_007_1512, w_006_150);
  nand2 I012_278(w_012_278, w_001_1002, w_006_289);
  not1 I012_279(w_012_279, w_005_824);
  or2  I012_281(w_012_281, w_008_032, w_008_219);
  or2  I012_284(w_012_284, w_008_190, w_008_560);
  or2  I012_287(w_012_287, w_010_287, w_011_034);
  and2 I012_288(w_012_288, w_001_253, w_003_160);
  or2  I012_289(w_012_289, w_009_062, w_011_623);
  nand2 I012_290(w_012_290, w_000_579, w_011_857);
  nand2 I012_292(w_012_292, w_002_407, w_002_497);
  not1 I012_293(w_012_293, w_003_185);
  or2  I012_294(w_012_294, w_003_020, w_009_108);
  or2  I012_295(w_012_295, w_001_108, w_007_174);
  and2 I012_297(w_012_297, w_009_023, w_000_1746);
  nand2 I012_298(w_012_298, w_007_1190, w_002_105);
  nand2 I012_302(w_012_302, w_006_107, w_006_252);
  or2  I012_304(w_012_304, w_011_105, w_006_342);
  not1 I012_305(w_012_305, w_008_504);
  and2 I012_307(w_012_307, w_011_402, w_000_1525);
  or2  I012_310(w_012_310, w_011_700, w_006_300);
  and2 I012_314(w_012_314, w_004_249, w_003_091);
  nand2 I012_316(w_012_316, w_005_1392, w_003_127);
  or2  I012_317(w_012_317, w_000_424, w_007_247);
  not1 I012_319(w_012_319, w_009_025);
  and2 I012_320(w_012_320, w_002_429, w_000_470);
  nand2 I012_322(w_012_322, w_006_043, w_007_900);
  not1 I012_323(w_012_323, w_005_292);
  or2  I012_324(w_012_324, w_008_681, w_005_126);
  not1 I012_326(w_012_326, w_008_461);
  nand2 I012_327(w_012_327, w_005_015, w_005_1218);
  nand2 I012_328(w_012_328, w_004_248, w_006_118);
  and2 I012_329(w_012_329, w_001_1193, w_011_181);
  and2 I012_330(w_012_330, w_008_825, w_009_045);
  nand2 I012_332(w_012_332, w_003_192, w_009_027);
  not1 I012_334(w_012_334, w_008_830);
  not1 I012_336(w_012_336, w_008_660);
  not1 I012_337(w_012_337, w_009_085);
  not1 I012_338(w_012_338, w_006_135);
  nand2 I012_339(w_012_339, w_005_1182, w_001_781);
  not1 I012_340(w_012_340, w_008_524);
  not1 I012_341(w_012_341, w_009_103);
  or2  I012_342(w_012_342, w_010_194, w_003_036);
  or2  I012_343(w_012_343, w_011_334, w_011_006);
  nand2 I012_345(w_012_345, w_000_599, w_001_366);
  not1 I012_346(w_012_346, w_008_196);
  and2 I012_348(w_012_348, w_000_1234, w_001_021);
  and2 I012_349(w_012_349, w_003_006, w_007_379);
  nand2 I012_350(w_012_350, w_006_229, w_007_865);
  nand2 I012_351(w_012_351, w_005_1519, w_007_573);
  or2  I012_353(w_012_353, w_008_022, w_009_061);
  and2 I012_355(w_012_355, w_010_384, w_000_1250);
  nand2 I012_356(w_012_356, w_007_005, w_003_130);
  nand2 I012_357(w_012_357, w_010_271, w_002_343);
  not1 I012_362(w_012_362, w_006_175);
  or2  I012_364(w_012_364, w_000_1808, w_007_439);
  and2 I012_366(w_012_366, w_002_211, w_009_049);
  and2 I012_368(w_012_368, w_004_996, w_003_078);
  not1 I012_369(w_012_369, w_005_1088);
  and2 I012_370(w_012_370, w_004_590, w_002_037);
  nand2 I012_371(w_012_371, w_006_197, w_006_217);
  and2 I012_372(w_012_372, w_000_827, w_008_813);
  not1 I012_373(w_012_373, w_009_080);
  nand2 I012_374(w_012_374, w_000_1730, w_004_171);
  nand2 I012_375(w_012_375, w_000_1519, w_010_333);
  or2  I012_376(w_012_376, w_003_243, w_001_248);
  or2  I012_377(w_012_377, w_008_285, w_001_898);
  nand2 I012_378(w_012_378, w_007_188, w_011_432);
  and2 I012_384(w_012_384, w_005_096, w_001_130);
  and2 I012_387(w_012_387, w_009_081, w_008_052);
  not1 I012_388(w_012_388, w_001_378);
  or2  I012_390(w_012_390, w_001_163, w_011_424);
  and2 I012_392(w_012_392, w_000_1701, w_008_386);
  or2  I012_393(w_012_393, w_000_1184, w_010_403);
  or2  I012_394(w_012_394, w_009_111, w_002_470);
  nand2 I012_395(w_012_395, w_004_1681, w_008_593);
  and2 I012_399(w_012_399, w_006_314, w_008_616);
  or2  I012_400(w_012_400, w_001_279, w_000_943);
  and2 I012_401(w_012_401, w_008_023, w_009_036);
  or2  I012_402(w_012_402, w_000_155, w_008_465);
  nand2 I012_403(w_012_403, w_004_062, w_007_559);
  or2  I012_404(w_012_404, w_003_081, w_006_132);
  and2 I012_405(w_012_405, w_006_074, w_006_078);
  nand2 I012_406(w_012_406, w_004_428, w_000_892);
  nand2 I012_407(w_012_407, w_008_026, w_003_061);
  nand2 I012_409(w_012_409, w_011_533, w_007_346);
  and2 I012_410(w_012_410, w_000_573, w_006_130);
  or2  I012_411(w_012_411, w_002_244, w_003_004);
  nand2 I012_412(w_012_412, w_010_138, w_011_711);
  or2  I012_413(w_012_413, w_002_439, w_009_081);
  nand2 I012_416(w_012_416, w_009_062, w_000_1823);
  nand2 I012_421(w_012_421, w_007_929, w_006_289);
  and2 I012_422(w_012_422, w_000_383, w_004_1361);
  or2  I012_425(w_012_425, w_009_107, w_005_094);
  or2  I012_426(w_012_426, w_000_163, w_000_1213);
  or2  I012_428(w_012_428, w_002_047, w_001_906);
  and2 I012_429(w_012_429, w_010_199, w_002_487);
  nand2 I012_430(w_012_430, w_005_528, w_007_378);
  or2  I012_431(w_012_431, w_008_051, w_008_556);
  nand2 I012_435(w_012_435, w_002_546, w_011_265);
  and2 I012_436(w_012_436, w_010_406, w_000_1902);
  and2 I012_438(w_012_438, w_004_459, w_009_016);
  nand2 I012_441(w_012_441, w_011_517, w_008_681);
  not1 I012_442(w_012_442, w_004_1681);
  nand2 I012_445(w_012_445, w_003_050, w_004_799);
  and2 I012_446(w_012_446, w_003_203, w_000_635);
  and2 I012_447(w_012_447, w_009_038, w_008_599);
  and2 I012_449(w_012_449, w_011_856, w_007_417);
  or2  I012_450(w_012_450, w_000_1698, w_005_1038);
  and2 I012_451(w_012_451, w_004_057, w_003_124);
  and2 I012_452(w_012_452, w_007_987, w_000_172);
  not1 I012_453(w_012_453, w_008_133);
  or2  I012_454(w_012_454, w_004_035, w_001_068);
  and2 I012_455(w_012_455, w_003_312, w_000_839);
  nand2 I012_459(w_012_459, w_001_062, w_007_549);
  and2 I012_460(w_012_460, w_008_682, w_009_076);
  and2 I012_461(w_012_461, w_010_172, w_000_1794);
  not1 I012_464(w_012_464, w_010_414);
  or2  I012_465(w_012_465, w_000_1489, w_005_362);
  nand2 I012_466(w_012_466, w_004_1263, w_003_016);
  not1 I012_467(w_012_467, w_001_1181);
  not1 I012_468(w_012_468, w_011_126);
  not1 I012_469(w_012_469, w_009_055);
  nand2 I012_470(w_012_470, w_010_219, w_004_015);
  or2  I012_471(w_012_471, w_008_619, w_004_787);
  or2  I012_472(w_012_472, w_006_212, w_002_531);
  not1 I012_474(w_012_474, w_006_113);
  nand2 I012_475(w_012_475, w_011_763, w_002_211);
  not1 I012_476(w_012_476, w_000_401);
  or2  I012_477(w_012_477, w_010_199, w_005_123);
  and2 I012_478(w_012_478, w_006_081, w_008_212);
  not1 I012_482(w_012_482, w_007_305);
  and2 I012_484(w_012_484, w_011_688, w_006_165);
  and2 I012_486(w_012_486, w_003_306, w_005_1410);
  or2  I012_487(w_012_487, w_009_039, w_002_205);
  not1 I012_488(w_012_488, w_010_093);
  nand2 I012_490(w_012_490, w_009_027, w_007_340);
  or2  I012_493(w_012_493, w_008_092, w_002_416);
  and2 I012_494(w_012_494, w_009_067, w_006_343);
  or2  I012_497(w_012_497, w_011_716, w_005_160);
  nand2 I012_500(w_012_500, w_011_426, w_006_221);
  and2 I012_502(w_012_502, w_002_387, w_002_434);
  not1 I012_503(w_012_503, w_004_187);
  nand2 I012_504(w_012_504, w_004_1788, w_000_947);
  nand2 I012_505(w_012_505, w_003_032, w_002_005);
  nand2 I012_506(w_012_506, w_008_175, w_002_403);
  or2  I012_507(w_012_507, w_002_587, w_011_751);
  or2  I012_508(w_012_508, w_002_332, w_009_048);
  and2 I012_509(w_012_509, w_003_118, w_010_207);
  or2  I012_510(w_012_510, w_001_1003, w_009_106);
  nand2 I012_511(w_012_511, w_001_1521, w_011_751);
  and2 I012_512(w_012_512, w_010_210, w_005_1469);
  and2 I012_513(w_012_513, w_006_131, w_011_853);
  not1 I012_514(w_012_514, w_004_663);
  nand2 I012_515(w_012_515, w_005_1159, w_003_008);
  nand2 I012_517(w_012_517, w_004_1784, w_010_193);
  nand2 I012_519(w_012_519, w_003_292, w_007_189);
  nand2 I012_520(w_012_520, w_006_011, w_002_390);
  not1 I012_521(w_012_521, w_001_183);
  not1 I012_522(w_012_522, w_008_143);
  nand2 I012_523(w_012_523, w_009_011, w_006_243);
  not1 I012_524(w_012_524, w_011_716);
  and2 I012_525(w_012_525, w_008_373, w_001_1429);
  nand2 I012_526(w_012_526, w_000_1392, w_002_163);
  and2 I012_527(w_012_527, w_007_128, w_010_191);
  nand2 I012_529(w_012_529, w_000_731, w_003_044);
  not1 I012_530(w_012_530, w_004_077);
  or2  I012_531(w_012_531, w_008_167, w_008_680);
  and2 I012_535(w_012_535, w_000_1498, w_005_1641);
  not1 I012_536(w_012_536, w_010_303);
  or2  I012_537(w_012_537, w_010_234, w_002_431);
  and2 I012_538(w_012_538, w_002_328, w_004_362);
  not1 I012_541(w_012_541, w_000_699);
  not1 I012_545(w_012_545, w_009_055);
  not1 I012_546(w_012_546, w_011_638);
  not1 I012_547(w_012_547, w_002_117);
  not1 I012_550(w_012_550, w_010_022);
  or2  I012_551(w_012_551, w_001_887, w_000_1904);
  nand2 I012_552(w_012_552, w_010_269, w_000_748);
  or2  I012_554(w_012_554, w_005_128, w_000_1652);
  or2  I012_555(w_012_555, w_006_002, w_005_411);
  and2 I012_556(w_012_556, w_008_209, w_008_317);
  nand2 I012_557(w_012_557, w_010_339, w_000_1905);
  or2  I012_558(w_012_558, w_000_246, w_004_1734);
  and2 I012_559(w_012_559, w_004_834, w_006_155);
  and2 I012_560(w_012_560, w_004_1292, w_005_197);
  and2 I012_561(w_012_561, w_006_206, w_006_315);
  nand2 I012_563(w_012_563, w_003_260, w_002_365);
  not1 I012_564(w_012_564, w_003_237);
  or2  I012_567(w_012_567, w_010_092, w_006_070);
  or2  I012_569(w_012_569, w_007_103, w_011_699);
  not1 I012_570(w_012_570, w_002_163);
  and2 I012_571(w_012_571, w_008_698, w_003_037);
  or2  I012_572(w_012_572, w_011_441, w_005_541);
  or2  I012_573(w_012_573, w_000_025, w_008_615);
  not1 I012_574(w_012_574, w_006_173);
  and2 I012_578(w_012_578, w_003_172, w_002_094);
  not1 I012_579(w_012_579, w_007_175);
  nand2 I012_580(w_012_580, w_007_200, w_011_182);
  nand2 I012_581(w_012_581, w_006_124, w_011_327);
  and2 I012_582(w_012_582, w_004_141, w_009_108);
  not1 I012_585(w_012_585, w_011_256);
  and2 I012_586(w_012_586, w_009_086, w_003_040);
  or2  I012_587(w_012_587, w_002_013, w_001_1521);
  and2 I012_588(w_012_588, w_011_137, w_003_094);
  or2  I012_589(w_012_589, w_007_907, w_006_051);
  or2  I012_590(w_012_590, w_007_734, w_002_010);
  and2 I012_591(w_012_591, w_010_367, w_002_194);
  nand2 I012_592(w_012_592, w_010_108, w_001_289);
  and2 I012_594(w_012_594, w_005_187, w_005_232);
  nand2 I012_596(w_012_596, w_009_000, w_010_277);
  and2 I012_597(w_012_597, w_010_121, w_003_308);
  nand2 I012_598(w_012_598, w_007_018, w_003_000);
  nand2 I012_599(w_012_599, w_011_067, w_002_094);
  nand2 I012_603(w_012_603, w_003_089, w_001_1163);
  or2  I012_607(w_012_607, w_003_035, w_008_216);
  or2  I012_608(w_012_608, w_011_071, w_010_288);
  not1 I012_609(w_012_609, w_007_1279);
  and2 I012_612(w_012_612, w_006_303, w_004_153);
  or2  I012_613(w_012_613, w_002_223, w_002_437);
  and2 I012_614(w_012_614, w_009_072, w_004_173);
  nand2 I012_616(w_012_616, w_003_302, w_005_394);
  or2  I012_617(w_012_617, w_010_118, w_009_039);
  not1 I012_618(w_012_618, w_010_005);
  or2  I012_619(w_012_619, w_006_194, w_003_120);
  or2  I012_620(w_012_620, w_009_093, w_010_326);
  not1 I012_621(w_012_621, w_006_156);
  and2 I012_625(w_012_625, w_005_156, w_006_279);
  not1 I012_626(w_012_626, w_009_071);
  nand2 I012_627(w_012_627, w_006_293, w_005_576);
  nand2 I012_628(w_012_628, w_004_1076, w_010_227);
  or2  I012_629(w_012_629, w_006_260, w_008_456);
  and2 I012_631(w_012_631, w_000_1334, w_001_601);
  or2  I012_632(w_012_632, w_007_288, w_003_256);
  and2 I012_633(w_012_633, w_011_582, w_001_1540);
  nand2 I012_635(w_012_635, w_010_205, w_008_300);
  nand2 I012_636(w_012_636, w_008_756, w_007_077);
  nand2 I012_637(w_012_637, w_000_1245, w_000_1906);
  nand2 I012_639(w_012_639, w_008_011, w_011_283);
  not1 I012_640(w_012_640, w_000_708);
  and2 I012_641(w_012_641, w_004_616, w_007_1310);
  nand2 I012_642(w_012_642, w_003_011, w_002_418);
  and2 I012_643(w_012_643, w_001_1065, w_004_1306);
  or2  I012_646(w_012_646, w_003_179, w_007_271);
  not1 I012_648(w_012_648, w_007_058);
  or2  I012_649(w_012_649, w_002_452, w_001_467);
  and2 I012_650(w_012_650, w_005_125, w_003_197);
  nand2 I012_652(w_012_652, w_002_205, w_004_1082);
  and2 I012_653(w_012_653, w_011_445, w_004_1599);
  or2  I012_654(w_012_654, w_000_194, w_007_1579);
  and2 I012_655(w_012_655, w_008_660, w_003_081);
  or2  I012_656(w_012_656, w_003_039, w_006_194);
  and2 I012_657(w_012_657, w_003_291, w_007_1341);
  or2  I012_659(w_012_659, w_010_262, w_003_210);
  or2  I012_660(w_012_660, w_000_1886, w_011_783);
  or2  I012_661(w_012_661, w_008_791, w_011_435);
  and2 I012_662(w_012_662, w_008_032, w_003_190);
  and2 I012_663(w_012_663, w_000_1377, w_003_227);
  nand2 I012_666(w_012_666, w_011_583, w_010_114);
  and2 I012_667(w_012_667, w_010_352, w_000_325);
  and2 I013_000(w_013_000, w_006_088, w_007_317);
  and2 I013_001(w_013_001, w_008_804, w_007_013);
  and2 I013_002(w_013_002, w_000_340, w_003_126);
  and2 I013_003(w_013_003, w_007_920, w_008_345);
  and2 I013_004(w_013_004, w_006_240, w_006_079);
  nand2 I013_006(w_013_006, w_005_1059, w_004_1448);
  not1 I013_008(w_013_008, w_007_270);
  not1 I013_009(w_013_009, w_012_020);
  nand2 I013_010(w_013_010, w_006_261, w_012_535);
  or2  I013_011(w_013_011, w_007_131, w_003_305);
  and2 I013_012(w_013_012, w_004_984, w_006_011);
  nand2 I013_013(w_013_013, w_011_798, w_006_186);
  not1 I013_014(w_013_014, w_009_091);
  not1 I013_015(w_013_015, w_009_009);
  nand2 I013_016(w_013_016, w_009_044, w_010_343);
  nand2 I013_017(w_013_017, w_005_313, w_012_608);
  or2  I013_018(w_013_018, w_006_032, w_007_1596);
  and2 I013_019(w_013_019, w_012_580, w_012_180);
  and2 I013_021(w_013_021, w_003_186, w_002_393);
  and2 I013_022(w_013_022, w_000_1904, w_005_1074);
  nand2 I013_023(w_013_023, w_003_187, w_003_299);
  and2 I013_024(w_013_024, w_005_661, w_000_1776);
  or2  I013_025(w_013_025, w_005_1553, w_012_350);
  or2  I013_026(w_013_026, w_000_959, w_010_337);
  not1 I013_027(w_013_027, w_009_012);
  and2 I013_028(w_013_028, w_012_618, w_012_236);
  not1 I013_029(w_013_029, w_006_278);
  or2  I013_030(w_013_030, w_009_025, w_005_1138);
  or2  I013_031(w_013_031, w_010_116, w_010_336);
  or2  I013_032(w_013_032, w_003_242, w_000_1644);
  nand2 I013_033(w_013_033, w_000_603, w_012_431);
  not1 I013_035(w_013_035, w_012_564);
  and2 I013_036(w_013_036, w_006_226, w_004_1138);
  or2  I013_038(w_013_038, w_005_1113, w_005_1369);
  or2  I013_040(w_013_040, w_008_513, w_003_080);
  or2  I013_041(w_013_041, w_001_1049, w_001_1195);
  and2 I013_043(w_013_043, w_007_109, w_009_089);
  not1 I013_044(w_013_044, w_005_944);
  nand2 I013_045(w_013_045, w_011_313, w_007_126);
  nand2 I013_046(w_013_046, w_003_204, w_008_200);
  or2  I013_047(w_013_047, w_011_388, w_012_031);
  or2  I013_048(w_013_048, w_000_562, w_005_872);
  and2 I013_049(w_013_049, w_004_764, w_007_411);
  or2  I013_050(w_013_050, w_006_268, w_011_852);
  or2  I013_051(w_013_051, w_012_345, w_000_1577);
  and2 I013_052(w_013_052, w_012_339, w_008_684);
  nand2 I013_053(w_013_053, w_006_248, w_000_1023);
  nand2 I013_054(w_013_054, w_005_160, w_002_144);
  and2 I013_055(w_013_055, w_007_975, w_010_309);
  nand2 I013_057(w_013_057, w_002_400, w_004_1706);
  or2  I013_058(w_013_058, w_004_1284, w_012_384);
  nand2 I013_059(w_013_059, w_009_061, w_009_030);
  or2  I013_060(w_013_060, w_011_173, w_005_188);
  or2  I013_061(w_013_061, w_009_109, w_004_286);
  and2 I013_062(w_013_062, w_003_280, w_001_252);
  nand2 I013_063(w_013_063, w_008_130, w_002_470);
  or2  I013_064(w_013_064, w_011_492, w_001_296);
  not1 I013_066(w_013_066, w_009_090);
  and2 I013_067(w_013_067, w_004_1191, w_011_161);
  and2 I013_068(w_013_068, w_003_216, w_004_1792);
  and2 I013_069(w_013_069, w_005_087, w_000_1907);
  or2  I013_070(w_013_070, w_005_316, w_001_984);
  not1 I013_072(w_013_072, w_008_315);
  or2  I013_073(w_013_073, w_007_1318, w_007_1230);
  or2  I013_074(w_013_074, w_005_1511, w_009_101);
  nand2 I013_075(w_013_075, w_000_918, w_005_153);
  or2  I013_076(w_013_076, w_006_142, w_008_749);
  not1 I013_077(w_013_077, w_012_598);
  not1 I013_078(w_013_078, w_003_000);
  or2  I013_080(w_013_080, w_012_240, w_002_304);
  or2  I013_081(w_013_081, w_002_571, w_006_044);
  nand2 I013_083(w_013_083, w_007_144, w_004_705);
  not1 I013_084(w_013_084, w_004_1535);
  nand2 I013_085(w_013_085, w_009_065, w_010_315);
  nand2 I013_086(w_013_086, w_007_1090, w_007_756);
  not1 I013_087(w_013_087, w_011_770);
  nand2 I013_088(w_013_088, w_000_1413, w_000_185);
  or2  I013_089(w_013_089, w_006_309, w_007_1406);
  and2 I013_090(w_013_090, w_001_1550, w_003_290);
  or2  I013_091(w_013_091, w_009_001, w_012_122);
  not1 I013_092(w_013_092, w_011_573);
  not1 I013_093(w_013_093, w_006_211);
  not1 I013_094(w_013_094, w_003_001);
  not1 I013_095(w_013_095, w_000_200);
  not1 I013_096(w_013_096, w_008_246);
  nand2 I013_097(w_013_097, w_003_226, w_000_1878);
  and2 I013_098(w_013_098, w_012_071, w_009_020);
  not1 I013_099(w_013_099, w_004_1095);
  nand2 I013_100(w_013_100, w_003_233, w_012_033);
  not1 I013_101(w_013_101, w_012_166);
  or2  I013_102(w_013_102, w_006_043, w_003_280);
  nand2 I013_103(w_013_103, w_012_051, w_011_365);
  not1 I013_104(w_013_104, w_003_271);
  nand2 I013_105(w_013_105, w_002_315, w_012_145);
  not1 I013_106(w_013_106, w_003_167);
  not1 I013_107(w_013_107, w_001_1299);
  nand2 I013_108(w_013_108, w_008_801, w_004_535);
  or2  I013_109(w_013_109, w_001_501, w_009_037);
  nand2 I013_110(w_013_110, w_011_461, w_005_032);
  not1 I013_111(w_013_111, w_003_081);
  not1 I013_112(w_013_112, w_002_128);
  and2 I013_113(w_013_113, w_009_040, w_000_612);
  and2 I013_114(w_013_114, w_005_059, w_002_088);
  or2  I013_115(w_013_115, w_012_077, w_004_1436);
  not1 I013_116(w_013_116, w_005_289);
  or2  I013_117(w_013_117, w_009_021, w_002_326);
  nand2 I013_118(w_013_118, w_010_133, w_006_158);
  not1 I013_119(w_013_119, w_008_453);
  not1 I013_120(w_013_120, w_004_607);
  nand2 I013_121(w_013_121, w_008_067, w_012_468);
  nand2 I013_122(w_013_122, w_011_009, w_008_825);
  nand2 I013_123(w_013_123, w_006_123, w_008_044);
  or2  I013_124(w_013_124, w_006_131, w_012_269);
  not1 I013_125(w_013_125, w_012_017);
  and2 I013_126(w_013_126, w_006_003, w_009_071);
  or2  I013_127(w_013_127, w_003_182, w_010_092);
  and2 I013_131(w_013_131, w_000_1093, w_006_295);
  nand2 I013_132(w_013_132, w_007_337, w_010_011);
  and2 I013_133(w_013_133, w_006_082, w_006_306);
  and2 I013_134(w_013_134, w_003_038, w_002_256);
  or2  I013_135(w_013_135, w_008_310, w_012_222);
  not1 I013_136(w_013_136, w_008_544);
  or2  I013_137(w_013_137, w_002_128, w_005_263);
  nand2 I013_139(w_013_139, w_005_160, w_009_083);
  or2  I013_140(w_013_140, w_004_430, w_007_105);
  and2 I013_141(w_013_141, w_009_001, w_002_092);
  and2 I013_142(w_013_142, w_002_072, w_001_1306);
  nand2 I013_143(w_013_143, w_001_895, w_004_152);
  not1 I013_144(w_013_144, w_003_303);
  or2  I013_145(w_013_145, w_000_864, w_010_082);
  or2  I013_147(w_013_147, w_008_185, w_005_408);
  or2  I013_148(w_013_148, w_009_040, w_008_326);
  nand2 I013_149(w_013_149, w_011_217, w_011_350);
  and2 I013_150(w_013_150, w_002_198, w_007_354);
  or2  I013_151(w_013_151, w_012_442, w_002_302);
  or2  I013_153(w_013_153, w_006_147, w_000_303);
  nand2 I013_154(w_013_154, w_007_1063, w_012_341);
  nand2 I013_155(w_013_155, w_009_008, w_009_012);
  or2  I013_156(w_013_156, w_008_702, w_003_037);
  and2 I013_159(w_013_159, w_011_522, w_001_1057);
  or2  I013_160(w_013_160, w_003_112, w_005_586);
  nand2 I013_161(w_013_161, w_006_219, w_009_109);
  nand2 I013_162(w_013_162, w_008_809, w_010_021);
  nand2 I013_163(w_013_163, w_001_1151, w_012_250);
  nand2 I013_164(w_013_164, w_004_771, w_004_1228);
  and2 I013_165(w_013_165, w_001_1278, w_004_670);
  nand2 I013_167(w_013_167, w_012_240, w_006_108);
  not1 I013_168(w_013_168, w_000_041);
  nand2 I013_169(w_013_169, w_010_062, w_011_620);
  nand2 I013_170(w_013_170, w_010_002, w_001_1067);
  not1 I013_171(w_013_171, w_005_296);
  not1 I013_172(w_013_172, w_008_709);
  and2 I013_173(w_013_173, w_012_613, w_004_931);
  and2 I013_174(w_013_174, w_006_282, w_010_096);
  and2 I013_175(w_013_175, w_007_382, w_007_120);
  or2  I013_176(w_013_176, w_007_579, w_000_1908);
  not1 I013_177(w_013_177, w_011_764);
  and2 I013_178(w_013_178, w_001_310, w_009_042);
  and2 I013_179(w_013_179, w_004_640, w_012_369);
  or2  I013_180(w_013_180, w_006_276, w_004_687);
  not1 I013_181(w_013_181, w_003_179);
  nand2 I013_182(w_013_182, w_011_669, w_005_362);
  nand2 I013_183(w_013_183, w_012_273, w_006_232);
  and2 I013_184(w_013_184, w_006_308, w_007_889);
  nand2 I013_185(w_013_185, w_004_1603, w_011_459);
  and2 I013_186(w_013_186, w_000_1181, w_006_092);
  or2  I013_187(w_013_187, w_011_051, w_007_110);
  nand2 I013_188(w_013_188, w_003_000, w_001_808);
  not1 I013_189(w_013_189, w_009_059);
  and2 I013_190(w_013_190, w_005_659, w_008_024);
  nand2 I013_191(w_013_191, w_002_590, w_005_029);
  not1 I013_192(w_013_192, w_004_516);
  nand2 I013_194(w_013_194, w_001_882, w_000_089);
  and2 I013_197(w_013_197, w_012_196, w_000_972);
  and2 I013_198(w_013_198, w_001_1667, w_002_011);
  not1 I013_199(w_013_199, w_011_097);
  nand2 I013_201(w_013_201, w_000_1676, w_002_491);
  nand2 I013_203(w_013_203, w_008_152, w_011_323);
  nand2 I013_205(w_013_205, w_012_655, w_004_1093);
  or2  I013_206(w_013_206, w_010_154, w_009_019);
  and2 I013_207(w_013_207, w_011_803, w_010_002);
  nand2 I013_209(w_013_209, w_004_1539, w_010_294);
  not1 I013_210(w_013_210, w_007_320);
  not1 I013_211(w_013_211, w_004_964);
  or2  I013_212(w_013_212, w_006_251, w_004_1645);
  and2 I013_214(w_013_214, w_006_009, w_006_125);
  or2  I013_215(w_013_215, w_003_257, w_009_046);
  and2 I013_216(w_013_216, w_002_397, w_000_470);
  nand2 I013_217(w_013_217, w_007_790, w_000_1403);
  not1 I013_219(w_013_219, w_004_1600);
  nand2 I013_221(w_013_221, w_006_265, w_012_502);
  not1 I013_222(w_013_222, w_010_304);
  and2 I013_223(w_013_223, w_007_1080, w_008_019);
  not1 I013_225(w_013_225, w_001_756);
  or2  I013_226(w_013_226, w_003_010, w_005_116);
  nand2 I013_227(w_013_227, w_009_081, w_002_237);
  or2  I013_228(w_013_228, w_009_034, w_008_678);
  or2  I013_229(w_013_229, w_005_982, w_001_065);
  not1 I013_230(w_013_230, w_009_100);
  and2 I013_231(w_013_231, w_009_087, w_005_832);
  nand2 I013_233(w_013_233, w_010_334, w_009_024);
  and2 I013_234(w_013_234, w_000_794, w_000_304);
  and2 I013_235(w_013_235, w_010_141, w_003_028);
  or2  I013_236(w_013_236, w_004_733, w_009_033);
  or2  I013_237(w_013_237, w_004_1035, w_009_028);
  not1 I013_239(w_013_239, w_012_272);
  and2 I013_240(w_013_240, w_010_135, w_002_108);
  or2  I013_242(w_013_242, w_001_1540, w_006_079);
  or2  I013_243(w_013_243, w_002_057, w_009_035);
  and2 I013_244(w_013_244, w_007_655, w_009_049);
  or2  I013_245(w_013_245, w_008_853, w_006_224);
  and2 I013_247(w_013_247, w_001_1282, w_007_082);
  or2  I013_248(w_013_248, w_006_019, w_002_357);
  nand2 I013_249(w_013_249, w_004_1398, w_006_146);
  or2  I013_250(w_013_250, w_005_1533, w_004_1321);
  nand2 I013_251(w_013_251, w_005_794, w_005_106);
  not1 I013_252(w_013_252, w_011_557);
  and2 I013_253(w_013_253, w_005_186, w_006_215);
  nand2 I013_254(w_013_254, w_001_994, w_003_239);
  or2  I013_255(w_013_255, w_007_822, w_011_125);
  or2  I013_257(w_013_257, w_006_198, w_006_110);
  and2 I013_258(w_013_258, w_011_579, w_003_182);
  and2 I013_259(w_013_259, w_012_314, w_011_015);
  not1 I013_260(w_013_260, w_004_830);
  and2 I013_261(w_013_261, w_009_029, w_011_833);
  not1 I013_263(w_013_263, w_012_659);
  nand2 I013_264(w_013_264, w_005_1209, w_008_464);
  or2  I013_265(w_013_265, w_008_530, w_002_156);
  and2 I013_266(w_013_266, w_003_105, w_007_030);
  nand2 I013_267(w_013_267, w_000_861, w_006_182);
  not1 I013_268(w_013_268, w_006_055);
  or2  I013_270(w_013_270, w_011_143, w_011_056);
  not1 I013_271(w_013_271, w_005_150);
  or2  I013_272(w_013_272, w_011_703, w_000_1527);
  nand2 I013_273(w_013_273, w_007_023, w_004_117);
  or2  I013_274(w_013_274, w_002_166, w_011_758);
  nand2 I013_275(w_013_275, w_012_572, w_011_065);
  or2  I013_278(w_013_278, w_006_022, w_005_089);
  or2  I013_279(w_013_279, w_005_293, w_004_121);
  nand2 I013_280(w_013_280, w_008_238, w_000_1172);
  nand2 I013_281(w_013_281, w_000_814, w_000_1119);
  nand2 I013_282(w_013_282, w_000_1184, w_002_239);
  nand2 I013_283(w_013_283, w_003_164, w_003_119);
  and2 I013_284(w_013_284, w_006_045, w_011_453);
  not1 I013_285(w_013_285, w_001_406);
  not1 I013_286(w_013_286, w_007_879);
  or2  I013_287(w_013_287, w_002_523, w_007_1349);
  and2 I013_288(w_013_288, w_007_515, w_004_078);
  not1 I013_289(w_013_289, w_006_153);
  and2 I013_290(w_013_290, w_012_180, w_002_333);
  not1 I013_291(w_013_291, w_007_915);
  or2  I013_292(w_013_292, w_005_574, w_011_344);
  not1 I013_293(w_013_293, w_006_026);
  nand2 I013_294(w_013_294, w_003_215, w_004_1641);
  and2 I013_295(w_013_295, w_008_110, w_001_432);
  or2  I013_296(w_013_296, w_011_022, w_004_1015);
  not1 I013_297(w_013_297, w_004_1863);
  and2 I013_298(w_013_298, w_004_1194, w_001_295);
  nand2 I013_299(w_013_299, w_006_189, w_006_135);
  nand2 I013_300(w_013_300, w_001_225, w_003_199);
  and2 I013_301(w_013_301, w_010_178, w_012_422);
  nand2 I013_302(w_013_302, w_002_190, w_009_007);
  or2  I013_303(w_013_303, w_000_1694, w_001_213);
  not1 I013_304(w_013_304, w_008_418);
  and2 I013_305(w_013_305, w_009_027, w_001_1387);
  nand2 I013_307(w_013_307, w_010_346, w_012_520);
  or2  I013_309(w_013_309, w_003_189, w_007_840);
  not1 I013_311(w_013_311, w_001_797);
  or2  I013_312(w_013_312, w_000_253, w_011_205);
  and2 I013_313(w_013_313, w_002_000, w_001_756);
  not1 I013_314(w_013_314, w_000_591);
  and2 I013_315(w_013_315, w_007_1507, w_004_159);
  not1 I013_316(w_013_316, w_006_096);
  and2 I013_318(w_013_318, w_004_190, w_009_056);
  nand2 I013_319(w_013_319, w_012_429, w_006_327);
  or2  I013_320(w_013_320, w_011_733, w_012_271);
  nand2 I013_321(w_013_321, w_001_862, w_010_027);
  and2 I013_323(w_013_323, w_003_182, w_006_283);
  not1 I013_324(w_013_324, w_001_374);
  and2 I013_325(w_013_325, w_000_1886, w_011_439);
  nand2 I013_326(w_013_326, w_006_086, w_005_504);
  and2 I013_327(w_013_327, w_006_095, w_007_025);
  not1 I013_328(w_013_328, w_006_182);
  not1 I013_330(w_013_330, w_009_008);
  nand2 I013_331(w_013_331, w_003_258, w_011_125);
  nand2 I013_332(w_013_332, w_000_363, w_002_114);
  not1 I013_335(w_013_335, w_007_756);
  not1 I013_336(w_013_336, w_005_1006);
  or2  I013_337(w_013_337, w_002_210, w_009_100);
  nand2 I013_338(w_013_338, w_002_146, w_003_036);
  nand2 I014_001(w_014_001, w_004_1694, w_009_105);
  and2 I014_002(w_014_002, w_007_699, w_002_023);
  and2 I014_003(w_014_003, w_006_139, w_001_518);
  not1 I014_005(w_014_005, w_012_278);
  and2 I014_008(w_014_008, w_008_085, w_005_1173);
  not1 I014_013(w_014_013, w_003_197);
  or2  I014_014(w_014_014, w_000_1370, w_005_109);
  nand2 I014_015(w_014_015, w_008_646, w_003_252);
  and2 I014_017(w_014_017, w_001_593, w_005_074);
  or2  I014_018(w_014_018, w_013_036, w_003_153);
  not1 I014_019(w_014_019, w_000_1304);
  and2 I014_020(w_014_020, w_001_173, w_007_384);
  nand2 I014_022(w_014_022, w_004_1301, w_012_580);
  not1 I014_023(w_014_023, w_008_188);
  nand2 I014_024(w_014_024, w_007_782, w_006_053);
  nand2 I014_025(w_014_025, w_003_153, w_006_240);
  not1 I014_027(w_014_027, w_005_611);
  nand2 I014_029(w_014_029, w_004_1040, w_003_262);
  nand2 I014_032(w_014_032, w_002_142, w_011_523);
  nand2 I014_038(w_014_038, w_007_921, w_003_159);
  or2  I014_040(w_014_040, w_011_378, w_006_080);
  not1 I014_041(w_014_041, w_002_103);
  nand2 I014_043(w_014_043, w_009_070, w_006_272);
  not1 I014_049(w_014_049, w_000_1910);
  nand2 I014_051(w_014_051, w_003_281, w_007_569);
  and2 I014_053(w_014_053, w_001_1111, w_008_088);
  or2  I014_055(w_014_055, w_007_342, w_013_205);
  not1 I014_056(w_014_056, w_011_164);
  nand2 I014_058(w_014_058, w_006_166, w_000_1885);
  or2  I014_059(w_014_059, w_000_504, w_007_517);
  and2 I014_060(w_014_060, w_001_605, w_004_1467);
  not1 I014_061(w_014_061, w_013_219);
  not1 I014_065(w_014_065, w_013_174);
  nand2 I014_070(w_014_070, w_011_228, w_009_057);
  not1 I014_072(w_014_072, w_002_258);
  and2 I014_074(w_014_074, w_008_518, w_011_752);
  nand2 I014_076(w_014_076, w_011_062, w_010_268);
  not1 I014_077(w_014_077, w_002_183);
  and2 I014_078(w_014_078, w_008_258, w_013_307);
  nand2 I014_079(w_014_079, w_008_660, w_011_128);
  nand2 I014_080(w_014_080, w_008_195, w_011_596);
  and2 I014_082(w_014_082, w_009_075, w_008_164);
  and2 I014_084(w_014_084, w_002_002, w_009_005);
  or2  I014_085(w_014_085, w_004_211, w_006_151);
  nand2 I014_086(w_014_086, w_005_322, w_001_1660);
  not1 I014_087(w_014_087, w_011_094);
  nand2 I014_089(w_014_089, w_001_017, w_012_305);
  nand2 I014_090(w_014_090, w_012_627, w_005_732);
  not1 I014_091(w_014_091, w_012_406);
  nand2 I014_092(w_014_092, w_002_097, w_006_056);
  or2  I014_093(w_014_093, w_009_093, w_008_379);
  nand2 I014_094(w_014_094, w_003_254, w_004_664);
  or2  I014_097(w_014_097, w_002_316, w_010_353);
  not1 I014_099(w_014_099, w_012_551);
  and2 I014_101(w_014_101, w_002_198, w_003_300);
  not1 I014_102(w_014_102, w_013_107);
  or2  I014_104(w_014_104, w_006_240, w_002_041);
  nand2 I014_106(w_014_106, w_010_188, w_008_172);
  or2  I014_107(w_014_107, w_008_199, w_009_024);
  or2  I014_108(w_014_108, w_012_509, w_012_181);
  and2 I014_109(w_014_109, w_012_560, w_002_546);
  or2  I014_110(w_014_110, w_006_134, w_001_1300);
  not1 I014_112(w_014_112, w_004_1865);
  and2 I014_115(w_014_115, w_010_316, w_010_371);
  and2 I014_116(w_014_116, w_006_197, w_000_1678);
  not1 I014_117(w_014_117, w_002_067);
  and2 I014_118(w_014_118, w_008_208, w_008_124);
  nand2 I014_119(w_014_119, w_011_389, w_005_650);
  not1 I014_121(w_014_121, w_003_110);
  nand2 I014_123(w_014_123, w_008_527, w_000_354);
  or2  I014_124(w_014_124, w_010_227, w_013_172);
  and2 I014_125(w_014_125, w_008_144, w_006_331);
  and2 I014_129(w_014_129, w_004_1786, w_001_291);
  and2 I014_130(w_014_130, w_002_349, w_004_151);
  or2  I014_131(w_014_131, w_000_098, w_009_090);
  or2  I014_132(w_014_132, w_007_085, w_008_474);
  or2  I014_133(w_014_133, w_006_257, w_010_217);
  not1 I014_136(w_014_136, w_006_123);
  or2  I014_138(w_014_138, w_011_125, w_012_490);
  and2 I014_140(w_014_140, w_008_231, w_012_061);
  or2  I014_142(w_014_142, w_005_1422, w_011_232);
  and2 I014_143(w_014_143, w_012_526, w_011_551);
  or2  I014_144(w_014_144, w_003_210, w_013_098);
  nand2 I014_145(w_014_145, w_010_127, w_002_300);
  not1 I014_147(w_014_147, w_011_188);
  nand2 I014_149(w_014_149, w_001_444, w_002_089);
  nand2 I014_150(w_014_150, w_011_350, w_006_090);
  or2  I014_151(w_014_151, w_006_184, w_008_436);
  not1 I014_154(w_014_154, w_002_246);
  nand2 I014_156(w_014_156, w_011_420, w_006_074);
  not1 I014_157(w_014_157, w_010_277);
  nand2 I014_158(w_014_158, w_000_1445, w_012_445);
  and2 I014_159(w_014_159, w_004_202, w_009_025);
  nand2 I014_160(w_014_160, w_008_683, w_013_136);
  or2  I014_161(w_014_161, w_013_210, w_001_397);
  not1 I014_163(w_014_163, w_012_453);
  and2 I014_164(w_014_164, w_006_305, w_000_1765);
  not1 I014_165(w_014_165, w_010_388);
  nand2 I014_167(w_014_167, w_012_143, w_006_176);
  or2  I014_168(w_014_168, w_003_123, w_012_618);
  and2 I014_169(w_014_169, w_006_088, w_002_509);
  nand2 I014_171(w_014_171, w_004_331, w_001_189);
  not1 I014_172(w_014_172, w_009_101);
  or2  I014_177(w_014_177, w_009_106, w_009_077);
  or2  I014_178(w_014_178, w_000_1208, w_000_1885);
  not1 I014_179(w_014_179, w_009_099);
  or2  I014_181(w_014_181, w_005_191, w_013_141);
  and2 I014_184(w_014_184, w_005_1663, w_007_183);
  not1 I014_189(w_014_189, w_007_295);
  or2  I014_191(w_014_191, w_003_066, w_005_1587);
  nand2 I014_193(w_014_193, w_011_036, w_012_221);
  not1 I014_194(w_014_194, w_007_704);
  not1 I014_195(w_014_195, w_009_053);
  and2 I014_196(w_014_196, w_000_972, w_013_229);
  and2 I014_197(w_014_197, w_002_175, w_008_527);
  and2 I014_199(w_014_199, w_002_194, w_007_158);
  not1 I014_203(w_014_203, w_011_142);
  not1 I014_204(w_014_204, w_011_741);
  not1 I014_205(w_014_205, w_008_437);
  and2 I014_208(w_014_208, w_000_517, w_005_1002);
  or2  I014_209(w_014_209, w_010_324, w_013_299);
  nand2 I014_210(w_014_210, w_009_058, w_001_669);
  or2  I014_211(w_014_211, w_007_095, w_003_030);
  or2  I014_212(w_014_212, w_009_067, w_007_147);
  or2  I014_213(w_014_213, w_009_066, w_004_1652);
  or2  I014_214(w_014_214, w_000_1436, w_000_1551);
  or2  I014_218(w_014_218, w_001_1397, w_012_451);
  or2  I014_219(w_014_219, w_005_890, w_006_165);
  or2  I014_221(w_014_221, w_003_110, w_009_018);
  and2 I014_223(w_014_223, w_000_075, w_005_709);
  not1 I014_225(w_014_225, w_008_442);
  nand2 I014_226(w_014_226, w_013_324, w_009_040);
  or2  I014_229(w_014_229, w_006_087, w_013_255);
  nand2 I014_232(w_014_232, w_006_279, w_008_612);
  not1 I014_234(w_014_234, w_001_1655);
  and2 I014_235(w_014_235, w_001_916, w_008_729);
  and2 I014_237(w_014_237, w_011_850, w_013_031);
  nand2 I014_239(w_014_239, w_009_052, w_007_313);
  nand2 I014_242(w_014_242, w_009_074, w_005_973);
  nand2 I014_243(w_014_243, w_003_234, w_003_224);
  nand2 I014_246(w_014_246, w_012_133, w_008_306);
  or2  I014_247(w_014_247, w_001_059, w_012_654);
  not1 I014_248(w_014_248, w_000_1807);
  or2  I014_249(w_014_249, w_005_1132, w_006_080);
  and2 I014_251(w_014_251, w_007_1351, w_009_083);
  nand2 I014_252(w_014_252, w_006_200, w_004_1463);
  or2  I014_255(w_014_255, w_009_030, w_004_340);
  not1 I014_256(w_014_256, w_008_148);
  and2 I014_257(w_014_257, w_002_240, w_002_335);
  and2 I014_258(w_014_258, w_012_662, w_001_116);
  nand2 I014_261(w_014_261, w_010_357, w_012_537);
  and2 I014_262(w_014_262, w_000_1230, w_004_321);
  not1 I014_263(w_014_263, w_003_017);
  nand2 I014_264(w_014_264, w_005_1025, w_001_1673);
  or2  I014_266(w_014_266, w_013_059, w_003_291);
  or2  I014_268(w_014_268, w_010_175, w_006_159);
  or2  I014_270(w_014_270, w_008_154, w_004_1641);
  and2 I014_271(w_014_271, w_008_038, w_004_1212);
  nand2 I014_272(w_014_272, w_004_213, w_006_189);
  or2  I014_273(w_014_273, w_001_502, w_002_049);
  and2 I014_274(w_014_274, w_001_1167, w_005_1171);
  not1 I014_276(w_014_276, w_001_143);
  and2 I014_277(w_014_277, w_008_297, w_008_038);
  nand2 I014_278(w_014_278, w_002_025, w_003_229);
  not1 I014_279(w_014_279, w_005_079);
  and2 I014_280(w_014_280, w_008_674, w_011_721);
  not1 I014_286(w_014_286, w_012_073);
  not1 I014_288(w_014_288, w_008_031);
  not1 I014_290(w_014_290, w_013_233);
  not1 I014_291(w_014_291, w_002_536);
  or2  I014_293(w_014_293, w_008_346, w_004_404);
  or2  I014_295(w_014_295, w_005_1121, w_000_1221);
  or2  I014_296(w_014_296, w_012_094, w_012_596);
  not1 I014_299(w_014_299, w_012_477);
  or2  I014_300(w_014_300, w_002_119, w_004_540);
  and2 I014_304(w_014_304, w_006_165, w_013_294);
  and2 I014_308(w_014_308, w_008_847, w_011_386);
  nand2 I014_309(w_014_309, w_009_080, w_001_929);
  nand2 I014_310(w_014_310, w_010_180, w_003_273);
  nand2 I014_311(w_014_311, w_002_579, w_001_240);
  nand2 I014_312(w_014_312, w_013_260, w_005_570);
  nand2 I014_313(w_014_313, w_010_036, w_003_276);
  and2 I014_314(w_014_314, w_012_262, w_000_1561);
  and2 I014_315(w_014_315, w_005_1557, w_000_531);
  not1 I014_316(w_014_316, w_001_1183);
  nand2 I014_318(w_014_318, w_007_808, w_013_250);
  and2 I014_319(w_014_319, w_004_1161, w_001_280);
  or2  I014_320(w_014_320, w_003_236, w_005_036);
  not1 I014_321(w_014_321, w_004_1624);
  not1 I014_322(w_014_322, w_009_061);
  not1 I014_323(w_014_323, w_000_020);
  not1 I014_324(w_014_324, w_012_545);
  nand2 I014_326(w_014_326, w_010_037, w_001_1637);
  nand2 I014_327(w_014_327, w_000_1312, w_009_092);
  nand2 I014_329(w_014_329, w_009_019, w_013_294);
  or2  I014_330(w_014_330, w_011_314, w_001_147);
  or2  I014_333(w_014_333, w_007_586, w_010_160);
  nand2 I014_334(w_014_334, w_003_288, w_006_030);
  or2  I014_335(w_014_335, w_011_623, w_009_006);
  nand2 I014_337(w_014_337, w_005_535, w_011_417);
  not1 I014_340(w_014_340, w_009_068);
  not1 I014_341(w_014_341, w_001_991);
  or2  I014_342(w_014_342, w_005_316, w_003_294);
  or2  I014_344(w_014_344, w_005_271, w_001_1458);
  not1 I014_345(w_014_345, w_002_299);
  not1 I014_349(w_014_349, w_002_079);
  and2 I014_352(w_014_352, w_013_327, w_010_178);
  or2  I014_353(w_014_353, w_005_077, w_012_040);
  not1 I014_359(w_014_359, w_003_249);
  and2 I014_360(w_014_360, w_007_1601, w_006_281);
  nand2 I014_361(w_014_361, w_007_477, w_004_375);
  not1 I014_362(w_014_362, w_000_1514);
  or2  I014_365(w_014_365, w_006_050, w_012_053);
  and2 I014_366(w_014_366, w_000_1238, w_012_007);
  not1 I014_370(w_014_370, w_012_377);
  not1 I014_372(w_014_372, w_009_063);
  or2  I014_375(w_014_375, w_012_042, w_012_191);
  or2  I014_376(w_014_376, w_006_322, w_000_1912);
  and2 I014_380(w_014_380, w_009_072, w_010_044);
  and2 I014_383(w_014_383, w_004_591, w_008_668);
  not1 I014_384(w_014_384, w_011_177);
  and2 I014_385(w_014_385, w_009_036, w_009_095);
  not1 I014_387(w_014_387, w_010_220);
  nand2 I014_390(w_014_390, w_009_047, w_010_012);
  nand2 I014_392(w_014_392, w_000_842, w_007_598);
  nand2 I014_393(w_014_393, w_008_238, w_003_076);
  nand2 I014_397(w_014_397, w_003_129, w_012_206);
  nand2 I014_398(w_014_398, w_013_245, w_011_836);
  not1 I014_402(w_014_402, w_009_035);
  or2  I014_403(w_014_403, w_004_894, w_008_579);
  nand2 I014_405(w_014_405, w_006_100, w_004_697);
  and2 I014_406(w_014_406, w_001_408, w_007_1510);
  not1 I014_411(w_014_411, w_005_907);
  or2  I014_412(w_014_412, w_010_011, w_003_053);
  not1 I014_416(w_014_416, w_004_848);
  nand2 I014_417(w_014_417, w_006_265, w_012_218);
  nand2 I014_420(w_014_420, w_011_588, w_009_111);
  not1 I014_422(w_014_422, w_007_654);
  nand2 I014_426(w_014_426, w_009_101, w_011_148);
  or2  I014_427(w_014_427, w_004_1719, w_000_1403);
  or2  I014_430(w_014_430, w_006_130, w_006_020);
  and2 I014_432(w_014_432, w_006_262, w_001_1121);
  and2 I014_433(w_014_433, w_010_084, w_011_738);
  or2  I014_434(w_014_434, w_011_493, w_008_807);
  and2 I014_436(w_014_436, w_005_1428, w_007_485);
  and2 I014_437(w_014_437, w_004_1839, w_010_012);
  not1 I014_438(w_014_438, w_000_152);
  or2  I014_439(w_014_439, w_013_254, w_007_102);
  nand2 I014_442(w_014_442, w_013_105, w_003_070);
  or2  I014_443(w_014_443, w_006_074, w_012_494);
  not1 I014_445(w_014_445, w_008_819);
  not1 I014_447(w_014_447, w_005_049);
  or2  I014_451(w_014_451, w_007_106, w_002_200);
  or2  I014_453(w_014_453, w_006_163, w_006_001);
  or2  I014_454(w_014_454, w_011_394, w_011_019);
  or2  I014_457(w_014_457, w_007_948, w_009_005);
  not1 I014_459(w_014_459, w_005_1175);
  not1 I014_461(w_014_461, w_004_507);
  and2 I014_465(w_014_465, w_004_1744, w_013_009);
  or2  I014_467(w_014_467, w_003_305, w_006_233);
  not1 I014_469(w_014_469, w_012_201);
  or2  I014_470(w_014_470, w_007_351, w_006_111);
  not1 I014_473(w_014_473, w_004_949);
  not1 I014_475(w_014_475, w_005_1596);
  nand2 I014_477(w_014_477, w_006_094, w_003_014);
  nand2 I014_478(w_014_478, w_012_227, w_013_022);
  not1 I014_481(w_014_481, w_009_028);
  not1 I014_483(w_014_483, w_006_209);
  nand2 I014_486(w_014_486, w_009_100, w_004_236);
  or2  I014_487(w_014_487, w_004_1865, w_013_106);
  nand2 I014_489(w_014_489, w_002_040, w_011_114);
  or2  I014_491(w_014_491, w_001_1633, w_013_184);
  and2 I014_492(w_014_492, w_008_102, w_007_953);
  or2  I014_495(w_014_495, w_008_315, w_012_174);
  or2  I014_500(w_014_500, w_003_097, w_005_400);
  and2 I014_502(w_014_502, w_010_103, w_010_331);
  nand2 I014_504(w_014_504, w_001_362, w_001_329);
  nand2 I014_505(w_014_505, w_013_063, w_003_025);
  or2  I014_506(w_014_506, w_006_119, w_003_047);
  nand2 I014_508(w_014_508, w_010_116, w_009_010);
  not1 I014_509(w_014_509, w_001_1568);
  and2 I014_512(w_014_512, w_012_153, w_007_208);
  and2 I014_516(w_014_516, w_009_046, w_006_291);
  and2 I014_517(w_014_517, w_010_129, w_000_970);
  nand2 I014_518(w_014_518, w_007_1446, w_001_427);
  nand2 I014_519(w_014_519, w_008_123, w_003_085);
  and2 I014_520(w_014_520, w_003_298, w_004_517);
  not1 I014_523(w_014_523, w_001_163);
  and2 I014_524(w_014_524, w_013_155, w_005_033);
  or2  I014_525(w_014_525, w_004_487, w_012_659);
  nand2 I014_526(w_014_526, w_001_022, w_001_1402);
  or2  I014_528(w_014_528, w_006_328, w_003_107);
  nand2 I014_529(w_014_529, w_000_070, w_006_268);
  not1 I014_532(w_014_532, w_005_577);
  or2  I014_533(w_014_533, w_006_289, w_003_289);
  nand2 I014_534(w_014_534, w_006_088, w_005_915);
  and2 I014_537(w_014_537, w_005_1093, w_007_657);
  not1 I014_540(w_014_540, w_010_147);
  not1 I014_543(w_014_543, w_001_143);
  nand2 I014_544(w_014_544, w_010_254, w_002_231);
  nand2 I014_545(w_014_545, w_005_137, w_003_128);
  or2  I014_547(w_014_547, w_013_088, w_005_790);
  and2 I014_551(w_014_551, w_005_713, w_006_240);
  and2 I014_556(w_014_556, w_003_130, w_008_421);
  or2  I014_560(w_014_560, w_002_389, w_006_139);
  not1 I014_561(w_014_561, w_012_059);
  or2  I014_565(w_014_565, w_002_530, w_010_379);
  nand2 I014_567(w_014_567, w_001_261, w_004_898);
  nand2 I014_569(w_014_569, w_012_475, w_008_098);
  nand2 I014_573(w_014_573, w_001_520, w_004_1169);
  nand2 I014_574(w_014_574, w_004_1472, w_011_738);
  and2 I014_576(w_014_576, w_002_434, w_009_076);
  not1 I014_577(w_014_577, w_006_111);
  and2 I014_578(w_014_578, w_012_375, w_009_071);
  not1 I014_579(w_014_579, w_002_559);
  not1 I014_581(w_014_581, w_009_046);
  and2 I014_582(w_014_582, w_011_037, w_000_424);
  nand2 I014_583(w_014_583, w_009_017, w_003_277);
  not1 I014_586(w_014_586, w_012_195);
  or2  I014_588(w_014_588, w_009_024, w_006_307);
  and2 I014_590(w_014_590, w_000_324, w_000_1913);
  or2  I014_598(w_014_598, w_003_202, w_009_073);
  nand2 I014_599(w_014_599, w_004_1907, w_002_136);
  not1 I014_601(w_014_601, w_009_023);
  or2  I014_604(w_014_604, w_003_178, w_000_1526);
  not1 I014_606(w_014_606, w_010_279);
  not1 I014_607(w_014_607, w_001_1502);
  not1 I014_609(w_014_609, w_002_169);
  or2  I014_611(w_014_611, w_011_262, w_000_069);
  not1 I014_613(w_014_613, w_010_278);
  or2  I014_614(w_014_614, w_004_1573, w_012_170);
  not1 I014_617(w_014_617, w_006_183);
  not1 I014_619(w_014_619, w_005_979);
  and2 I014_623(w_014_623, w_011_819, w_003_086);
  and2 I014_624(w_014_624, w_005_628, w_005_1588);
  not1 I014_626(w_014_626, w_010_190);
  or2  I014_629(w_014_629, w_007_1402, w_003_269);
  or2  I014_632(w_014_632, w_009_065, w_011_079);
  or2  I014_636(w_014_636, w_006_269, w_005_534);
  or2  I014_639(w_014_639, w_002_025, w_011_755);
  not1 I014_640(w_014_640, w_002_113);
  not1 I014_641(w_014_641, w_010_247);
  and2 I014_643(w_014_643, w_013_167, w_009_077);
  not1 I014_644(w_014_644, w_011_559);
  and2 I014_646(w_014_646, w_013_067, w_006_056);
  and2 I014_648(w_014_648, w_002_264, w_006_111);
  and2 I014_649(w_014_649, w_007_418, w_005_025);
  not1 I014_650(w_014_650, w_002_192);
  or2  I014_651(w_014_651, w_001_663, w_005_154);
  not1 I014_652(w_014_652, w_006_281);
  and2 I014_653(w_014_653, w_005_533, w_005_1132);
  nand2 I014_654(w_014_654, w_007_894, w_004_209);
  nand2 I014_659(w_014_659, w_000_1177, w_003_266);
  nand2 I014_661(w_014_661, w_001_1568, w_013_185);
  nand2 I014_662(w_014_662, w_004_1679, w_012_328);
  or2  I014_663(w_014_663, w_007_1198, w_006_104);
  nand2 I014_664(w_014_664, w_009_084, w_004_139);
  or2  I014_666(w_014_666, w_008_678, w_001_1571);
  nand2 I014_668(w_014_668, w_008_694, w_004_313);
  or2  I014_672(w_014_672, w_003_002, w_010_080);
  and2 I014_673(w_014_673, w_009_061, w_009_019);
  and2 I014_677(w_014_677, w_002_047, w_011_573);
  not1 I014_685(w_014_685, w_011_216);
  nand2 I014_686(w_014_686, w_006_272, w_005_769);
  or2  I014_688(w_014_688, w_011_464, w_000_1916);
  and2 I014_690(w_014_690, w_009_105, w_000_080);
  or2  I014_691(w_014_691, w_005_730, w_009_006);
  not1 I014_692(w_014_692, w_006_116);
  or2  I014_696(w_014_696, w_012_505, w_000_1917);
  nand2 I014_702(w_014_702, w_000_1222, w_006_225);
  nand2 I014_703(w_014_703, w_006_172, w_005_857);
  and2 I014_704(w_014_704, w_011_163, w_005_932);
  and2 I014_707(w_014_707, w_011_782, w_001_273);
  or2  I014_708(w_014_708, w_002_131, w_005_1364);
  not1 I014_709(w_014_709, w_005_1348);
  not1 I014_711(w_014_711, w_005_369);
  and2 I014_713(w_014_713, w_010_369, w_003_045);
  not1 I014_716(w_014_716, w_006_055);
  or2  I014_717(w_014_717, w_001_1314, w_011_407);
  not1 I014_719(w_014_719, w_011_490);
  and2 I014_721(w_014_721, w_011_203, w_008_003);
  and2 I014_722(w_014_722, w_002_082, w_007_289);
  not1 I014_723(w_014_723, w_010_244);
  nand2 I014_726(w_014_726, w_003_319, w_000_809);
  or2  I014_728(w_014_728, w_006_160, w_000_576);
  and2 I014_729(w_014_729, w_009_032, w_006_148);
  not1 I014_732(w_014_732, w_006_044);
  or2  I014_734(w_014_734, w_004_1753, w_011_328);
  and2 I014_736(w_014_736, w_001_423, w_002_550);
  and2 I014_738(w_014_738, w_002_100, w_006_197);
  not1 I014_740(w_014_740, w_001_806);
  not1 I014_745(w_014_745, w_005_1582);
  or2  I014_746(w_014_746, w_010_098, w_008_408);
  and2 I014_752(w_014_752, w_012_212, w_001_182);
  or2  I014_755(w_014_755, w_009_027, w_006_117);
  not1 I014_757(w_014_757, w_000_365);
  or2  I014_767(w_014_767, w_008_059, w_012_425);
  or2  I014_768(w_014_768, w_000_1494, w_006_110);
  or2  I014_772(w_014_772, w_011_347, w_003_076);
  not1 I014_777(w_014_777, w_005_156);
  nand2 I014_780(w_014_780, w_010_126, w_006_226);
  not1 I014_784(w_014_784, w_004_764);
  not1 I014_787(w_014_787, w_006_162);
  nand2 I014_793(w_014_793, w_012_202, w_005_741);
  not1 I014_795(w_014_795, w_002_216);
  nand2 I014_796(w_014_796, w_004_207, w_002_187);
  and2 I014_798(w_014_798, w_010_055, w_001_1437);
  or2  I014_801(w_014_801, w_010_322, w_013_303);
  not1 I014_805(w_014_805, w_005_897);
  or2  I014_806(w_014_806, w_006_174, w_009_013);
  or2  I014_807(w_014_807, w_003_131, w_001_674);
  and2 I014_808(w_014_808, w_009_079, w_008_070);
  nand2 I014_809(w_014_809, w_011_687, w_005_434);
  or2  I014_810(w_014_810, w_003_062, w_011_480);
  or2  I014_814(w_014_814, w_009_089, w_000_1907);
  and2 I014_815(w_014_815, w_008_059, w_004_1549);
  or2  I014_819(w_014_819, w_006_193, w_007_673);
  or2  I014_821(w_014_821, w_004_361, w_013_018);
  not1 I014_822(w_014_822, w_006_225);
  or2  I014_823(w_014_823, w_004_1228, w_006_214);
  nand2 I014_824(w_014_824, w_007_884, w_010_116);
  nand2 I014_825(w_014_825, w_011_532, w_010_312);
  or2  I014_826(w_014_826, w_004_1021, w_001_445);
  and2 I014_829(w_014_829, w_012_446, w_006_330);
  and2 I014_830(w_014_830, w_011_879, w_012_641);
  not1 I014_831(w_014_831, w_010_369);
  and2 I015_000(w_015_000, w_010_059, w_008_008);
  and2 I015_001(w_015_001, w_005_1553, w_001_1185);
  not1 I015_002(w_015_002, w_011_154);
  and2 I015_003(w_015_003, w_010_311, w_009_077);
  or2  I015_004(w_015_004, w_001_1557, w_009_101);
  and2 I015_005(w_015_005, w_007_138, w_007_761);
  not1 I015_006(w_015_006, w_003_079);
  not1 I015_007(w_015_007, w_013_098);
  nand2 I015_008(w_015_008, w_013_170, w_007_483);
  not1 I015_010(w_015_010, w_010_032);
  or2  I015_011(w_015_011, w_003_099, w_001_1532);
  nand2 I015_012(w_015_012, w_014_793, w_006_301);
  nand2 I015_013(w_015_013, w_009_079, w_012_184);
  not1 I015_014(w_015_014, w_002_126);
  or2  I015_015(w_015_015, w_007_517, w_002_567);
  not1 I015_016(w_015_016, w_012_345);
  not1 I015_017(w_015_017, w_011_324);
  nand2 I015_019(w_015_019, w_009_005, w_008_139);
  and2 I015_020(w_015_020, w_008_735, w_002_027);
  or2  I015_021(w_015_021, w_013_045, w_011_051);
  not1 I015_022(w_015_022, w_003_172);
  and2 I015_023(w_015_023, w_010_357, w_010_061);
  and2 I015_024(w_015_024, w_013_288, w_000_425);
  or2  I015_025(w_015_025, w_002_327, w_003_281);
  and2 I015_026(w_015_026, w_011_353, w_005_039);
  and2 I015_027(w_015_027, w_014_078, w_013_173);
  or2  I015_030(w_015_030, w_001_1637, w_005_146);
  not1 I015_031(w_015_031, w_006_331);
  or2  I015_032(w_015_032, w_009_012, w_003_093);
  or2  I015_033(w_015_033, w_000_799, w_001_1390);
  or2  I015_034(w_015_034, w_014_239, w_003_010);
  nand2 I015_035(w_015_035, w_003_041, w_000_101);
  nand2 I015_036(w_015_036, w_000_474, w_008_151);
  and2 I015_038(w_015_038, w_012_139, w_010_411);
  and2 I015_039(w_015_039, w_008_533, w_006_203);
  and2 I015_040(w_015_040, w_012_330, w_013_290);
  and2 I015_041(w_015_041, w_011_705, w_013_053);
  not1 I015_042(w_015_042, w_001_1390);
  and2 I015_043(w_015_043, w_001_203, w_006_327);
  not1 I015_044(w_015_044, w_012_328);
  not1 I015_045(w_015_045, w_001_1487);
  not1 I015_046(w_015_046, w_001_1379);
  and2 I015_047(w_015_047, w_010_001, w_014_385);
  nand2 I015_048(w_015_048, w_007_157, w_011_838);
  nand2 I015_049(w_015_049, w_006_092, w_008_224);
  or2  I015_050(w_015_050, w_010_242, w_008_569);
  or2  I015_052(w_015_052, w_003_277, w_002_421);
  and2 I015_053(w_015_053, w_000_612, w_011_816);
  and2 I015_055(w_015_055, w_007_874, w_004_1647);
  nand2 I015_056(w_015_056, w_002_080, w_011_189);
  nand2 I015_057(w_015_057, w_009_100, w_004_1836);
  not1 I015_058(w_015_058, w_002_410);
  and2 I015_059(w_015_059, w_005_371, w_014_023);
  nand2 I015_060(w_015_060, w_002_503, w_005_1022);
  or2  I015_061(w_015_061, w_007_478, w_013_201);
  and2 I015_062(w_015_062, w_002_286, w_003_205);
  not1 I015_064(w_015_064, w_005_504);
  or2  I015_065(w_015_065, w_007_237, w_006_127);
  and2 I015_066(w_015_066, w_012_478, w_003_097);
  or2  I015_067(w_015_067, w_008_719, w_012_104);
  or2  I015_068(w_015_068, w_011_006, w_013_030);
  not1 I015_069(w_015_069, w_002_039);
  or2  I015_070(w_015_070, w_008_382, w_012_169);
  and2 I015_071(w_015_071, w_002_505, w_014_677);
  nand2 I015_073(w_015_073, w_010_155, w_012_441);
  or2  I015_074(w_015_074, w_012_180, w_009_092);
  or2  I015_075(w_015_075, w_012_106, w_000_1238);
  or2  I015_076(w_015_076, w_009_017, w_002_228);
  nand2 I015_077(w_015_077, w_006_033, w_011_543);
  not1 I015_078(w_015_078, w_002_405);
  or2  I015_079(w_015_079, w_000_746, w_014_160);
  or2  I015_080(w_015_080, w_003_161, w_013_167);
  or2  I015_081(w_015_081, w_008_098, w_001_045);
  not1 I015_082(w_015_082, w_008_770);
  nand2 I015_083(w_015_083, w_003_133, w_006_312);
  and2 I015_084(w_015_084, w_013_073, w_000_523);
  not1 I015_086(w_015_086, w_001_914);
  and2 I015_087(w_015_087, w_011_035, w_001_098);
  and2 I015_088(w_015_088, w_001_1062, w_014_242);
  and2 I015_089(w_015_089, w_007_253, w_009_110);
  not1 I015_090(w_015_090, w_000_878);
  nand2 I015_091(w_015_091, w_005_1303, w_010_324);
  nand2 I015_093(w_015_093, w_013_273, w_001_1319);
  and2 I015_094(w_015_094, w_009_074, w_001_466);
  not1 I015_097(w_015_097, w_002_236);
  and2 I015_099(w_015_099, w_012_239, w_006_304);
  or2  I015_100(w_015_100, w_014_311, w_008_384);
  or2  I015_101(w_015_101, w_002_014, w_006_024);
  nand2 I015_103(w_015_103, w_003_137, w_008_264);
  nand2 I015_104(w_015_104, w_010_010, w_005_262);
  and2 I015_105(w_015_105, w_013_149, w_012_249);
  and2 I015_106(w_015_106, w_011_141, w_000_1921);
  and2 I015_108(w_015_108, w_008_857, w_007_781);
  or2  I015_110(w_015_110, w_011_112, w_002_363);
  or2  I015_112(w_015_112, w_008_662, w_012_580);
  and2 I015_113(w_015_113, w_013_107, w_006_205);
  or2  I015_115(w_015_115, w_001_1152, w_013_160);
  or2  I015_116(w_015_116, w_008_213, w_005_538);
  nand2 I015_117(w_015_117, w_009_043, w_008_144);
  or2  I015_118(w_015_118, w_002_247, w_004_1319);
  nand2 I015_119(w_015_119, w_006_262, w_003_259);
  nand2 I015_120(w_015_120, w_000_1782, w_004_819);
  and2 I015_122(w_015_122, w_009_009, w_002_417);
  not1 I015_124(w_015_124, w_013_103);
  or2  I015_125(w_015_125, w_009_019, w_007_1615);
  or2  I015_126(w_015_126, w_002_560, w_013_124);
  or2  I015_127(w_015_127, w_002_096, w_007_1094);
  and2 I015_128(w_015_128, w_000_1667, w_000_1316);
  and2 I015_129(w_015_129, w_009_007, w_012_399);
  or2  I015_130(w_015_130, w_004_1270, w_007_1377);
  or2  I015_131(w_015_131, w_006_081, w_005_926);
  or2  I015_133(w_015_133, w_000_824, w_007_037);
  not1 I015_134(w_015_134, w_014_239);
  or2  I015_135(w_015_135, w_006_187, w_005_131);
  nand2 I015_136(w_015_136, w_009_085, w_014_074);
  nand2 I015_137(w_015_137, w_006_083, w_009_082);
  and2 I015_138(w_015_138, w_014_576, w_002_323);
  not1 I015_140(w_015_140, w_013_225);
  or2  I015_141(w_015_141, w_004_817, w_000_481);
  and2 I015_142(w_015_142, w_013_287, w_001_452);
  and2 I015_143(w_015_143, w_008_013, w_004_1204);
  not1 I015_144(w_015_144, w_013_174);
  nand2 I015_146(w_015_146, w_011_039, w_009_104);
  and2 I015_147(w_015_147, w_012_635, w_002_065);
  not1 I015_149(w_015_149, w_006_266);
  not1 I015_150(w_015_150, w_006_167);
  not1 I015_151(w_015_151, w_004_1511);
  not1 I015_152(w_015_152, w_003_164);
  or2  I015_153(w_015_153, w_000_1218, w_000_901);
  and2 I015_154(w_015_154, w_004_553, w_003_183);
  and2 I015_155(w_015_155, w_011_102, w_012_056);
  or2  I015_157(w_015_157, w_008_759, w_003_277);
  not1 I015_158(w_015_158, w_014_556);
  and2 I015_159(w_015_159, w_010_342, w_000_1655);
  nand2 I015_160(w_015_160, w_001_908, w_008_110);
  or2  I015_161(w_015_161, w_011_626, w_014_784);
  and2 I015_162(w_015_162, w_011_176, w_000_355);
  nand2 I015_163(w_015_163, w_010_357, w_006_015);
  or2  I015_164(w_015_164, w_001_203, w_014_685);
  or2  I015_165(w_015_165, w_013_242, w_010_286);
  or2  I015_166(w_015_166, w_000_782, w_013_188);
  or2  I015_168(w_015_168, w_009_049, w_000_869);
  and2 I015_169(w_015_169, w_002_338, w_008_688);
  not1 I015_170(w_015_170, w_011_141);
  nand2 I015_171(w_015_171, w_002_590, w_010_229);
  or2  I015_172(w_015_172, w_005_1041, w_000_867);
  nand2 I015_173(w_015_173, w_013_076, w_010_156);
  or2  I015_174(w_015_174, w_005_025, w_013_141);
  not1 I015_176(w_015_176, w_007_589);
  nand2 I015_177(w_015_177, w_000_483, w_011_787);
  not1 I015_178(w_015_178, w_013_090);
  or2  I015_181(w_015_181, w_001_1346, w_002_009);
  and2 I015_183(w_015_183, w_002_566, w_002_317);
  nand2 I015_184(w_015_184, w_005_1528, w_009_024);
  not1 I015_185(w_015_185, w_012_459);
  or2  I015_186(w_015_186, w_012_035, w_009_107);
  nand2 I015_187(w_015_187, w_005_1404, w_012_003);
  not1 I015_188(w_015_188, w_006_262);
  nand2 I015_189(w_015_189, w_007_436, w_012_236);
  or2  I015_190(w_015_190, w_014_732, w_004_379);
  and2 I015_191(w_015_191, w_009_036, w_007_126);
  not1 I015_192(w_015_192, w_011_209);
  and2 I015_193(w_015_193, w_008_400, w_000_337);
  and2 I015_194(w_015_194, w_005_066, w_010_012);
  and2 I015_195(w_015_195, w_008_151, w_011_293);
  not1 I015_196(w_015_196, w_008_750);
  not1 I015_198(w_015_198, w_012_105);
  and2 I015_199(w_015_199, w_010_189, w_005_151);
  nand2 I015_200(w_015_200, w_014_611, w_007_738);
  and2 I015_201(w_015_201, w_004_831, w_013_169);
  or2  I015_203(w_015_203, w_003_296, w_000_143);
  not1 I015_204(w_015_204, w_003_076);
  or2  I015_205(w_015_205, w_000_1117, w_007_1247);
  and2 I015_206(w_015_206, w_013_054, w_003_102);
  or2  I015_207(w_015_207, w_002_324, w_005_1577);
  nand2 I015_208(w_015_208, w_003_178, w_006_263);
  or2  I015_209(w_015_209, w_009_025, w_001_535);
  or2  I015_210(w_015_210, w_001_1030, w_001_274);
  not1 I015_211(w_015_211, w_014_257);
  nand2 I015_212(w_015_212, w_007_1504, w_000_1495);
  not1 I015_213(w_015_213, w_010_269);
  and2 I015_214(w_015_214, w_013_081, w_003_267);
  nand2 I015_216(w_015_216, w_014_204, w_013_236);
  or2  I015_217(w_015_217, w_007_1606, w_001_048);
  and2 I015_218(w_015_218, w_001_305, w_012_579);
  and2 I015_219(w_015_219, w_004_1410, w_010_040);
  nand2 I015_220(w_015_220, w_008_707, w_014_252);
  nand2 I015_221(w_015_221, w_005_560, w_004_192);
  nand2 I015_222(w_015_222, w_008_151, w_012_169);
  or2  I015_223(w_015_223, w_004_1633, w_000_732);
  nand2 I015_224(w_015_224, w_007_1173, w_002_378);
  and2 I015_225(w_015_225, w_009_088, w_010_386);
  not1 I015_226(w_015_226, w_001_190);
  not1 I015_227(w_015_227, w_007_1316);
  or2  I015_228(w_015_228, w_005_201, w_009_022);
  nand2 I015_229(w_015_229, w_009_031, w_011_846);
  and2 I015_230(w_015_230, w_000_1363, w_004_942);
  and2 I015_232(w_015_232, w_003_116, w_011_790);
  not1 I015_234(w_015_234, w_006_132);
  not1 I015_235(w_015_235, w_007_714);
  or2  I015_236(w_015_236, w_008_664, w_010_247);
  or2  I015_237(w_015_237, w_002_210, w_009_072);
  nand2 I015_238(w_015_238, w_012_324, w_000_1698);
  or2  I015_240(w_015_240, w_011_303, w_008_605);
  not1 I015_241(w_015_241, w_006_226);
  and2 I015_242(w_015_242, w_005_668, w_011_749);
  or2  I015_243(w_015_243, w_006_034, w_009_083);
  nand2 I015_244(w_015_244, w_010_039, w_005_612);
  nand2 I015_245(w_015_245, w_006_310, w_005_838);
  and2 I015_246(w_015_246, w_004_1235, w_003_095);
  nand2 I015_247(w_015_247, w_003_237, w_004_931);
  nand2 I015_248(w_015_248, w_007_1206, w_004_043);
  nand2 I015_249(w_015_249, w_008_677, w_004_1814);
  and2 I015_250(w_015_250, w_003_164, w_003_283);
  and2 I015_251(w_015_251, w_013_031, w_005_673);
  not1 I015_252(w_015_252, w_001_022);
  or2  I015_253(w_015_253, w_011_479, w_010_380);
  and2 I015_254(w_015_254, w_014_084, w_007_1567);
  not1 I015_255(w_015_255, w_011_194);
  not1 I015_256(w_015_256, w_011_639);
  and2 I015_257(w_015_257, w_005_199, w_008_591);
  not1 I015_258(w_015_258, w_008_184);
  and2 I015_259(w_015_259, w_007_1574, w_011_414);
  or2  I015_260(w_015_260, w_003_263, w_006_070);
  and2 I015_261(w_015_261, w_013_118, w_010_185);
  not1 I015_262(w_015_262, w_009_110);
  and2 I015_264(w_015_264, w_013_170, w_009_056);
  and2 I015_265(w_015_265, w_009_032, w_010_201);
  nand2 I015_266(w_015_266, w_013_287, w_001_283);
  nand2 I015_267(w_015_267, w_014_043, w_004_884);
  not1 I015_268(w_015_268, w_014_248);
  not1 I015_270(w_015_270, w_002_584);
  not1 I015_271(w_015_271, w_001_010);
  not1 I015_273(w_015_273, w_012_058);
  or2  I015_274(w_015_274, w_004_842, w_008_507);
  and2 I015_275(w_015_275, w_012_191, w_006_152);
  and2 I015_276(w_015_276, w_000_076, w_001_866);
  and2 I015_277(w_015_277, w_006_008, w_010_131);
  not1 I015_278(w_015_278, w_011_064);
  or2  I015_279(w_015_279, w_011_653, w_009_033);
  nand2 I015_280(w_015_280, w_006_308, w_011_757);
  not1 I015_281(w_015_281, w_004_130);
  not1 I015_282(w_015_282, w_008_673);
  nand2 I015_283(w_015_283, w_009_013, w_004_200);
  nand2 I015_285(w_015_285, w_011_685, w_004_1893);
  and2 I015_286(w_015_286, w_006_298, w_009_084);
  and2 I015_287(w_015_287, w_008_566, w_012_339);
  nand2 I015_288(w_015_288, w_000_1218, w_003_252);
  and2 I015_289(w_015_289, w_012_557, w_007_1246);
  nand2 I015_290(w_015_290, w_004_1799, w_010_197);
  and2 I015_291(w_015_291, w_003_015, w_009_044);
  nand2 I015_293(w_015_293, w_005_398, w_000_1888);
  or2  I016_000(w_016_000, w_010_272, w_010_401);
  and2 I016_001(w_016_001, w_012_043, w_008_203);
  not1 I016_002(w_016_002, w_011_354);
  and2 I016_003(w_016_003, w_000_1230, w_009_095);
  nand2 I016_004(w_016_004, w_005_580, w_008_419);
  nand2 I016_005(w_016_005, w_007_663, w_014_661);
  or2  I016_006(w_016_006, w_014_567, w_006_248);
  nand2 I016_007(w_016_007, w_000_1758, w_000_253);
  not1 I016_008(w_016_008, w_008_808);
  and2 I016_009(w_016_009, w_003_234, w_008_802);
  and2 I016_010(w_016_010, w_001_1666, w_015_128);
  not1 I016_011(w_016_011, w_007_058);
  or2  I016_012(w_016_012, w_014_721, w_008_818);
  not1 I016_013(w_016_013, w_006_059);
  and2 I016_014(w_016_014, w_015_260, w_009_077);
  not1 I016_015(w_016_015, w_006_007);
  not1 I016_016(w_016_016, w_014_432);
  or2  I016_017(w_016_017, w_008_599, w_004_032);
  not1 I016_018(w_016_018, w_007_295);
  and2 I016_019(w_016_019, w_013_338, w_011_739);
  and2 I016_020(w_016_020, w_012_455, w_007_1103);
  or2  I016_021(w_016_021, w_002_275, w_004_313);
  and2 I016_022(w_016_022, w_002_217, w_006_289);
  not1 I016_023(w_016_023, w_004_593);
  nand2 I016_024(w_016_024, w_012_410, w_004_476);
  and2 I016_025(w_016_025, w_011_395, w_004_1224);
  or2  I016_026(w_016_026, w_015_259, w_005_1228);
  not1 I016_027(w_016_027, w_013_331);
  and2 I016_028(w_016_028, w_015_146, w_008_696);
  nand2 I016_029(w_016_029, w_010_206, w_009_092);
  not1 I016_030(w_016_030, w_014_077);
  or2  I016_031(w_016_031, w_010_056, w_009_039);
  nand2 I016_032(w_016_032, w_004_1234, w_000_813);
  and2 I016_033(w_016_033, w_015_012, w_009_027);
  nand2 I016_034(w_016_034, w_006_158, w_015_090);
  or2  I016_035(w_016_035, w_007_102, w_012_002);
  not1 I016_036(w_016_036, w_005_670);
  and2 I016_037(w_016_037, w_003_299, w_002_120);
  nand2 I016_038(w_016_038, w_011_389, w_014_560);
  or2  I017_002(w_017_002, w_004_715, w_011_107);
  or2  I017_003(w_017_003, w_002_297, w_005_170);
  not1 I017_005(w_017_005, w_000_1922);
  and2 I017_006(w_017_006, w_016_002, w_011_136);
  and2 I017_007(w_017_007, w_013_074, w_005_1668);
  not1 I017_010(w_017_010, w_008_364);
  and2 I017_012(w_017_012, w_012_316, w_003_226);
  or2  I017_013(w_017_013, w_014_810, w_001_128);
  and2 I017_014(w_017_014, w_015_074, w_000_1923);
  and2 I017_016(w_017_016, w_002_020, w_012_395);
  and2 I017_017(w_017_017, w_014_740, w_007_1479);
  nand2 I017_018(w_017_018, w_010_273, w_004_191);
  not1 I017_019(w_017_019, w_007_977);
  and2 I017_020(w_017_020, w_016_015, w_010_405);
  or2  I017_022(w_017_022, w_007_1349, w_008_251);
  or2  I017_023(w_017_023, w_012_376, w_016_010);
  and2 I017_029(w_017_029, w_016_012, w_012_002);
  not1 I017_032(w_017_032, w_003_256);
  or2  I017_033(w_017_033, w_002_044, w_002_475);
  or2  I017_034(w_017_034, w_008_092, w_012_616);
  not1 I017_036(w_017_036, w_015_264);
  nand2 I017_038(w_017_038, w_010_365, w_008_352);
  or2  I017_040(w_017_040, w_002_390, w_016_030);
  not1 I017_044(w_017_044, w_011_533);
  or2  I017_045(w_017_045, w_010_043, w_003_097);
  not1 I017_046(w_017_046, w_012_656);
  nand2 I017_047(w_017_047, w_014_308, w_016_010);
  nand2 I017_052(w_017_052, w_008_779, w_016_014);
  and2 I017_057(w_017_057, w_014_397, w_009_068);
  or2  I017_059(w_017_059, w_007_1446, w_008_396);
  or2  I017_075(w_017_075, w_004_1703, w_016_002);
  not1 I017_077(w_017_077, w_011_542);
  and2 I017_084(w_017_084, w_000_1675, w_013_301);
  and2 I017_085(w_017_085, w_004_407, w_003_217);
  not1 I017_087(w_017_087, w_009_054);
  and2 I017_088(w_017_088, w_006_127, w_007_1366);
  nand2 I017_089(w_017_089, w_002_068, w_003_127);
  not1 I017_100(w_017_100, w_004_1716);
  not1 I017_102(w_017_102, w_008_112);
  nand2 I017_106(w_017_106, w_011_097, w_001_991);
  and2 I017_117(w_017_117, w_002_439, w_009_023);
  not1 I017_124(w_017_124, w_009_039);
  and2 I017_133(w_017_133, w_002_139, w_013_048);
  or2  I017_141(w_017_141, w_014_461, w_004_068);
  or2  I017_142(w_017_142, w_004_1111, w_013_135);
  or2  I017_143(w_017_143, w_011_318, w_009_073);
  and2 I017_150(w_017_150, w_000_1262, w_007_1269);
  not1 I017_155(w_017_155, w_008_195);
  and2 I017_158(w_017_158, w_006_166, w_006_007);
  and2 I017_159(w_017_159, w_001_1417, w_016_030);
  nand2 I017_162(w_017_162, w_013_076, w_013_303);
  and2 I017_171(w_017_171, w_011_101, w_014_578);
  and2 I017_174(w_017_174, w_004_990, w_009_024);
  nand2 I017_179(w_017_179, w_010_269, w_003_198);
  nand2 I017_183(w_017_183, w_001_1571, w_010_030);
  nand2 I017_194(w_017_194, w_014_179, w_007_014);
  or2  I017_197(w_017_197, w_013_094, w_009_047);
  nand2 I017_198(w_017_198, w_016_038, w_008_862);
  nand2 I017_203(w_017_203, w_001_1264, w_013_030);
  or2  I017_205(w_017_205, w_014_070, w_004_877);
  and2 I017_211(w_017_211, w_003_248, w_007_934);
  and2 I017_214(w_017_214, w_013_085, w_014_780);
  nand2 I017_218(w_017_218, w_008_475, w_009_086);
  nand2 I017_225(w_017_225, w_005_258, w_010_304);
  and2 I017_229(w_017_229, w_005_458, w_004_251);
  nand2 I017_234(w_017_234, w_008_093, w_002_342);
  not1 I017_236(w_017_236, w_001_542);
  not1 I017_240(w_017_240, w_006_258);
  and2 I017_244(w_017_244, w_001_949, w_015_006);
  nand2 I017_251(w_017_251, w_003_237, w_000_1925);
  not1 I017_253(w_017_253, w_015_040);
  not1 I017_254(w_017_254, w_016_019);
  and2 I017_264(w_017_264, w_003_122, w_001_1633);
  nand2 I017_269(w_017_269, w_016_015, w_014_219);
  nand2 I017_282(w_017_282, w_014_433, w_005_287);
  not1 I017_288(w_017_288, w_013_235);
  nand2 I017_299(w_017_299, w_013_295, w_007_171);
  nand2 I017_300(w_017_300, w_014_329, w_003_187);
  and2 I017_303(w_017_303, w_005_775, w_010_159);
  nand2 I017_305(w_017_305, w_016_021, w_000_417);
  nand2 I017_307(w_017_307, w_007_1321, w_008_506);
  and2 I017_315(w_017_315, w_006_276, w_008_450);
  or2  I017_317(w_017_317, w_000_279, w_012_348);
  not1 I017_322(w_017_322, w_001_1462);
  or2  I017_324(w_017_324, w_015_056, w_010_111);
  and2 I017_325(w_017_325, w_015_254, w_010_342);
  and2 I017_326(w_017_326, w_008_038, w_013_155);
  not1 I017_333(w_017_333, w_015_226);
  and2 I017_334(w_017_334, w_002_240, w_012_581);
  not1 I017_335(w_017_335, w_015_273);
  and2 I017_346(w_017_346, w_012_054, w_009_043);
  or2  I017_352(w_017_352, w_005_032, w_010_022);
  not1 I017_360(w_017_360, w_009_106);
  or2  I017_366(w_017_366, w_006_104, w_001_172);
  not1 I017_368(w_017_368, w_016_029);
  or2  I017_373(w_017_373, w_002_572, w_013_307);
  nand2 I017_381(w_017_381, w_013_154, w_014_027);
  not1 I017_384(w_017_384, w_004_384);
  and2 I017_385(w_017_385, w_016_020, w_013_123);
  and2 I017_386(w_017_386, w_002_176, w_007_1215);
  or2  I017_390(w_017_390, w_011_829, w_009_098);
  nand2 I017_393(w_017_393, w_007_1048, w_000_1555);
  nand2 I017_396(w_017_396, w_000_1692, w_013_151);
  not1 I017_397(w_017_397, w_005_1061);
  and2 I017_398(w_017_398, w_003_050, w_016_022);
  and2 I017_404(w_017_404, w_016_022, w_001_626);
  not1 I017_408(w_017_408, w_013_140);
  or2  I017_411(w_017_411, w_001_261, w_015_285);
  or2  I017_413(w_017_413, w_004_960, w_015_171);
  or2  I017_417(w_017_417, w_001_1225, w_016_000);
  not1 I017_427(w_017_427, w_008_850);
  not1 I017_428(w_017_428, w_005_556);
  or2  I017_429(w_017_429, w_000_1219, w_016_005);
  and2 I017_432(w_017_432, w_013_174, w_002_248);
  not1 I017_434(w_017_434, w_002_352);
  not1 I017_436(w_017_436, w_014_547);
  nand2 I017_442(w_017_442, w_000_332, w_003_224);
  or2  I017_446(w_017_446, w_003_289, w_007_152);
  or2  I017_450(w_017_450, w_006_306, w_007_1593);
  or2  I017_457(w_017_457, w_002_034, w_003_105);
  nand2 I017_459(w_017_459, w_012_049, w_002_522);
  or2  I017_468(w_017_468, w_009_073, w_007_1337);
  or2  I017_471(w_017_471, w_000_791, w_007_1566);
  or2  I017_472(w_017_472, w_006_305, w_010_015);
  nand2 I017_476(w_017_476, w_001_121, w_004_085);
  nand2 I017_478(w_017_478, w_000_1027, w_001_814);
  and2 I017_479(w_017_479, w_015_288, w_006_300);
  nand2 I017_482(w_017_482, w_010_131, w_014_249);
  nand2 I017_485(w_017_485, w_007_398, w_001_163);
  not1 I017_491(w_017_491, w_005_106);
  or2  I017_502(w_017_502, w_002_503, w_015_226);
  and2 I017_507(w_017_507, w_004_1595, w_006_263);
  or2  I017_508(w_017_508, w_010_091, w_015_255);
  nand2 I017_513(w_017_513, w_006_179, w_009_087);
  not1 I017_524(w_017_524, w_014_639);
  nand2 I017_525(w_017_525, w_012_530, w_012_524);
  or2  I017_528(w_017_528, w_007_720, w_009_012);
  or2  I017_534(w_017_534, w_013_021, w_012_628);
  not1 I017_539(w_017_539, w_002_125);
  nand2 I017_540(w_017_540, w_002_017, w_005_134);
  and2 I017_549(w_017_549, w_002_502, w_009_073);
  and2 I017_551(w_017_551, w_016_029, w_016_003);
  nand2 I017_556(w_017_556, w_009_013, w_000_1232);
  or2  I017_558(w_017_558, w_005_094, w_006_154);
  or2  I017_562(w_017_562, w_004_1589, w_012_472);
  and2 I017_589(w_017_589, w_005_268, w_016_030);
  and2 I017_595(w_017_595, w_004_991, w_000_1397);
  not1 I017_602(w_017_602, w_012_652);
  nand2 I017_605(w_017_605, w_011_704, w_011_574);
  and2 I017_615(w_017_615, w_014_169, w_005_320);
  nand2 I017_616(w_017_616, w_006_184, w_015_055);
  not1 I017_619(w_017_619, w_016_012);
  and2 I017_622(w_017_622, w_009_010, w_004_775);
  not1 I017_623(w_017_623, w_010_028);
  and2 I017_624(w_017_624, w_006_174, w_011_071);
  nand2 I017_631(w_017_631, w_016_013, w_011_219);
  not1 I017_633(w_017_633, w_015_235);
  and2 I017_644(w_017_644, w_009_081, w_004_280);
  not1 I017_647(w_017_647, w_012_059);
  nand2 I017_649(w_017_649, w_009_014, w_003_247);
  not1 I017_664(w_017_664, w_010_078);
  or2  I017_665(w_017_665, w_015_035, w_000_778);
  and2 I017_666(w_017_666, w_016_009, w_005_222);
  or2  I017_673(w_017_673, w_000_1199, w_004_1605);
  nand2 I017_675(w_017_675, w_008_210, w_014_274);
  or2  I017_677(w_017_677, w_002_017, w_006_102);
  or2  I017_678(w_017_678, w_009_083, w_015_186);
  and2 I017_681(w_017_681, w_012_154, w_000_1362);
  nand2 I017_684(w_017_684, w_011_163, w_008_198);
  or2  I017_685(w_017_685, w_005_1309, w_006_293);
  not1 I017_687(w_017_687, w_003_019);
  and2 I017_691(w_017_691, w_013_316, w_004_1080);
  nand2 I017_694(w_017_694, w_005_617, w_009_009);
  nand2 I017_697(w_017_697, w_012_020, w_014_626);
  and2 I017_702(w_017_702, w_003_112, w_013_163);
  not1 I017_703(w_017_703, w_003_209);
  not1 I017_704(w_017_704, w_000_435);
  or2  I017_707(w_017_707, w_006_216, w_011_339);
  not1 I017_713(w_017_713, w_010_238);
  not1 I017_722(w_017_722, w_001_1343);
  nand2 I017_723(w_017_723, w_009_085, w_007_147);
  or2  I017_730(w_017_730, w_005_809, w_000_1057);
  or2  I017_732(w_017_732, w_013_331, w_016_011);
  or2  I017_734(w_017_734, w_015_184, w_003_052);
  and2 I017_736(w_017_736, w_002_252, w_002_555);
  and2 I017_740(w_017_740, w_008_833, w_013_072);
  not1 I017_742(w_017_742, w_005_1293);
  nand2 I017_743(w_017_743, w_008_776, w_011_196);
  nand2 I017_744(w_017_744, w_005_1398, w_014_131);
  or2  I017_748(w_017_748, w_014_315, w_009_068);
  nand2 I017_753(w_017_753, w_007_105, w_007_168);
  nand2 I017_773(w_017_773, w_013_006, w_005_172);
  and2 I017_774(w_017_774, w_002_554, w_010_102);
  or2  I017_777(w_017_777, w_009_035, w_015_195);
  not1 I017_779(w_017_779, w_003_105);
  and2 I017_781(w_017_781, w_013_164, w_010_221);
  not1 I017_798(w_017_798, w_012_156);
  and2 I017_804(w_017_804, w_013_154, w_006_102);
  nand2 I017_805(w_017_805, w_013_320, w_015_285);
  nand2 I017_809(w_017_809, w_012_587, w_007_288);
  or2  I017_812(w_017_812, w_010_213, w_016_009);
  and2 I017_813(w_017_813, w_008_688, w_006_207);
  nand2 I017_821(w_017_821, w_001_216, w_008_166);
  nand2 I017_838(w_017_838, w_013_163, w_003_172);
  and2 I017_841(w_017_841, w_014_526, w_016_000);
  nand2 I017_845(w_017_845, w_004_633, w_004_1321);
  nand2 I017_846(w_017_846, w_003_105, w_014_509);
  and2 I017_847(w_017_847, w_010_384, w_011_126);
  or2  I017_851(w_017_851, w_015_113, w_013_148);
  nand2 I017_858(w_017_858, w_015_240, w_004_884);
  or2  I017_863(w_017_863, w_016_010, w_009_111);
  not1 I017_864(w_017_864, w_015_115);
  nand2 I017_867(w_017_867, w_016_003, w_000_1842);
  nand2 I017_871(w_017_871, w_016_006, w_014_650);
  or2  I017_873(w_017_873, w_012_399, w_011_474);
  or2  I017_875(w_017_875, w_014_024, w_012_222);
  and2 I017_885(w_017_885, w_014_330, w_003_075);
  or2  I017_891(w_017_891, w_009_047, w_007_1243);
  or2  I017_895(w_017_895, w_007_1460, w_008_772);
  not1 I017_896(w_017_896, w_015_286);
  and2 I017_899(w_017_899, w_008_829, w_000_1054);
  and2 I017_902(w_017_902, w_014_060, w_015_168);
  nand2 I017_903(w_017_903, w_005_911, w_012_394);
  nand2 I017_905(w_017_905, w_015_065, w_014_544);
  and2 I017_914(w_017_914, w_012_612, w_012_450);
  nand2 I017_917(w_017_917, w_001_1325, w_010_233);
  not1 I017_921(w_017_921, w_001_074);
  nand2 I017_929(w_017_929, w_014_099, w_001_1653);
  nand2 I017_932(w_017_932, w_012_599, w_016_013);
  and2 I017_933(w_017_933, w_006_127, w_014_304);
  and2 I017_935(w_017_935, w_003_281, w_009_044);
  not1 I017_944(w_017_944, w_008_074);
  or2  I017_947(w_017_947, w_001_597, w_009_053);
  and2 I017_950(w_017_950, w_013_090, w_003_120);
  or2  I017_953(w_017_953, w_013_192, w_007_1315);
  nand2 I017_956(w_017_956, w_014_525, w_013_177);
  nand2 I017_960(w_017_960, w_011_877, w_010_050);
  nand2 I017_967(w_017_967, w_002_494, w_010_112);
  nand2 I017_975(w_017_975, w_002_130, w_009_031);
  nand2 I017_977(w_017_977, w_015_042, w_012_141);
  and2 I017_982(w_017_982, w_004_790, w_009_068);
  and2 I017_984(w_017_984, w_009_017, w_006_209);
  and2 I017_985(w_017_985, w_011_548, w_008_222);
  nand2 I017_990(w_017_990, w_011_849, w_010_055);
  nand2 I017_998(w_017_998, w_011_735, w_009_017);
  nand2 I017_1000(w_017_1000, w_005_1274, w_007_357);
  not1 I017_1001(w_017_1001, w_002_126);
  or2  I017_1005(w_017_1005, w_001_1527, w_014_740);
  or2  I017_1006(w_017_1006, w_013_225, w_003_004);
  nand2 I017_1008(w_017_1008, w_011_560, w_008_082);
  and2 I017_1014(w_017_1014, w_003_233, w_011_483);
  and2 I017_1020(w_017_1020, w_008_002, w_007_101);
  not1 I017_1023(w_017_1023, w_013_323);
  not1 I017_1026(w_017_1026, w_010_397);
  and2 I017_1031(w_017_1031, w_007_313, w_013_081);
  and2 I017_1036(w_017_1036, w_006_191, w_015_177);
  and2 I017_1041(w_017_1041, w_011_035, w_012_262);
  or2  I017_1043(w_017_1043, w_012_132, w_003_219);
  and2 I017_1047(w_017_1047, w_009_107, w_004_496);
  and2 I017_1049(w_017_1049, w_013_125, w_014_532);
  nand2 I017_1051(w_017_1051, w_010_167, w_011_247);
  and2 I017_1058(w_017_1058, w_000_1074, w_005_1264);
  nand2 I017_1059(w_017_1059, w_007_603, w_002_160);
  and2 I017_1060(w_017_1060, w_010_176, w_008_759);
  and2 I017_1065(w_017_1065, w_015_225, w_015_116);
  not1 I017_1067(w_017_1067, w_011_088);
  nand2 I017_1070(w_017_1070, w_014_078, w_008_147);
  nand2 I017_1071(w_017_1071, w_013_083, w_001_737);
  nand2 I017_1074(w_017_1074, w_014_808, w_008_235);
  or2  I017_1077(w_017_1077, w_002_285, w_012_302);
  nand2 I017_1079(w_017_1079, w_005_127, w_001_1264);
  or2  I017_1092(w_017_1092, w_009_046, w_013_153);
  and2 I017_1098(w_017_1098, w_015_086, w_000_693);
  and2 I017_1101(w_017_1101, w_014_777, w_014_273);
  not1 I017_1103(w_017_1103, w_011_751);
  or2  I017_1104(w_017_1104, w_014_316, w_013_114);
  or2  I017_1109(w_017_1109, w_013_263, w_014_668);
  and2 I017_1111(w_017_1111, w_011_445, w_005_1101);
  not1 I017_1113(w_017_1113, w_009_055);
  not1 I017_1116(w_017_1116, w_012_246);
  and2 I017_1123(w_017_1123, w_005_640, w_010_237);
  nand2 I017_1126(w_017_1126, w_003_005, w_005_1181);
  or2  I017_1128(w_017_1128, w_011_316, w_006_045);
  not1 I017_1129(w_017_1129, w_008_195);
  and2 I017_1131(w_017_1131, w_009_005, w_001_906);
  or2  I017_1133(w_017_1133, w_010_246, w_006_249);
  and2 I017_1135(w_017_1135, w_004_1811, w_002_189);
  and2 I017_1139(w_017_1139, w_002_048, w_007_1444);
  not1 I017_1140(w_017_1140, w_005_037);
  not1 I017_1143(w_017_1143, w_001_1485);
  not1 I017_1145(w_017_1145, w_004_868);
  and2 I017_1153(w_017_1153, w_013_010, w_001_746);
  not1 I017_1163(w_017_1163, w_005_565);
  or2  I017_1165(w_017_1165, w_009_095, w_004_513);
  nand2 I017_1179(w_017_1179, w_007_1069, w_003_151);
  not1 I017_1182(w_017_1182, w_005_1645);
  or2  I017_1195(w_017_1195, w_002_461, w_009_035);
  or2  I017_1201(w_017_1201, w_000_1839, w_007_523);
  and2 I017_1206(w_017_1206, w_012_187, w_007_1454);
  or2  I017_1207(w_017_1207, w_014_191, w_001_1522);
  nand2 I017_1214(w_017_1214, w_013_230, w_004_001);
  nand2 I017_1216(w_017_1216, w_010_119, w_009_065);
  not1 I017_1218(w_017_1218, w_007_590);
  or2  I017_1220(w_017_1220, w_004_888, w_000_622);
  or2  I017_1223(w_017_1223, w_006_018, w_005_173);
  or2  I017_1224(w_017_1224, w_013_126, w_007_001);
  nand2 I017_1226(w_017_1226, w_004_1130, w_007_330);
  or2  I017_1227(w_017_1227, w_004_1463, w_014_663);
  and2 I017_1231(w_017_1231, w_005_1187, w_002_590);
  and2 I017_1232(w_017_1232, w_016_011, w_005_378);
  and2 I017_1237(w_017_1237, w_014_082, w_002_082);
  or2  I017_1238(w_017_1238, w_005_1266, w_009_030);
  or2  I017_1240(w_017_1240, w_014_349, w_006_060);
  not1 I017_1241(w_017_1241, w_001_668);
  not1 I017_1242(w_017_1242, w_003_182);
  nand2 I017_1244(w_017_1244, w_011_733, w_002_429);
  and2 I017_1246(w_017_1246, w_014_078, w_015_262);
  nand2 I017_1250(w_017_1250, w_000_1406, w_007_927);
  nand2 I017_1262(w_017_1262, w_013_263, w_013_050);
  not1 I017_1269(w_017_1269, w_015_220);
  and2 I017_1271(w_017_1271, w_007_349, w_011_320);
  and2 I017_1280(w_017_1280, w_000_540, w_000_327);
  or2  I017_1284(w_017_1284, w_013_066, w_008_560);
  or2  I017_1288(w_017_1288, w_004_229, w_003_158);
  not1 I017_1301(w_017_1301, w_008_799);
  nand2 I017_1308(w_017_1308, w_011_056, w_011_403);
  and2 I017_1310(w_017_1310, w_014_133, w_002_167);
  not1 I017_1312(w_017_1312, w_002_288);
  or2  I017_1322(w_017_1322, w_015_050, w_012_142);
  or2  I017_1325(w_017_1325, w_014_133, w_006_264);
  not1 I017_1327(w_017_1327, w_007_1307);
  or2  I017_1333(w_017_1333, w_016_016, w_012_330);
  or2  I017_1336(w_017_1336, w_010_259, w_002_027);
  not1 I017_1340(w_017_1340, w_010_174);
  nand2 I017_1348(w_017_1348, w_007_193, w_006_309);
  not1 I017_1351(w_017_1351, w_013_319);
  and2 I017_1354(w_017_1354, w_004_1248, w_005_196);
  not1 I017_1357(w_017_1357, w_006_218);
  not1 I017_1365(w_017_1365, w_010_080);
  not1 I017_1366(w_017_1366, w_013_216);
  or2  I017_1369(w_017_1369, w_007_734, w_002_067);
  or2  I017_1370(w_017_1370, w_012_085, w_008_741);
  not1 I017_1372(w_017_1372, w_014_123);
  and2 I017_1373(w_017_1373, w_001_010, w_000_1079);
  not1 I017_1374(w_017_1374, w_010_284);
  nand2 I017_1379(w_017_1379, w_016_025, w_016_028);
  or2  I017_1380(w_017_1380, w_000_1913, w_012_637);
  nand2 I017_1381(w_017_1381, w_005_605, w_004_1352);
  and2 I017_1383(w_017_1383, w_011_043, w_000_1472);
  or2  I017_1388(w_017_1388, w_008_703, w_001_042);
  nand2 I017_1391(w_017_1391, w_000_412, w_005_1297);
  or2  I017_1392(w_017_1392, w_008_237, w_010_175);
  not1 I017_1393(w_017_1393, w_009_072);
  and2 I017_1396(w_017_1396, w_009_071, w_004_1382);
  and2 I017_1397(w_017_1397, w_016_038, w_006_293);
  or2  I017_1400(w_017_1400, w_006_261, w_011_496);
  nand2 I017_1402(w_017_1402, w_006_286, w_010_025);
  nand2 I017_1407(w_017_1407, w_003_314, w_000_059);
  not1 I017_1410(w_017_1410, w_014_002);
  not1 I017_1416(w_017_1416, w_004_235);
  or2  I017_1419(w_017_1419, w_006_106, w_011_510);
  and2 I017_1421(w_017_1421, w_008_312, w_013_144);
  and2 I017_1422(w_017_1422, w_013_170, w_004_1216);
  or2  I017_1423(w_017_1423, w_016_008, w_009_080);
  not1 I017_1430(w_017_1430, w_009_007);
  not1 I017_1439(w_017_1439, w_013_180);
  nand2 I017_1443(w_017_1443, w_008_823, w_005_302);
  not1 I017_1445(w_017_1445, w_002_326);
  not1 I017_1448(w_017_1448, w_014_191);
  or2  I017_1449(w_017_1449, w_014_652, w_006_225);
  and2 I017_1453(w_017_1453, w_014_526, w_000_053);
  nand2 I017_1457(w_017_1457, w_008_353, w_012_243);
  and2 I017_1460(w_017_1460, w_013_247, w_006_285);
  and2 I017_1464(w_017_1464, w_014_459, w_014_359);
  nand2 I017_1469(w_017_1469, w_016_027, w_012_633);
  not1 I017_1480(w_017_1480, w_012_466);
  nand2 I017_1497(w_017_1497, w_007_026, w_000_1317);
  or2  I017_1504(w_017_1504, w_000_1435, w_013_125);
  nand2 I017_1505(w_017_1505, w_013_197, w_009_067);
  and2 I017_1517(w_017_1517, w_016_012, w_015_084);
  or2  I017_1530(w_017_1530, w_013_031, w_002_101);
  not1 I017_1531(w_017_1531, w_016_001);
  and2 I017_1533(w_017_1533, w_007_1597, w_002_184);
  nand2 I017_1534(w_017_1534, w_007_1397, w_006_170);
  nand2 I017_1541(w_017_1541, w_008_555, w_012_330);
  and2 I017_1550(w_017_1550, w_008_788, w_009_040);
  nand2 I017_1552(w_017_1552, w_016_011, w_007_144);
  nand2 I017_1556(w_017_1556, w_011_708, w_013_141);
  and2 I017_1557(w_017_1557, w_012_629, w_009_110);
  not1 I017_1563(w_017_1563, w_005_1187);
  or2  I017_1575(w_017_1575, w_007_036, w_012_147);
  not1 I017_1576(w_017_1576, w_005_713);
  and2 I017_1578(w_017_1578, w_012_511, w_008_151);
  and2 I017_1583(w_017_1583, w_007_925, w_015_078);
  and2 I017_1586(w_017_1586, w_003_188, w_009_091);
  and2 I017_1588(w_017_1588, w_015_225, w_015_000);
  not1 I017_1591(w_017_1591, w_012_000);
  and2 I017_1595(w_017_1595, w_012_349, w_006_282);
  not1 I017_1598(w_017_1598, w_013_122);
  or2  I017_1606(w_017_1606, w_016_026, w_002_511);
  and2 I017_1607(w_017_1607, w_013_013, w_000_1861);
  not1 I017_1612(w_017_1612, w_009_071);
  not1 I017_1622(w_017_1622, w_007_871);
  nand2 I017_1626(w_017_1626, w_002_063, w_013_331);
  and2 I017_1630(w_017_1630, w_011_553, w_002_276);
  not1 I017_1633(w_017_1633, w_006_073);
  not1 I017_1636(w_017_1636, w_000_715);
  and2 I017_1639(w_017_1639, w_004_035, w_011_229);
  or2  I017_1640(w_017_1640, w_009_043, w_006_128);
  nand2 I017_1645(w_017_1645, w_007_526, w_010_020);
  or2  I017_1646(w_017_1646, w_004_017, w_004_310);
  nand2 I017_1654(w_017_1654, w_016_026, w_006_059);
  nand2 I017_1655(w_017_1655, w_012_054, w_004_680);
  and2 I017_1656(w_017_1656, w_014_225, w_004_823);
  not1 I017_1658(w_017_1658, w_013_106);
  or2  I017_1665(w_017_1665, w_016_007, w_010_175);
  and2 I017_1666(w_017_1666, w_016_021, w_016_019);
  nand2 I017_1670(w_017_1670, w_006_063, w_013_004);
  or2  I017_1671(w_017_1671, w_008_013, w_015_074);
  or2  I017_1672(w_017_1672, w_000_1007, w_010_155);
  or2  I017_1679(w_017_1679, w_012_065, w_012_425);
  nand2 I017_1686(w_017_1686, w_003_280, w_012_332);
  or2  I017_1689(w_017_1689, w_004_1089, w_003_317);
  nand2 I017_1694(w_017_1694, w_002_008, w_007_194);
  not1 I017_1706(w_017_1706, w_004_1686);
  and2 I017_1707(w_017_1707, w_014_161, w_005_242);
  or2  I017_1710(w_017_1710, w_003_106, w_012_617);
  or2  I017_1715(w_017_1715, w_012_467, w_012_044);
  and2 I017_1718(w_017_1718, w_007_817, w_000_311);
  and2 I017_1727(w_017_1727, w_016_003, w_016_025);
  or2  I017_1729(w_017_1729, w_000_379, w_006_096);
  not1 I017_1732(w_017_1732, w_010_174);
  nand2 I017_1738(w_017_1738, w_009_111, w_014_015);
  nand2 I017_1743(w_017_1743, w_014_719, w_010_387);
  and2 I017_1750(w_017_1750, w_005_883, w_007_687);
  or2  I017_1753(w_017_1753, w_002_071, w_016_022);
  nand2 I017_1763(w_017_1763, w_015_074, w_009_100);
  nand2 I017_1768(w_017_1768, w_008_014, w_008_133);
  not1 I017_1778(w_017_1778, w_007_049);
  or2  I017_1792(w_017_1792, w_012_329, w_015_188);
  and2 I017_1797(w_017_1797, w_008_117, w_005_702);
  nand2 I017_1802(w_017_1802, w_010_065, w_004_1130);
  or2  I017_1809(w_017_1809, w_010_118, w_013_110);
  not1 I017_1814(w_017_1814, w_006_187);
  nand2 I017_1816(w_017_1816, w_005_971, w_002_373);
  and2 I017_1818(w_017_1818, w_007_1436, w_008_696);
  and2 I017_1822(w_017_1822, w_001_1211, w_001_311);
  nand2 I017_1823(w_017_1823, w_003_045, w_005_079);
  not1 I017_1828(w_017_1828, w_011_159);
  and2 I017_1831(w_017_1831, w_002_421, w_014_352);
  not1 I017_1839(w_017_1839, w_011_471);
  or2  I017_1852(w_017_1852, w_000_1370, w_002_546);
  and2 I017_1857(w_017_1857, w_006_154, w_004_1338);
  nand2 I017_1860(w_017_1860, w_004_746, w_009_066);
  or2  I017_1866(w_017_1866, w_000_511, w_007_618);
  and2 I017_1870(w_017_1870, w_005_817, w_001_035);
  not1 I017_1871(w_017_1871, w_011_210);
  not1 I017_1873(w_017_1873, w_001_873);
  and2 I017_1877(w_017_1877, w_014_008, w_014_469);
  nand2 I017_1878(w_017_1878, w_016_004, w_012_099);
  not1 I017_1881(w_017_1881, w_006_215);
  nand2 I017_1882(w_017_1882, w_006_025, w_000_632);
  not1 I017_1885(w_017_1885, w_001_150);
  or2  I017_1888(w_017_1888, w_013_215, w_006_302);
  or2  I017_1893(w_017_1893, w_000_406, w_013_206);
  or2  I017_1895(w_017_1895, w_012_342, w_010_365);
  nand2 I017_1900(w_017_1900, w_015_293, w_002_121);
  nand2 I017_1903(w_017_1903, w_016_038, w_016_027);
  nand2 I017_1910(w_017_1910, w_011_525, w_009_011);
  and2 I017_1911(w_017_1911, w_009_045, w_008_260);
  or2  I017_1913(w_017_1913, w_016_030, w_003_073);
  and2 I017_1923(w_017_1923, w_001_783, w_002_047);
  not1 I017_1924(w_017_1924, w_004_025);
  not1 I017_1935(w_017_1935, w_002_490);
  and2 I017_1937(w_017_1937, w_016_030, w_006_182);
  or2  I017_1945(w_017_1945, w_000_1099, w_005_213);
  and2 I017_1947(w_017_1947, w_005_562, w_009_049);
  and2 I018_003(w_018_003, w_001_032, w_000_046);
  or2  I018_004(w_018_004, w_013_073, w_011_002);
  nand2 I018_005(w_018_005, w_016_034, w_001_152);
  and2 I018_006(w_018_006, w_000_296, w_000_151);
  or2  I018_007(w_018_007, w_010_138, w_005_790);
  and2 I018_008(w_018_008, w_006_070, w_007_1600);
  not1 I018_009(w_018_009, w_011_085);
  not1 I018_010(w_018_010, w_009_024);
  nand2 I018_011(w_018_011, w_004_813, w_004_1078);
  or2  I018_012(w_018_012, w_001_283, w_006_125);
  nand2 I018_013(w_018_013, w_004_493, w_006_086);
  nand2 I018_014(w_018_014, w_016_007, w_002_382);
  not1 I018_015(w_018_015, w_007_1118);
  or2  I018_016(w_018_016, w_015_155, w_016_001);
  nand2 I018_017(w_018_017, w_007_266, w_003_293);
  and2 I018_018(w_018_018, w_005_363, w_017_386);
  not1 I018_019(w_018_019, w_005_584);
  and2 I018_021(w_018_021, w_014_574, w_001_162);
  and2 I018_022(w_018_022, w_008_106, w_011_257);
  not1 I018_024(w_018_024, w_016_000);
  not1 I018_025(w_018_025, w_004_558);
  nand2 I018_026(w_018_026, w_008_691, w_000_598);
  or2  I018_027(w_018_027, w_006_300, w_007_484);
  and2 I018_028(w_018_028, w_003_242, w_017_211);
  not1 I018_029(w_018_029, w_005_1534);
  nand2 I018_030(w_018_030, w_006_282, w_002_452);
  not1 I018_031(w_018_031, w_014_226);
  and2 I018_032(w_018_032, w_015_256, w_002_185);
  nand2 I018_033(w_018_033, w_011_107, w_003_193);
  not1 I018_035(w_018_035, w_017_373);
  or2  I018_036(w_018_036, w_010_338, w_011_669);
  nand2 I018_037(w_018_037, w_015_035, w_015_015);
  or2  I018_038(w_018_038, w_010_212, w_004_003);
  nand2 I018_039(w_018_039, w_004_323, w_010_089);
  not1 I018_040(w_018_040, w_014_767);
  nand2 I018_041(w_018_041, w_004_1100, w_017_556);
  and2 I018_043(w_018_043, w_009_041, w_017_046);
  and2 I018_044(w_018_044, w_014_777, w_007_268);
  nand2 I018_045(w_018_045, w_017_1743, w_005_1205);
  nand2 I018_046(w_018_046, w_009_088, w_001_1589);
  not1 I018_047(w_018_047, w_013_168);
  not1 I018_048(w_018_048, w_017_288);
  or2  I018_049(w_018_049, w_004_547, w_006_141);
  nand2 I018_050(w_018_050, w_013_186, w_016_003);
  not1 I018_052(w_018_052, w_012_371);
  and2 I018_054(w_018_054, w_016_025, w_017_1671);
  and2 I018_055(w_018_055, w_009_057, w_015_271);
  not1 I018_056(w_018_056, w_017_052);
  not1 I018_057(w_018_057, w_001_1671);
  not1 I018_059(w_018_059, w_011_404);
  and2 I018_061(w_018_061, w_017_1831, w_012_406);
  or2  I018_063(w_018_063, w_004_383, w_011_163);
  or2  I018_064(w_018_064, w_012_618, w_007_125);
  not1 I018_065(w_018_065, w_003_271);
  and2 I018_066(w_018_066, w_014_291, w_008_713);
  nand2 I018_067(w_018_067, w_003_200, w_013_270);
  nand2 I018_068(w_018_068, w_005_009, w_001_427);
  not1 I018_069(w_018_069, w_010_158);
  and2 I018_070(w_018_070, w_012_294, w_005_1033);
  and2 I018_071(w_018_071, w_017_1340, w_003_256);
  not1 I018_072(w_018_072, w_006_088);
  not1 I018_073(w_018_073, w_003_163);
  or2  I018_075(w_018_075, w_002_119, w_002_367);
  not1 I018_077(w_018_077, w_017_1895);
  and2 I018_078(w_018_078, w_010_210, w_002_162);
  nand2 I018_079(w_018_079, w_004_1319, w_007_048);
  nand2 I018_080(w_018_080, w_007_186, w_016_023);
  and2 I018_081(w_018_081, w_004_017, w_012_370);
  nand2 I018_082(w_018_082, w_012_589, w_000_1686);
  and2 I018_084(w_018_084, w_000_1481, w_008_059);
  nand2 I018_085(w_018_085, w_003_126, w_006_231);
  not1 I018_086(w_018_086, w_004_550);
  and2 I018_087(w_018_087, w_000_641, w_012_143);
  nand2 I018_088(w_018_088, w_004_1849, w_016_025);
  nand2 I018_089(w_018_089, w_014_519, w_000_1929);
  and2 I018_090(w_018_090, w_014_465, w_017_282);
  nand2 I018_091(w_018_091, w_005_1558, w_002_063);
  and2 I018_092(w_018_092, w_007_1584, w_000_551);
  and2 I018_094(w_018_094, w_010_054, w_015_087);
  not1 I018_097(w_018_097, w_010_007);
  or2  I018_098(w_018_098, w_013_205, w_004_1780);
  nand2 I018_100(w_018_100, w_017_1043, w_001_784);
  not1 I018_101(w_018_101, w_014_341);
  not1 I018_102(w_018_102, w_007_1562);
  or2  I018_103(w_018_103, w_014_119, w_016_016);
  and2 I018_104(w_018_104, w_006_313, w_010_035);
  nand2 I018_105(w_018_105, w_003_037, w_003_074);
  not1 I018_107(w_018_107, w_014_601);
  nand2 I018_108(w_018_108, w_005_257, w_009_069);
  not1 I018_109(w_018_109, w_014_447);
  or2  I018_110(w_018_110, w_015_242, w_001_814);
  nand2 I018_111(w_018_111, w_000_422, w_003_044);
  and2 I018_112(w_018_112, w_006_135, w_013_231);
  not1 I018_113(w_018_113, w_001_142);
  not1 I018_114(w_018_114, w_008_495);
  not1 I018_115(w_018_115, w_013_319);
  nand2 I018_117(w_018_117, w_014_504, w_002_189);
  nand2 I018_118(w_018_118, w_004_494, w_006_126);
  or2  I018_119(w_018_119, w_000_062, w_001_1437);
  and2 I018_120(w_018_120, w_003_107, w_007_769);
  or2  I018_121(w_018_121, w_015_129, w_001_601);
  and2 I018_122(w_018_122, w_008_564, w_017_006);
  or2  I018_124(w_018_124, w_017_102, w_007_1173);
  and2 I018_125(w_018_125, w_000_1435, w_009_007);
  nand2 I018_127(w_018_127, w_016_031, w_012_123);
  or2  I018_128(w_018_128, w_001_073, w_000_940);
  nand2 I018_129(w_018_129, w_005_1087, w_011_333);
  or2  I018_131(w_018_131, w_013_033, w_000_194);
  and2 I018_132(w_018_132, w_012_125, w_015_137);
  and2 I018_133(w_018_133, w_002_483, w_006_019);
  not1 I018_134(w_018_134, w_015_106);
  or2  I018_135(w_018_135, w_015_222, w_000_084);
  and2 I018_136(w_018_136, w_009_069, w_009_059);
  or2  I018_137(w_018_137, w_010_214, w_006_323);
  or2  I018_138(w_018_138, w_004_1558, w_014_370);
  nand2 I018_139(w_018_139, w_009_041, w_011_411);
  and2 I018_140(w_018_140, w_015_244, w_006_256);
  not1 I018_141(w_018_141, w_014_823);
  nand2 I018_142(w_018_142, w_012_240, w_015_174);
  or2  I018_143(w_018_143, w_004_657, w_013_124);
  not1 I018_144(w_018_144, w_017_847);
  nand2 I018_145(w_018_145, w_004_757, w_003_262);
  or2  I018_146(w_018_146, w_012_096, w_004_1110);
  and2 I018_147(w_018_147, w_000_588, w_013_180);
  nand2 I018_148(w_018_148, w_009_012, w_008_139);
  and2 I018_149(w_018_149, w_003_241, w_009_101);
  nand2 I018_150(w_018_150, w_002_139, w_011_018);
  and2 I018_151(w_018_151, w_000_1398, w_016_004);
  and2 I018_152(w_018_152, w_009_080, w_010_031);
  not1 I018_153(w_018_153, w_017_1639);
  and2 I018_155(w_018_155, w_008_742, w_008_577);
  and2 I018_156(w_018_156, w_017_1366, w_011_550);
  nand2 I018_157(w_018_157, w_002_326, w_003_136);
  not1 I018_158(w_018_158, w_001_1662);
  not1 I018_159(w_018_159, w_008_670);
  nand2 I018_160(w_018_160, w_002_517, w_012_035);
  and2 I018_161(w_018_161, w_006_215, w_010_070);
  nand2 I018_162(w_018_162, w_016_025, w_005_539);
  or2  I018_163(w_018_163, w_003_305, w_008_133);
  or2  I018_165(w_018_165, w_013_155, w_013_250);
  and2 I018_167(w_018_167, w_002_053, w_006_002);
  or2  I018_168(w_018_168, w_015_221, w_004_1153);
  not1 I018_170(w_018_170, w_009_060);
  nand2 I018_171(w_018_171, w_001_299, w_015_264);
  and2 I018_172(w_018_172, w_008_426, w_001_1066);
  nand2 I018_175(w_018_175, w_004_1296, w_003_165);
  nand2 I018_176(w_018_176, w_011_850, w_010_237);
  nand2 I018_178(w_018_178, w_009_037, w_005_243);
  not1 I018_180(w_018_180, w_006_273);
  and2 I018_181(w_018_181, w_013_060, w_009_041);
  or2  I018_182(w_018_182, w_011_538, w_004_990);
  or2  I018_183(w_018_183, w_012_175, w_016_024);
  nand2 I018_184(w_018_184, w_008_271, w_003_233);
  not1 I018_186(w_018_186, w_001_742);
  or2  I018_187(w_018_187, w_005_1088, w_017_1732);
  and2 I018_189(w_018_189, w_008_152, w_013_118);
  or2  I018_190(w_018_190, w_009_036, w_015_133);
  and2 I018_191(w_018_191, w_000_1122, w_001_226);
  not1 I018_192(w_018_192, w_015_142);
  or2  I018_193(w_018_193, w_014_118, w_000_1732);
  not1 I018_194(w_018_194, w_017_1816);
  nand2 I018_195(w_018_195, w_008_166, w_008_352);
  not1 I018_196(w_018_196, w_016_002);
  nand2 I018_197(w_018_197, w_001_1664, w_004_337);
  or2  I018_198(w_018_198, w_003_229, w_015_059);
  nand2 I018_200(w_018_200, w_002_302, w_005_546);
  not1 I018_201(w_018_201, w_005_078);
  not1 I018_202(w_018_202, w_004_172);
  not1 I018_203(w_018_203, w_014_168);
  nand2 I018_204(w_018_204, w_014_619, w_006_043);
  and2 I018_205(w_018_205, w_006_209, w_015_160);
  and2 I018_206(w_018_206, w_010_161, w_011_796);
  or2  I018_207(w_018_207, w_016_005, w_005_1257);
  not1 I018_209(w_018_209, w_003_101);
  not1 I018_210(w_018_210, w_003_216);
  and2 I018_211(w_018_211, w_009_059, w_016_035);
  or2  I018_212(w_018_212, w_005_1548, w_005_1584);
  or2  I018_213(w_018_213, w_009_008, w_007_577);
  or2  I018_214(w_018_214, w_009_046, w_001_1270);
  and2 I018_215(w_018_215, w_000_1789, w_010_222);
  nand2 I018_216(w_018_216, w_013_327, w_007_1194);
  and2 I018_218(w_018_218, w_001_400, w_002_039);
  and2 I018_219(w_018_219, w_000_1642, w_016_036);
  nand2 I018_220(w_018_220, w_017_012, w_006_202);
  nand2 I018_221(w_018_221, w_010_382, w_014_454);
  nand2 I018_222(w_018_222, w_015_193, w_004_980);
  or2  I018_223(w_018_223, w_014_617, w_014_208);
  not1 I018_224(w_018_224, w_014_708);
  not1 I018_225(w_018_225, w_015_171);
  not1 I018_226(w_018_226, w_015_165);
  not1 I018_227(w_018_227, w_002_259);
  nand2 I018_228(w_018_228, w_015_271, w_014_017);
  or2  I018_229(w_018_229, w_011_509, w_009_034);
  or2  I018_230(w_018_230, w_002_264, w_005_687);
  not1 I018_231(w_018_231, w_013_087);
  nand2 I018_232(w_018_232, w_003_048, w_001_082);
  or2  I018_233(w_018_233, w_006_038, w_012_155);
  or2  I018_234(w_018_234, w_012_340, w_008_170);
  nand2 I018_235(w_018_235, w_004_187, w_004_1221);
  and2 I018_236(w_018_236, w_011_371, w_015_157);
  and2 I018_237(w_018_237, w_003_204, w_012_266);
  nand2 I018_239(w_018_239, w_009_098, w_012_625);
  not1 I018_240(w_018_240, w_007_1033);
  not1 I018_241(w_018_241, w_015_027);
  not1 I018_242(w_018_242, w_000_1742);
  not1 I018_243(w_018_243, w_013_027);
  not1 I018_244(w_018_244, w_015_228);
  nand2 I018_245(w_018_245, w_005_120, w_016_036);
  or2  I018_246(w_018_246, w_008_157, w_009_064);
  not1 I018_248(w_018_248, w_012_341);
  nand2 I018_249(w_018_249, w_016_007, w_007_1596);
  nand2 I018_250(w_018_250, w_013_139, w_014_372);
  or2  I018_251(w_018_251, w_009_021, w_016_029);
  and2 I018_252(w_018_252, w_014_690, w_004_220);
  or2  I018_253(w_018_253, w_011_872, w_002_363);
  or2  I018_254(w_018_254, w_006_270, w_013_090);
  nand2 I018_255(w_018_255, w_013_337, w_014_286);
  or2  I018_256(w_018_256, w_013_307, w_004_1478);
  and2 I018_257(w_018_257, w_011_543, w_003_302);
  and2 I018_258(w_018_258, w_013_230, w_000_1327);
  nand2 I018_259(w_018_259, w_017_446, w_005_124);
  not1 I018_260(w_018_260, w_011_870);
  and2 I018_261(w_018_261, w_004_524, w_005_1079);
  or2  I018_262(w_018_262, w_000_197, w_015_191);
  or2  I018_263(w_018_263, w_017_845, w_005_1117);
  or2  I018_264(w_018_264, w_008_699, w_011_783);
  or2  I018_265(w_018_265, w_009_003, w_006_002);
  or2  I018_266(w_018_266, w_012_465, w_009_033);
  nand2 I018_267(w_018_267, w_001_1637, w_000_763);
  or2  I018_268(w_018_268, w_015_257, w_006_128);
  not1 I018_269(w_018_269, w_001_476);
  and2 I018_271(w_018_271, w_012_490, w_001_1101);
  or2  I018_272(w_018_272, w_008_238, w_002_180);
  and2 I018_273(w_018_273, w_010_035, w_014_117);
  and2 I018_274(w_018_274, w_012_376, w_017_1945);
  nand2 I018_275(w_018_275, w_006_074, w_006_179);
  not1 I018_276(w_018_276, w_008_211);
  and2 I018_278(w_018_278, w_010_132, w_001_522);
  or2  I018_279(w_018_279, w_002_460, w_015_142);
  nand2 I018_280(w_018_280, w_011_795, w_010_307);
  and2 I018_281(w_018_281, w_007_1095, w_007_601);
  or2  I018_282(w_018_282, w_013_165, w_007_327);
  not1 I019_000(w_019_000, w_011_159);
  or2  I019_001(w_019_001, w_017_236, w_007_325);
  or2  I019_002(w_019_002, w_012_378, w_016_014);
  not1 I019_005(w_019_005, w_009_095);
  nand2 I019_010(w_019_010, w_008_646, w_002_486);
  or2  I019_011(w_019_011, w_001_700, w_018_252);
  not1 I019_014(w_019_014, w_008_707);
  and2 I019_019(w_019_019, w_003_139, w_011_383);
  and2 I019_020(w_019_020, w_014_020, w_015_164);
  not1 I019_021(w_019_021, w_004_325);
  not1 I019_023(w_019_023, w_013_295);
  nand2 I019_024(w_019_024, w_003_135, w_017_1388);
  and2 I019_025(w_019_025, w_003_122, w_018_151);
  and2 I019_027(w_019_027, w_008_646, w_015_181);
  and2 I019_028(w_019_028, w_017_1430, w_012_016);
  or2  I019_030(w_019_030, w_015_122, w_012_484);
  or2  I019_031(w_019_031, w_012_279, w_017_404);
  nand2 I019_032(w_019_032, w_017_846, w_017_411);
  nand2 I019_040(w_019_040, w_014_029, w_006_009);
  nand2 I019_055(w_019_055, w_018_078, w_005_328);
  and2 I019_058(w_019_058, w_002_064, w_018_280);
  not1 I019_062(w_019_062, w_005_816);
  nand2 I019_071(w_019_071, w_010_246, w_004_1123);
  nand2 I019_074(w_019_074, w_005_1276, w_012_327);
  and2 I019_077(w_019_077, w_012_008, w_007_1449);
  or2  I019_080(w_019_080, w_006_055, w_017_1658);
  nand2 I019_081(w_019_081, w_011_501, w_000_694);
  and2 I019_082(w_019_082, w_016_017, w_000_389);
  not1 I019_083(w_019_083, w_010_273);
  not1 I019_085(w_019_085, w_013_328);
  not1 I019_089(w_019_089, w_000_964);
  or2  I019_090(w_019_090, w_006_189, w_003_280);
  not1 I019_091(w_019_091, w_002_382);
  or2  I019_092(w_019_092, w_012_636, w_002_259);
  not1 I019_097(w_019_097, w_007_058);
  or2  I019_099(w_019_099, w_016_015, w_017_1893);
  not1 I019_101(w_019_101, w_003_031);
  not1 I019_105(w_019_105, w_010_306);
  nand2 I019_106(w_019_106, w_006_063, w_012_201);
  not1 I019_110(w_019_110, w_013_311);
  not1 I019_113(w_019_113, w_012_643);
  nand2 I019_115(w_019_115, w_018_006, w_004_086);
  nand2 I019_122(w_019_122, w_001_955, w_017_1533);
  not1 I019_123(w_019_123, w_018_114);
  and2 I019_124(w_019_124, w_012_141, w_006_191);
  not1 I019_127(w_019_127, w_000_036);
  not1 I019_128(w_019_128, w_014_013);
  and2 I019_130(w_019_130, w_008_386, w_001_1001);
  not1 I019_132(w_019_132, w_010_048);
  not1 I019_133(w_019_133, w_012_541);
  nand2 I019_135(w_019_135, w_012_598, w_002_306);
  not1 I019_139(w_019_139, w_008_290);
  not1 I019_141(w_019_141, w_005_800);
  or2  I019_142(w_019_142, w_004_1394, w_000_766);
  and2 I019_144(w_019_144, w_017_434, w_014_225);
  not1 I019_145(w_019_145, w_016_008);
  or2  I019_150(w_019_150, w_012_119, w_015_046);
  nand2 I019_151(w_019_151, w_010_008, w_005_1309);
  not1 I019_152(w_019_152, w_000_1902);
  not1 I019_153(w_019_153, w_005_769);
  and2 I019_161(w_019_161, w_010_366, w_011_204);
  and2 I019_164(w_019_164, w_016_004, w_018_054);
  nand2 I019_165(w_019_165, w_017_697, w_006_001);
  nand2 I019_167(w_019_167, w_016_009, w_002_292);
  and2 I019_176(w_019_176, w_012_293, w_004_1732);
  nand2 I019_183(w_019_183, w_010_005, w_000_111);
  or2  I019_188(w_019_188, w_018_111, w_008_484);
  nand2 I019_189(w_019_189, w_015_203, w_018_215);
  nand2 I019_190(w_019_190, w_018_043, w_015_243);
  and2 I019_191(w_019_191, w_005_281, w_008_821);
  or2  I019_192(w_019_192, w_000_1551, w_017_1591);
  and2 I019_201(w_019_201, w_018_077, w_003_114);
  or2  I019_202(w_019_202, w_011_258, w_001_266);
  or2  I019_204(w_019_204, w_013_227, w_000_1390);
  and2 I019_205(w_019_205, w_017_1877, w_015_134);
  nand2 I019_206(w_019_206, w_006_242, w_002_163);
  or2  I019_209(w_019_209, w_003_039, w_006_190);
  nand2 I019_212(w_019_212, w_005_160, w_004_1063);
  nand2 I019_213(w_019_213, w_006_194, w_010_386);
  nand2 I019_216(w_019_216, w_012_506, w_016_023);
  not1 I019_219(w_019_219, w_015_067);
  or2  I019_220(w_019_220, w_018_278, w_003_257);
  nand2 I019_222(w_019_222, w_017_100, w_011_267);
  not1 I019_225(w_019_225, w_001_1100);
  not1 I019_229(w_019_229, w_002_523);
  or2  I019_230(w_019_230, w_000_1264, w_018_253);
  nand2 I019_232(w_019_232, w_008_395, w_001_451);
  or2  I019_234(w_019_234, w_009_038, w_014_322);
  not1 I019_237(w_019_237, w_008_085);
  or2  I019_239(w_019_239, w_003_001, w_010_196);
  not1 I019_240(w_019_240, w_007_1390);
  not1 I019_244(w_019_244, w_018_124);
  not1 I019_246(w_019_246, w_008_766);
  nand2 I019_250(w_019_250, w_014_808, w_004_872);
  or2  I019_252(w_019_252, w_008_680, w_014_685);
  not1 I019_253(w_019_253, w_004_635);
  nand2 I019_257(w_019_257, w_010_231, w_004_202);
  nand2 I019_259(w_019_259, w_016_038, w_010_082);
  and2 I019_262(w_019_262, w_006_153, w_010_235);
  or2  I019_269(w_019_269, w_017_1480, w_014_582);
  or2  I019_273(w_019_273, w_018_112, w_005_1078);
  not1 I019_277(w_019_277, w_015_144);
  and2 I019_278(w_019_278, w_001_138, w_017_1123);
  or2  I019_279(w_019_279, w_010_054, w_014_663);
  and2 I019_284(w_019_284, w_009_093, w_014_406);
  nand2 I019_287(w_019_287, w_010_402, w_002_086);
  or2  I019_288(w_019_288, w_000_110, w_015_164);
  or2  I019_289(w_019_289, w_012_637, w_013_102);
  and2 I019_290(w_019_290, w_009_076, w_015_262);
  and2 I019_292(w_019_292, w_003_160, w_017_1246);
  or2  I019_294(w_019_294, w_008_308, w_000_1625);
  and2 I019_296(w_019_296, w_002_028, w_007_604);
  not1 I019_297(w_019_297, w_016_006);
  and2 I019_298(w_019_298, w_018_036, w_014_234);
  nand2 I019_302(w_019_302, w_016_035, w_013_294);
  or2  I019_303(w_019_303, w_001_610, w_013_289);
  nand2 I019_304(w_019_304, w_004_758, w_000_296);
  and2 I019_305(w_019_305, w_009_102, w_002_033);
  or2  I019_310(w_019_310, w_013_315, w_010_168);
  not1 I019_317(w_019_317, w_016_005);
  or2  I019_326(w_019_326, w_001_298, w_006_193);
  and2 I019_328(w_019_328, w_014_107, w_010_158);
  not1 I019_329(w_019_329, w_004_1186);
  not1 I019_331(w_019_331, w_014_221);
  not1 I019_338(w_019_338, w_001_302);
  not1 I019_339(w_019_339, w_005_055);
  or2  I019_340(w_019_340, w_014_014, w_005_1082);
  and2 I019_342(w_019_342, w_016_025, w_013_279);
  and2 I019_343(w_019_343, w_005_1581, w_007_1340);
  nand2 I019_344(w_019_344, w_015_289, w_002_069);
  or2  I019_347(w_019_347, w_005_1480, w_002_034);
  nand2 I019_350(w_019_350, w_015_270, w_017_1280);
  nand2 I019_353(w_019_353, w_001_852, w_010_166);
  and2 I019_358(w_019_358, w_006_274, w_002_274);
  nand2 I019_359(w_019_359, w_013_292, w_012_168);
  nand2 I019_360(w_019_360, w_002_335, w_014_801);
  nand2 I019_361(w_019_361, w_017_1237, w_007_1494);
  or2  I019_365(w_019_365, w_003_308, w_001_1305);
  not1 I019_368(w_019_368, w_006_236);
  not1 I019_369(w_019_369, w_013_307);
  not1 I019_374(w_019_374, w_016_031);
  nand2 I019_377(w_019_377, w_008_165, w_014_049);
  nand2 I019_383(w_019_383, w_007_796, w_014_041);
  not1 I019_385(w_019_385, w_003_293);
  or2  I019_386(w_019_386, w_002_583, w_004_1663);
  and2 I019_387(w_019_387, w_006_186, w_013_087);
  or2  I019_389(w_019_389, w_010_266, w_009_083);
  not1 I019_391(w_019_391, w_005_341);
  not1 I019_395(w_019_395, w_015_290);
  nand2 I019_397(w_019_397, w_009_051, w_007_1123);
  nand2 I019_401(w_019_401, w_005_1526, w_001_864);
  or2  I019_402(w_019_402, w_016_023, w_002_493);
  or2  I019_404(w_019_404, w_006_132, w_007_119);
  not1 I019_405(w_019_405, w_003_017);
  and2 I019_406(w_019_406, w_005_911, w_010_074);
  nand2 I019_407(w_019_407, w_007_1536, w_004_1843);
  not1 I019_409(w_019_409, w_001_246);
  not1 I019_411(w_019_411, w_004_046);
  not1 I019_415(w_019_415, w_005_179);
  not1 I019_416(w_019_416, w_002_420);
  nand2 I019_417(w_019_417, w_010_088, w_017_742);
  not1 I019_419(w_019_419, w_013_016);
  not1 I019_420(w_019_420, w_017_1001);
  or2  I019_423(w_019_423, w_004_1001, w_015_222);
  nand2 I019_428(w_019_428, w_002_222, w_008_472);
  and2 I019_430(w_019_430, w_001_1005, w_002_119);
  and2 I019_436(w_019_436, w_016_036, w_002_083);
  nand2 I019_437(w_019_437, w_001_294, w_000_277);
  or2  I019_438(w_019_438, w_005_898, w_010_239);
  not1 I019_439(w_019_439, w_006_033);
  or2  I019_441(w_019_441, w_001_1440, w_002_399);
  or2  I019_445(w_019_445, w_017_315, w_011_802);
  nand2 I019_449(w_019_449, w_000_257, w_009_019);
  not1 I019_450(w_019_450, w_011_009);
  nand2 I019_451(w_019_451, w_013_176, w_009_104);
  or2  I019_459(w_019_459, w_000_1598, w_009_044);
  not1 I019_463(w_019_463, w_003_018);
  not1 I019_465(w_019_465, w_008_861);
  or2  I019_467(w_019_467, w_000_741, w_000_1121);
  or2  I019_470(w_019_470, w_003_086, w_011_633);
  nand2 I019_474(w_019_474, w_009_083, w_017_1336);
  not1 I019_476(w_019_476, w_009_007);
  or2  I019_478(w_019_478, w_016_036, w_013_064);
  not1 I019_480(w_019_480, w_005_1010);
  or2  I019_481(w_019_481, w_011_109, w_011_297);
  or2  I019_482(w_019_482, w_016_012, w_005_578);
  nand2 I019_485(w_019_485, w_009_026, w_015_249);
  nand2 I019_486(w_019_486, w_010_373, w_016_035);
  and2 I019_487(w_019_487, w_002_167, w_002_046);
  not1 I019_488(w_019_488, w_011_695);
  or2  I019_491(w_019_491, w_004_788, w_017_685);
  not1 I019_494(w_019_494, w_013_338);
  and2 I019_499(w_019_499, w_000_1239, w_017_1689);
  nand2 I019_500(w_019_500, w_012_574, w_002_205);
  and2 I019_504(w_019_504, w_018_117, w_009_030);
  not1 I019_505(w_019_505, w_004_701);
  and2 I019_507(w_019_507, w_003_207, w_014_279);
  and2 I019_512(w_019_512, w_017_1923, w_010_325);
  or2  I019_514(w_019_514, w_015_241, w_016_006);
  nand2 I019_516(w_019_516, w_001_824, w_018_129);
  or2  I019_519(w_019_519, w_011_163, w_004_1664);
  not1 I019_521(w_019_521, w_002_551);
  or2  I019_524(w_019_524, w_007_1148, w_017_384);
  not1 I019_525(w_019_525, w_011_624);
  nand2 I019_526(w_019_526, w_004_555, w_018_193);
  or2  I019_527(w_019_527, w_004_104, w_014_276);
  or2  I019_530(w_019_530, w_006_023, w_001_1627);
  nand2 I019_537(w_019_537, w_001_1241, w_017_1023);
  nand2 I019_538(w_019_538, w_007_224, w_009_023);
  not1 I019_543(w_019_543, w_007_441);
  nand2 I019_544(w_019_544, w_005_1464, w_014_097);
  and2 I019_545(w_019_545, w_004_952, w_012_233);
  not1 I019_547(w_019_547, w_003_116);
  or2  I019_551(w_019_551, w_018_226, w_004_383);
  or2  I019_552(w_019_552, w_016_038, w_018_242);
  or2  I019_553(w_019_553, w_015_093, w_008_314);
  not1 I019_556(w_019_556, w_015_227);
  nand2 I019_558(w_019_558, w_011_848, w_006_154);
  or2  I019_559(w_019_559, w_002_027, w_010_191);
  nand2 I019_560(w_019_560, w_016_004, w_016_019);
  not1 I019_563(w_019_563, w_002_523);
  or2  I019_568(w_019_568, w_003_282, w_016_036);
  not1 I019_569(w_019_569, w_006_063);
  and2 I019_571(w_019_571, w_014_664, w_009_005);
  nand2 I019_573(w_019_573, w_007_555, w_008_618);
  or2  I019_575(w_019_575, w_017_1818, w_001_1580);
  nand2 I019_577(w_019_577, w_009_100, w_000_869);
  and2 I019_580(w_019_580, w_010_165, w_013_090);
  nand2 I019_583(w_019_583, w_011_256, w_017_1612);
  not1 I019_585(w_019_585, w_010_405);
  nand2 I019_586(w_019_586, w_008_817, w_002_042);
  not1 I019_590(w_019_590, w_002_291);
  and2 I019_593(w_019_593, w_008_071, w_007_1022);
  not1 I019_595(w_019_595, w_010_095);
  or2  I019_596(w_019_596, w_007_1190, w_014_487);
  and2 I019_597(w_019_597, w_017_953, w_008_426);
  nand2 I019_598(w_019_598, w_005_497, w_001_322);
  not1 I019_599(w_019_599, w_017_1576);
  and2 I019_601(w_019_601, w_005_165, w_000_523);
  or2  I019_604(w_019_604, w_005_204, w_004_472);
  not1 I019_608(w_019_608, w_008_095);
  or2  I019_610(w_019_610, w_018_137, w_014_115);
  not1 I019_613(w_019_613, w_015_170);
  and2 I019_614(w_019_614, w_014_023, w_011_466);
  not1 I019_615(w_019_615, w_003_081);
  or2  I019_617(w_019_617, w_011_350, w_003_051);
  nand2 I019_618(w_019_618, w_010_006, w_008_638);
  or2  I019_619(w_019_619, w_001_1661, w_004_1604);
  or2  I019_625(w_019_625, w_000_556, w_018_210);
  not1 I019_627(w_019_627, w_007_104);
  and2 I019_629(w_019_629, w_013_095, w_004_1868);
  nand2 I019_631(w_019_631, w_011_429, w_003_233);
  not1 I019_632(w_019_632, w_008_298);
  nand2 I019_633(w_019_633, w_006_302, w_013_001);
  and2 I019_637(w_019_637, w_016_030, w_001_250);
  not1 I019_643(w_019_643, w_007_060);
  and2 I019_647(w_019_647, w_007_664, w_012_194);
  not1 I019_648(w_019_648, w_007_017);
  and2 I019_655(w_019_655, w_018_071, w_002_179);
  nand2 I019_656(w_019_656, w_009_056, w_000_975);
  not1 I019_657(w_019_657, w_011_580);
  not1 I019_659(w_019_659, w_005_398);
  not1 I019_665(w_019_665, w_006_256);
  not1 I019_666(w_019_666, w_010_260);
  nand2 I019_668(w_019_668, w_013_029, w_011_482);
  not1 I019_671(w_019_671, w_014_232);
  or2  I019_673(w_019_673, w_013_253, w_013_205);
  nand2 I019_675(w_019_675, w_004_172, w_008_423);
  not1 I019_682(w_019_682, w_004_1086);
  or2  I019_689(w_019_689, w_013_315, w_002_247);
  nand2 I019_691(w_019_691, w_012_488, w_007_367);
  not1 I019_692(w_019_692, w_008_081);
  nand2 I019_695(w_019_695, w_001_295, w_004_850);
  or2  I019_699(w_019_699, w_010_272, w_003_058);
  nand2 I019_700(w_019_700, w_000_1766, w_018_158);
  and2 I019_701(w_019_701, w_013_190, w_004_011);
  nand2 I019_702(w_019_702, w_008_348, w_005_014);
  or2  I019_705(w_019_705, w_002_519, w_003_066);
  and2 I019_706(w_019_706, w_006_316, w_004_540);
  not1 I019_707(w_019_707, w_003_182);
  or2  I019_709(w_019_709, w_005_1251, w_012_157);
  not1 I019_710(w_019_710, w_018_066);
  nand2 I019_717(w_019_717, w_016_030, w_012_189);
  nand2 I019_718(w_019_718, w_010_105, w_000_1568);
  not1 I019_721(w_019_721, w_009_034);
  not1 I019_722(w_019_722, w_000_940);
  or2  I019_723(w_019_723, w_016_018, w_014_745);
  nand2 I019_724(w_019_724, w_013_028, w_005_1393);
  not1 I019_726(w_019_726, w_017_1729);
  or2  I019_729(w_019_729, w_008_799, w_014_734);
  nand2 I019_732(w_019_732, w_015_223, w_016_025);
  or2  I019_745(w_019_745, w_008_108, w_012_569);
  and2 I019_748(w_019_748, w_018_157, w_012_515);
  or2  I019_753(w_019_753, w_016_019, w_001_430);
  or2  I019_754(w_019_754, w_008_661, w_008_841);
  nand2 I019_755(w_019_755, w_001_1044, w_000_1612);
  nand2 I019_756(w_019_756, w_010_274, w_013_069);
  not1 I019_757(w_019_757, w_004_1420);
  nand2 I019_761(w_019_761, w_001_769, w_014_205);
  or2  I019_763(w_019_763, w_009_022, w_002_122);
  nand2 I019_766(w_019_766, w_012_310, w_002_360);
  nand2 I019_770(w_019_770, w_012_465, w_008_694);
  or2  I019_771(w_019_771, w_008_317, w_011_496);
  nand2 I019_772(w_019_772, w_012_597, w_006_101);
  or2  I019_773(w_019_773, w_015_117, w_009_047);
  not1 I019_775(w_019_775, w_006_294);
  and2 I019_776(w_019_776, w_012_509, w_001_805);
  nand2 I019_778(w_019_778, w_015_151, w_009_066);
  nand2 I019_782(w_019_782, w_006_166, w_016_030);
  nand2 I019_783(w_019_783, w_009_110, w_012_276);
  and2 I019_784(w_019_784, w_000_1147, w_012_388);
  or2  I019_786(w_019_786, w_006_134, w_012_199);
  and2 I019_790(w_019_790, w_005_1495, w_012_482);
  nand2 I019_791(w_019_791, w_014_060, w_002_176);
  and2 I019_797(w_019_797, w_009_013, w_016_013);
  not1 I019_800(w_019_800, w_009_005);
  or2  I019_808(w_019_808, w_000_021, w_008_748);
  and2 I019_812(w_019_812, w_010_262, w_003_304);
  nand2 I019_814(w_019_814, w_002_335, w_000_163);
  and2 I019_815(w_019_815, w_006_056, w_012_346);
  and2 I019_817(w_019_817, w_012_102, w_009_052);
  not1 I019_819(w_019_819, w_005_1480);
  or2  I019_825(w_019_825, w_005_1540, w_002_075);
  not1 I019_831(w_019_831, w_008_359);
  and2 I019_834(w_019_834, w_009_079, w_007_118);
  not1 I019_836(w_019_836, w_001_666);
  or2  I019_842(w_019_842, w_017_036, w_013_030);
  not1 I019_843(w_019_843, w_015_283);
  nand2 I019_844(w_019_844, w_010_214, w_008_064);
  or2  I019_845(w_019_845, w_001_346, w_007_863);
  not1 I019_849(w_019_849, w_013_235);
  not1 I019_858(w_019_858, w_011_551);
  or2  I019_859(w_019_859, w_011_384, w_012_087);
  not1 I019_860(w_019_860, w_016_005);
  or2  I019_864(w_019_864, w_009_109, w_016_031);
  nand2 I019_865(w_019_865, w_005_376, w_009_003);
  and2 I019_866(w_019_866, w_002_081, w_006_194);
  not1 I019_868(w_019_868, w_005_747);
  not1 I019_876(w_019_876, w_001_020);
  nand2 I019_877(w_019_877, w_003_118, w_015_015);
  or2  I019_879(w_019_879, w_000_1333, w_015_188);
  or2  I019_881(w_019_881, w_011_039, w_015_142);
  nand2 I019_882(w_019_882, w_004_1727, w_015_050);
  or2  I019_888(w_019_888, w_000_1857, w_016_007);
  or2  I019_890(w_019_890, w_015_207, w_002_526);
  or2  I019_893(w_019_893, w_000_1585, w_018_071);
  nand2 I019_894(w_019_894, w_015_047, w_000_1018);
  nand2 I019_897(w_019_897, w_003_031, w_004_1112);
  not1 I019_898(w_019_898, w_017_1445);
  or2  I019_900(w_019_900, w_002_193, w_001_1674);
  nand2 I019_905(w_019_905, w_001_1453, w_011_108);
  and2 I019_908(w_019_908, w_014_495, w_010_049);
  not1 I019_909(w_019_909, w_004_952);
  and2 I019_917(w_019_917, w_011_163, w_002_406);
  nand2 I019_918(w_019_918, w_018_205, w_010_323);
  not1 I019_920(w_019_920, w_014_110);
  not1 I019_926(w_019_926, w_002_177);
  nand2 I019_951(w_019_951, w_002_340, w_008_831);
  not1 I019_953(w_019_953, w_014_040);
  and2 I019_958(w_019_958, w_007_1187, w_011_122);
  and2 I019_960(w_019_960, w_011_020, w_016_006);
  nand2 I019_962(w_019_962, w_015_230, w_001_279);
  or2  I019_965(w_019_965, w_000_1590, w_006_243);
  and2 I019_968(w_019_968, w_009_029, w_008_646);
  or2  I019_975(w_019_975, w_007_1600, w_011_575);
  nand2 I019_978(w_019_978, w_007_1350, w_010_391);
  or2  I019_980(w_019_980, w_015_084, w_002_028);
  nand2 I019_994(w_019_994, w_000_1931, w_005_286);
  and2 I019_1007(w_019_1007, w_006_121, w_006_301);
  and2 I019_1008(w_019_1008, w_010_242, w_008_172);
  or2  I019_1017(w_019_1017, w_012_646, w_012_221);
  or2  I019_1019(w_019_1019, w_001_1307, w_004_1092);
  and2 I019_1021(w_019_1021, w_005_1090, w_009_080);
  and2 I019_1022(w_019_1022, w_004_782, w_005_136);
  and2 I019_1026(w_019_1026, w_014_181, w_003_138);
  or2  I019_1029(w_019_1029, w_009_021, w_016_036);
  or2  I019_1031(w_019_1031, w_016_012, w_006_058);
  or2  I019_1036(w_019_1036, w_016_002, w_011_803);
  not1 I019_1037(w_019_1037, w_014_194);
  and2 I019_1040(w_019_1040, w_004_1689, w_007_697);
  not1 I019_1048(w_019_1048, w_001_1216);
  and2 I019_1057(w_019_1057, w_018_235, w_006_063);
  nand2 I019_1059(w_019_1059, w_002_497, w_002_198);
  nand2 I019_1060(w_019_1060, w_006_295, w_016_034);
  or2  I019_1070(w_019_1070, w_014_209, w_005_1424);
  not1 I019_1073(w_019_1073, w_003_297);
  and2 I019_1074(w_019_1074, w_017_1839, w_016_016);
  and2 I019_1082(w_019_1082, w_006_207, w_005_1219);
  not1 I019_1084(w_019_1084, w_008_261);
  nand2 I019_1085(w_019_1085, w_014_087, w_012_036);
  nand2 I019_1086(w_019_1086, w_006_271, w_015_214);
  or2  I019_1089(w_019_1089, w_012_122, w_000_700);
  and2 I019_1097(w_019_1097, w_004_056, w_006_146);
  or2  I020_007(w_020_007, w_008_463, w_003_224);
  or2  I020_014(w_020_014, w_012_372, w_013_272);
  nand2 I020_015(w_020_015, w_009_028, w_006_310);
  not1 I020_017(w_020_017, w_016_016);
  and2 I020_020(w_020_020, w_017_1288, w_008_355);
  nand2 I020_028(w_020_028, w_015_030, w_014_360);
  and2 I020_029(w_020_029, w_001_772, w_011_811);
  nand2 I020_030(w_020_030, w_019_089, w_000_736);
  nand2 I020_032(w_020_032, w_014_024, w_006_339);
  nand2 I020_039(w_020_039, w_008_285, w_001_589);
  nand2 I020_041(w_020_041, w_017_398, w_015_081);
  nand2 I020_045(w_020_045, w_006_300, w_016_010);
  and2 I020_063(w_020_063, w_006_063, w_014_008);
  not1 I020_064(w_020_064, w_011_635);
  nand2 I020_068(w_020_068, w_009_021, w_018_017);
  and2 I020_074(w_020_074, w_006_258, w_001_1496);
  not1 I020_075(w_020_075, w_014_666);
  not1 I020_085(w_020_085, w_011_150);
  and2 I020_092(w_020_092, w_014_473, w_005_144);
  nand2 I020_093(w_020_093, w_012_157, w_012_027);
  nand2 I020_096(w_020_096, w_010_038, w_019_167);
  nand2 I020_106(w_020_106, w_011_026, w_000_879);
  or2  I020_107(w_020_107, w_009_023, w_004_1187);
  and2 I020_111(w_020_111, w_008_248, w_001_020);
  nand2 I020_112(w_020_112, w_000_1819, w_011_619);
  or2  I020_114(w_020_114, w_011_815, w_018_054);
  nand2 I020_116(w_020_116, w_014_422, w_001_1632);
  or2  I020_117(w_020_117, w_006_275, w_009_014);
  or2  I020_121(w_020_121, w_003_108, w_000_387);
  not1 I020_123(w_020_123, w_001_201);
  and2 I020_133(w_020_133, w_018_088, w_019_115);
  not1 I020_134(w_020_134, w_004_1840);
  nand2 I020_135(w_020_135, w_015_006, w_011_428);
  nand2 I020_138(w_020_138, w_007_555, w_015_002);
  and2 I020_139(w_020_139, w_008_233, w_011_676);
  not1 I020_151(w_020_151, w_015_192);
  and2 I020_152(w_020_152, w_017_194, w_010_330);
  and2 I020_154(w_020_154, w_002_267, w_010_245);
  or2  I020_160(w_020_160, w_015_171, w_006_305);
  not1 I020_162(w_020_162, w_008_594);
  nand2 I020_164(w_020_164, w_005_1197, w_007_115);
  or2  I020_171(w_020_171, w_011_209, w_005_1426);
  or2  I020_174(w_020_174, w_012_573, w_014_237);
  and2 I020_176(w_020_176, w_012_039, w_014_072);
  nand2 I020_178(w_020_178, w_002_426, w_004_1781);
  nand2 I020_182(w_020_182, w_010_275, w_016_010);
  or2  I020_183(w_020_183, w_002_351, w_003_114);
  not1 I020_191(w_020_191, w_003_130);
  nand2 I020_193(w_020_193, w_006_320, w_014_809);
  nand2 I020_196(w_020_196, w_013_156, w_008_739);
  not1 I020_201(w_020_201, w_012_525);
  not1 I020_203(w_020_203, w_000_832);
  not1 I020_204(w_020_204, w_019_385);
  and2 I020_209(w_020_209, w_015_137, w_007_1078);
  and2 I020_210(w_020_210, w_010_208, w_012_538);
  or2  I020_217(w_020_217, w_005_1149, w_010_315);
  nand2 I020_219(w_020_219, w_003_290, w_006_325);
  nand2 I020_220(w_020_220, w_019_831, w_018_073);
  and2 I020_227(w_020_227, w_012_218, w_018_132);
  or2  I020_228(w_020_228, w_011_757, w_001_041);
  or2  I020_229(w_020_229, w_003_000, w_001_1186);
  nand2 I020_231(w_020_231, w_018_227, w_001_897);
  not1 I020_239(w_020_239, w_007_628);
  not1 I020_240(w_020_240, w_012_364);
  and2 I020_243(w_020_243, w_012_384, w_017_002);
  nand2 I020_244(w_020_244, w_012_454, w_006_104);
  not1 I020_249(w_020_249, w_019_499);
  not1 I020_250(w_020_250, w_011_135);
  or2  I020_252(w_020_252, w_008_058, w_018_161);
  or2  I020_256(w_020_256, w_017_034, w_011_667);
  or2  I020_265(w_020_265, w_000_1745, w_017_047);
  and2 I020_269(w_020_269, w_009_036, w_005_912);
  not1 I020_274(w_020_274, w_000_851);
  not1 I020_277(w_020_277, w_016_023);
  nand2 I020_278(w_020_278, w_001_1302, w_006_184);
  not1 I020_286(w_020_286, w_000_501);
  nand2 I020_288(w_020_288, w_013_270, w_015_023);
  or2  I020_289(w_020_289, w_017_562, w_019_302);
  or2  I020_290(w_020_290, w_010_224, w_014_293);
  not1 I020_292(w_020_292, w_003_258);
  or2  I020_293(w_020_293, w_005_1652, w_018_206);
  or2  I020_295(w_020_295, w_001_1301, w_002_423);
  nand2 I020_296(w_020_296, w_002_420, w_012_388);
  not1 I020_298(w_020_298, w_016_009);
  and2 I020_301(w_020_301, w_005_1424, w_018_091);
  not1 I020_304(w_020_304, w_010_211);
  and2 I020_305(w_020_305, w_019_504, w_001_1462);
  nand2 I020_308(w_020_308, w_009_024, w_016_018);
  nand2 I020_312(w_020_312, w_009_000, w_016_007);
  and2 I020_314(w_020_314, w_009_036, w_016_035);
  or2  I020_315(w_020_315, w_007_713, w_008_025);
  nand2 I020_317(w_020_317, w_008_662, w_005_1536);
  nand2 I020_323(w_020_323, w_019_361, w_019_627);
  nand2 I020_325(w_020_325, w_009_040, w_017_1031);
  or2  I020_327(w_020_327, w_010_090, w_009_063);
  not1 I020_330(w_020_330, w_013_325);
  or2  I020_332(w_020_332, w_009_042, w_019_298);
  nand2 I020_333(w_020_333, w_005_1140, w_012_171);
  nand2 I020_338(w_020_338, w_009_079, w_018_082);
  nand2 I020_342(w_020_342, w_010_014, w_017_1241);
  or2  I020_343(w_020_343, w_013_111, w_003_267);
  nand2 I020_348(w_020_348, w_010_131, w_005_1662);
  and2 I020_350(w_020_350, w_015_002, w_006_329);
  and2 I020_351(w_020_351, w_017_084, w_015_135);
  or2  I020_354(w_020_354, w_014_588, w_012_356);
  or2  I020_355(w_020_355, w_009_019, w_004_554);
  not1 I020_358(w_020_358, w_000_405);
  nand2 I020_359(w_020_359, w_004_1231, w_004_206);
  not1 I020_360(w_020_360, w_016_029);
  not1 I020_366(w_020_366, w_011_832);
  or2  I020_369(w_020_369, w_013_109, w_016_014);
  not1 I020_371(w_020_371, w_000_1086);
  nand2 I020_373(w_020_373, w_007_1077, w_017_1715);
  not1 I020_375(w_020_375, w_009_080);
  and2 I020_376(w_020_376, w_012_029, w_002_095);
  nand2 I020_377(w_020_377, w_004_011, w_006_178);
  and2 I020_379(w_020_379, w_001_1108, w_004_056);
  nand2 I020_381(w_020_381, w_012_061, w_001_031);
  not1 I020_383(w_020_383, w_001_090);
  nand2 I020_385(w_020_385, w_006_031, w_003_287);
  or2  I020_387(w_020_387, w_010_153, w_012_122);
  not1 I020_388(w_020_388, w_014_196);
  not1 I020_395(w_020_395, w_005_263);
  and2 I020_397(w_020_397, w_007_689, w_000_517);
  not1 I020_399(w_020_399, w_006_140);
  nand2 I020_401(w_020_401, w_002_217, w_016_001);
  and2 I020_404(w_020_404, w_016_004, w_016_018);
  or2  I020_405(w_020_405, w_011_718, w_016_029);
  not1 I020_416(w_020_416, w_014_533);
  or2  I020_422(w_020_422, w_014_094, w_008_163);
  and2 I020_423(w_020_423, w_014_426, w_017_1070);
  not1 I020_430(w_020_430, w_003_273);
  not1 I020_431(w_020_431, w_016_017);
  and2 I020_439(w_020_439, w_017_1421, w_011_094);
  or2  I020_440(w_020_440, w_018_201, w_003_243);
  nand2 I020_441(w_020_441, w_006_283, w_012_618);
  or2  I020_445(w_020_445, w_015_105, w_001_1284);
  not1 I020_448(w_020_448, w_012_133);
  not1 I020_449(w_020_449, w_002_324);
  or2  I020_452(w_020_452, w_014_723, w_014_167);
  nand2 I020_453(w_020_453, w_019_1082, w_017_155);
  nand2 I020_456(w_020_456, w_011_715, w_013_335);
  and2 I020_457(w_020_457, w_004_1682, w_019_082);
  or2  I020_460(w_020_460, w_018_144, w_013_172);
  or2  I020_464(w_020_464, w_009_036, w_011_453);
  not1 I020_465(w_020_465, w_016_012);
  or2  I020_466(w_020_466, w_015_033, w_007_1206);
  and2 I020_469(w_020_469, w_003_148, w_018_231);
  not1 I020_473(w_020_473, w_019_279);
  nand2 I020_476(w_020_476, w_000_174, w_010_160);
  not1 I020_478(w_020_478, w_001_174);
  and2 I020_480(w_020_480, w_009_082, w_011_057);
  not1 I020_483(w_020_483, w_001_1083);
  not1 I020_485(w_020_485, w_005_1636);
  nand2 I020_487(w_020_487, w_006_185, w_012_052);
  and2 I020_488(w_020_488, w_005_1581, w_007_1257);
  nand2 I020_490(w_020_490, w_016_005, w_008_739);
  not1 I020_493(w_020_493, w_017_1588);
  or2  I020_494(w_020_494, w_004_469, w_006_284);
  and2 I020_498(w_020_498, w_014_543, w_013_212);
  nand2 I020_500(w_020_500, w_000_503, w_001_1636);
  and2 I020_503(w_020_503, w_003_008, w_011_861);
  not1 I020_507(w_020_507, w_016_005);
  nand2 I020_510(w_020_510, w_004_1811, w_014_261);
  and2 I020_516(w_020_516, w_009_051, w_012_567);
  and2 I020_517(w_020_517, w_015_024, w_008_061);
  not1 I020_518(w_020_518, w_013_203);
  or2  I020_519(w_020_519, w_012_460, w_011_791);
  nand2 I020_520(w_020_520, w_002_034, w_019_552);
  or2  I020_521(w_020_521, w_018_110, w_001_989);
  not1 I020_525(w_020_525, w_018_269);
  and2 I020_527(w_020_527, w_001_292, w_003_046);
  not1 I020_528(w_020_528, w_013_040);
  and2 I020_538(w_020_538, w_008_110, w_005_919);
  not1 I020_539(w_020_539, w_007_1515);
  or2  I020_544(w_020_544, w_014_590, w_014_573);
  not1 I020_545(w_020_545, w_014_716);
  and2 I020_546(w_020_546, w_013_147, w_003_189);
  or2  I020_549(w_020_549, w_019_209, w_019_601);
  nand2 I020_551(w_020_551, w_017_702, w_005_140);
  or2  I020_557(w_020_557, w_009_084, w_006_275);
  not1 I020_559(w_020_559, w_015_224);
  not1 I020_569(w_020_569, w_016_010);
  and2 I020_572(w_020_572, w_014_641, w_016_019);
  and2 I020_573(w_020_573, w_018_265, w_019_575);
  not1 I020_579(w_020_579, w_001_418);
  nand2 I020_581(w_020_581, w_004_1749, w_005_094);
  nand2 I020_582(w_020_582, w_014_157, w_019_1086);
  not1 I020_583(w_020_583, w_011_619);
  or2  I020_585(w_020_585, w_016_037, w_002_360);
  not1 I020_589(w_020_589, w_007_1500);
  nand2 I020_591(w_020_591, w_014_402, w_014_502);
  nand2 I020_593(w_020_593, w_017_1396, w_009_096);
  and2 I020_597(w_020_597, w_016_030, w_019_122);
  or2  I020_598(w_020_598, w_005_050, w_017_1727);
  or2  I020_599(w_020_599, w_011_273, w_016_010);
  and2 I020_603(w_020_603, w_019_1070, w_007_174);
  nand2 I020_606(w_020_606, w_016_013, w_011_757);
  nand2 I020_611(w_020_611, w_014_278, w_011_040);
  and2 I020_612(w_020_612, w_010_080, w_012_071);
  not1 I020_614(w_020_614, w_009_077);
  or2  I020_620(w_020_620, w_016_001, w_003_231);
  nand2 I020_622(w_020_622, w_014_014, w_019_845);
  not1 I020_628(w_020_628, w_000_490);
  or2  I020_629(w_020_629, w_014_663, w_018_243);
  or2  I020_630(w_020_630, w_013_285, w_007_1619);
  and2 I020_631(w_020_631, w_001_721, w_002_156);
  not1 I020_643(w_020_643, w_004_970);
  not1 I020_648(w_020_648, w_006_242);
  nand2 I020_649(w_020_649, w_006_288, w_011_685);
  nand2 I020_650(w_020_650, w_007_539, w_006_036);
  nand2 I020_651(w_020_651, w_003_025, w_004_000);
  not1 I020_652(w_020_652, w_017_665);
  and2 I020_658(w_020_658, w_010_346, w_012_112);
  or2  I020_659(w_020_659, w_012_650, w_003_197);
  or2  I020_662(w_020_662, w_014_722, w_013_028);
  or2  I020_663(w_020_663, w_000_1191, w_019_374);
  or2  I020_664(w_020_664, w_007_837, w_006_239);
  nand2 I020_667(w_020_667, w_009_035, w_003_040);
  nand2 I020_668(w_020_668, w_012_154, w_013_077);
  and2 I020_671(w_020_671, w_008_627, w_001_420);
  or2  I020_673(w_020_673, w_004_1865, w_004_746);
  or2  I020_674(w_020_674, w_007_1458, w_008_031);
  or2  I020_676(w_020_676, w_003_104, w_017_905);
  and2 I020_677(w_020_677, w_001_1105, w_000_1423);
  not1 I020_685(w_020_685, w_012_049);
  and2 I020_687(w_020_687, w_018_214, w_015_031);
  nand2 I020_692(w_020_692, w_017_896, w_001_1532);
  and2 I020_694(w_020_694, w_007_202, w_004_914);
  nand2 I020_696(w_020_696, w_013_156, w_017_1065);
  or2  I020_701(w_020_701, w_008_379, w_004_1417);
  not1 I020_714(w_020_714, w_013_183);
  nand2 I020_717(w_020_717, w_003_131, w_019_304);
  nand2 I020_720(w_020_720, w_011_081, w_001_627);
  and2 I020_722(w_020_722, w_011_551, w_008_049);
  and2 I020_727(w_020_727, w_013_035, w_014_300);
  not1 I020_730(w_020_730, w_011_573);
  or2  I020_734(w_020_734, w_017_016, w_010_272);
  not1 I020_742(w_020_742, w_002_537);
  not1 I020_745(w_020_745, w_012_143);
  and2 I020_746(w_020_746, w_010_099, w_006_109);
  or2  I020_750(w_020_750, w_004_615, w_002_218);
  and2 I020_752(w_020_752, w_008_421, w_000_1026);
  not1 I020_753(w_020_753, w_001_643);
  nand2 I020_755(w_020_755, w_016_027, w_004_436);
  nand2 I020_764(w_020_764, w_017_1497, w_004_1102);
  not1 I020_766(w_020_766, w_015_052);
  or2  I020_772(w_020_772, w_000_1556, w_008_017);
  not1 I020_776(w_020_776, w_015_042);
  nand2 I020_777(w_020_777, w_016_011, w_008_474);
  and2 I020_784(w_020_784, w_004_1516, w_008_158);
  and2 I020_792(w_020_792, w_013_266, w_019_374);
  or2  I020_793(w_020_793, w_019_387, w_005_093);
  nand2 I020_794(w_020_794, w_013_236, w_003_020);
  or2  I020_796(w_020_796, w_005_1353, w_014_056);
  not1 I020_806(w_020_806, w_009_044);
  or2  I020_808(w_020_808, w_017_1031, w_010_360);
  nand2 I020_811(w_020_811, w_018_148, w_000_515);
  and2 I020_821(w_020_821, w_018_207, w_004_527);
  or2  I020_830(w_020_830, w_016_037, w_001_783);
  nand2 I020_839(w_020_839, w_009_006, w_018_160);
  or2  I020_842(w_020_842, w_009_100, w_007_1087);
  not1 I020_843(w_020_843, w_007_421);
  nand2 I020_846(w_020_846, w_017_038, w_001_1199);
  nand2 I020_857(w_020_857, w_017_393, w_013_115);
  and2 I020_858(w_020_858, w_012_250, w_013_178);
  and2 I020_860(w_020_860, w_013_207, w_004_080);
  and2 I020_867(w_020_867, w_005_466, w_004_1132);
  and2 I020_869(w_020_869, w_017_704, w_010_248);
  or2  I020_870(w_020_870, w_010_026, w_006_141);
  or2  I020_875(w_020_875, w_017_018, w_005_1134);
  not1 I020_880(w_020_880, w_008_207);
  and2 I020_886(w_020_886, w_007_035, w_001_639);
  not1 I020_887(w_020_887, w_005_873);
  and2 I020_892(w_020_892, w_007_085, w_001_235);
  and2 I020_895(w_020_895, w_010_045, w_008_252);
  not1 I020_897(w_020_897, w_015_155);
  not1 I020_905(w_020_905, w_016_029);
  or2  I020_915(w_020_915, w_015_097, w_006_228);
  not1 I020_922(w_020_922, w_000_1410);
  or2  I020_923(w_020_923, w_002_445, w_017_1460);
  and2 I020_924(w_020_924, w_019_246, w_015_077);
  not1 I020_929(w_020_929, w_013_309);
  or2  I020_934(w_020_934, w_016_015, w_004_1810);
  and2 I020_937(w_020_937, w_011_875, w_018_137);
  nand2 I020_939(w_020_939, w_005_005, w_015_183);
  or2  I020_941(w_020_941, w_002_030, w_007_1244);
  and2 I020_946(w_020_946, w_001_909, w_000_1347);
  not1 I020_949(w_020_949, w_003_296);
  nand2 I020_951(w_020_951, w_014_258, w_006_238);
  nand2 I020_961(w_020_961, w_003_045, w_001_294);
  and2 I020_976(w_020_976, w_014_453, w_006_006);
  and2 I020_979(w_020_979, w_012_139, w_000_1438);
  and2 I020_981(w_020_981, w_007_353, w_016_006);
  nand2 I020_983(w_020_983, w_000_1407, w_002_199);
  nand2 I020_986(w_020_986, w_010_304, w_005_546);
  and2 I020_989(w_020_989, w_019_756, w_011_003);
  or2  I020_991(w_020_991, w_001_492, w_011_871);
  and2 I020_993(w_020_993, w_001_377, w_002_095);
  not1 I020_994(w_020_994, w_002_497);
  or2  I020_995(w_020_995, w_015_200, w_017_1866);
  nand2 I020_1001(w_020_1001, w_014_411, w_019_909);
  nand2 I020_1017(w_020_1017, w_004_007, w_003_078);
  and2 I020_1020(w_020_1020, w_002_278, w_007_1276);
  not1 I020_1021(w_020_1021, w_018_057);
  nand2 I020_1030(w_020_1030, w_016_030, w_018_145);
  nand2 I020_1038(w_020_1038, w_004_921, w_004_027);
  nand2 I020_1040(w_020_1040, w_007_747, w_005_156);
  not1 I020_1043(w_020_1043, w_003_079);
  not1 I020_1053(w_020_1053, w_009_044);
  and2 I020_1060(w_020_1060, w_006_190, w_005_069);
  or2  I020_1062(w_020_1062, w_007_1402, w_000_098);
  or2  I020_1063(w_020_1063, w_016_036, w_018_195);
  or2  I020_1068(w_020_1068, w_019_553, w_010_358);
  and2 I020_1072(w_020_1072, w_003_284, w_013_227);
  nand2 I020_1084(w_020_1084, w_012_582, w_011_010);
  or2  I020_1085(w_020_1085, w_005_768, w_011_232);
  not1 I020_1091(w_020_1091, w_016_023);
  not1 I020_1095(w_020_1095, w_012_564);
  and2 I020_1097(w_020_1097, w_002_089, w_008_065);
  not1 I020_1108(w_020_1108, w_011_006);
  not1 I020_1115(w_020_1115, w_002_158);
  not1 I020_1120(w_020_1120, w_005_1080);
  nand2 I020_1121(w_020_1121, w_014_807, w_003_231);
  and2 I020_1125(w_020_1125, w_005_850, w_005_1044);
  not1 I020_1129(w_020_1129, w_011_077);
  nand2 I020_1131(w_020_1131, w_012_137, w_014_108);
  nand2 I020_1139(w_020_1139, w_019_568, w_014_520);
  and2 I020_1143(w_020_1143, w_009_059, w_001_1158);
  nand2 I020_1144(w_020_1144, w_014_072, w_006_257);
  or2  I020_1147(w_020_1147, w_001_102, w_003_213);
  nand2 I020_1151(w_020_1151, w_017_141, w_004_1687);
  and2 I020_1155(w_020_1155, w_006_125, w_004_1682);
  or2  I020_1163(w_020_1163, w_009_046, w_010_236);
  not1 I020_1166(w_020_1166, w_006_282);
  nand2 I020_1176(w_020_1176, w_009_064, w_014_027);
  nand2 I020_1189(w_020_1189, w_018_161, w_018_028);
  nand2 I020_1191(w_020_1191, w_017_1244, w_012_430);
  and2 I020_1194(w_020_1194, w_013_109, w_012_172);
  nand2 I020_1196(w_020_1196, w_016_031, w_005_1118);
  not1 I020_1198(w_020_1198, w_008_230);
  nand2 I020_1202(w_020_1202, w_012_106, w_014_276);
  not1 I020_1215(w_020_1215, w_015_141);
  and2 I020_1219(w_020_1219, w_012_077, w_003_079);
  nand2 I020_1222(w_020_1222, w_001_084, w_011_565);
  not1 I020_1225(w_020_1225, w_007_967);
  nand2 I020_1235(w_020_1235, w_011_718, w_015_048);
  not1 I020_1245(w_020_1245, w_017_903);
  not1 I020_1255(w_020_1255, w_011_856);
  nand2 I020_1258(w_020_1258, w_011_398, w_014_003);
  or2  I020_1263(w_020_1263, w_005_1283, w_008_456);
  and2 I020_1265(w_020_1265, w_001_1268, w_007_330);
  not1 I021_000(w_021_000, w_010_122);
  or2  I021_001(w_021_001, w_004_229, w_010_168);
  or2  I021_002(w_021_002, w_001_1226, w_018_110);
  not1 I021_003(w_021_003, w_020_017);
  or2  I021_005(w_021_005, w_004_979, w_003_319);
  and2 I021_006(w_021_006, w_013_038, w_012_085);
  and2 I021_007(w_021_007, w_001_1159, w_007_292);
  not1 I021_009(w_021_009, w_020_014);
  and2 I021_010(w_021_010, w_020_934, w_009_021);
  nand2 I021_011(w_021_011, w_014_243, w_002_020);
  not1 I021_013(w_021_013, w_017_932);
  and2 I021_015(w_021_015, w_020_171, w_017_002);
  and2 I021_016(w_021_016, w_006_308, w_020_1196);
  and2 I021_018(w_021_018, w_014_392, w_015_188);
  and2 I021_019(w_021_019, w_011_350, w_010_034);
  or2  I021_020(w_021_020, w_006_011, w_005_849);
  nand2 I021_021(w_021_021, w_017_1111, w_015_209);
  not1 I021_022(w_021_022, w_018_281);
  not1 I021_023(w_021_023, w_017_326);
  not1 I021_024(w_021_024, w_010_079);
  not1 I021_025(w_021_025, w_004_039);
  nand2 I021_026(w_021_026, w_010_403, w_015_052);
  and2 I021_027(w_021_027, w_003_289, w_005_159);
  nand2 I021_028(w_021_028, w_006_042, w_002_555);
  and2 I021_033(w_021_033, w_013_149, w_005_331);
  not1 I021_034(w_021_034, w_010_097);
  or2  I021_035(w_021_035, w_014_632, w_007_1295);
  not1 I021_036(w_021_036, w_000_938);
  or2  I021_037(w_021_037, w_005_858, w_010_188);
  or2  I021_041(w_021_041, w_001_1106, w_001_1457);
  not1 I021_042(w_021_042, w_008_752);
  or2  I021_044(w_021_044, w_012_626, w_003_170);
  not1 I021_045(w_021_045, w_006_024);
  not1 I021_046(w_021_046, w_017_975);
  or2  I021_047(w_021_047, w_005_1619, w_020_092);
  and2 I021_048(w_021_048, w_018_269, w_017_1893);
  and2 I021_049(w_021_049, w_011_215, w_005_1114);
  and2 I021_050(w_021_050, w_011_272, w_001_742);
  or2  I021_051(w_021_051, w_013_008, w_012_216);
  and2 I021_053(w_021_053, w_012_591, w_019_563);
  nand2 I021_054(w_021_054, w_016_001, w_000_366);
  or2  I021_055(w_021_055, w_015_023, w_015_150);
  not1 I021_057(w_021_057, w_010_392);
  and2 I021_058(w_021_058, w_011_064, w_003_116);
  nand2 I021_060(w_021_060, w_003_017, w_019_723);
  and2 I021_061(w_021_061, w_014_831, w_002_502);
  and2 I021_063(w_021_063, w_020_630, w_018_183);
  and2 I021_064(w_021_064, w_008_129, w_012_372);
  and2 I021_065(w_021_065, w_009_013, w_002_553);
  nand2 I021_066(w_021_066, w_001_1613, w_008_126);
  not1 I021_068(w_021_068, w_001_065);
  and2 I021_069(w_021_069, w_003_223, w_005_1278);
  or2  I021_071(w_021_071, w_010_149, w_012_494);
  not1 I021_072(w_021_072, w_012_067);
  or2  I021_073(w_021_073, w_011_700, w_019_754);
  or2  I021_074(w_021_074, w_008_205, w_010_178);
  and2 I021_075(w_021_075, w_011_553, w_007_1502);
  or2  I021_076(w_021_076, w_012_464, w_018_119);
  or2  I021_077(w_021_077, w_016_009, w_005_599);
  or2  I021_078(w_021_078, w_017_429, w_020_063);
  and2 I021_079(w_021_079, w_011_058, w_017_1262);
  and2 I021_080(w_021_080, w_013_252, w_000_867);
  and2 I021_081(w_021_081, w_013_001, w_015_285);
  nand2 I021_082(w_021_082, w_018_031, w_016_004);
  not1 I021_083(w_021_083, w_016_010);
  not1 I021_084(w_021_084, w_001_1585);
  nand2 I021_085(w_021_085, w_016_014, w_015_030);
  nand2 I021_086(w_021_086, w_005_1384, w_000_1118);
  and2 I021_087(w_021_087, w_013_010, w_001_573);
  nand2 I021_088(w_021_088, w_012_598, w_011_203);
  or2  I021_089(w_021_089, w_008_270, w_002_556);
  or2  I021_090(w_021_090, w_018_165, w_002_171);
  and2 I021_091(w_021_091, w_017_502, w_004_1578);
  and2 I021_092(w_021_092, w_010_171, w_012_314);
  or2  I021_093(w_021_093, w_011_020, w_011_782);
  or2  I021_094(w_021_094, w_007_1234, w_014_055);
  not1 I021_095(w_021_095, w_019_710);
  or2  I021_096(w_021_096, w_000_1556, w_010_086);
  nand2 I021_097(w_021_097, w_012_288, w_006_338);
  not1 I021_099(w_021_099, w_018_108);
  not1 I021_100(w_021_100, w_003_016);
  not1 I021_101(w_021_101, w_001_263);
  and2 I021_102(w_021_102, w_012_238, w_008_477);
  or2  I021_103(w_021_103, w_018_165, w_009_097);
  not1 I021_104(w_021_104, w_013_236);
  nand2 I021_105(w_021_105, w_001_890, w_006_219);
  not1 I021_107(w_021_107, w_001_1681);
  not1 I021_111(w_021_111, w_009_067);
  or2  I021_112(w_021_112, w_008_750, w_007_1468);
  not1 I021_115(w_021_115, w_008_108);
  or2  I021_116(w_021_116, w_003_039, w_003_316);
  or2  I021_117(w_021_117, w_011_091, w_012_006);
  nand2 I021_118(w_021_118, w_002_552, w_018_249);
  not1 I021_119(w_021_119, w_005_173);
  not1 I021_120(w_021_120, w_019_514);
  or2  I021_122(w_021_122, w_020_075, w_006_126);
  or2  I021_123(w_021_123, w_007_1502, w_006_340);
  nand2 I021_124(w_021_124, w_015_062, w_009_037);
  and2 I021_126(w_021_126, w_017_006, w_002_273);
  or2  I021_128(w_021_128, w_019_105, w_013_053);
  nand2 I021_129(w_021_129, w_016_018, w_015_031);
  not1 I021_130(w_021_130, w_012_163);
  or2  I021_132(w_021_132, w_006_166, w_015_293);
  or2  I021_134(w_021_134, w_002_579, w_013_038);
  and2 I021_135(w_021_135, w_000_1328, w_012_227);
  or2  I021_136(w_021_136, w_015_059, w_011_347);
  and2 I021_137(w_021_137, w_010_295, w_016_017);
  nand2 I021_138(w_021_138, w_014_150, w_012_122);
  and2 I021_139(w_021_139, w_004_768, w_009_073);
  and2 I021_140(w_021_140, w_020_685, w_005_187);
  not1 I021_141(w_021_141, w_019_978);
  not1 I021_142(w_021_142, w_010_225);
  nand2 I021_143(w_021_143, w_002_048, w_015_213);
  or2  I021_144(w_021_144, w_003_180, w_001_1130);
  and2 I021_145(w_021_145, w_013_112, w_006_292);
  and2 I021_147(w_021_147, w_015_209, w_003_283);
  nand2 I021_148(w_021_148, w_001_1613, w_010_303);
  nand2 I021_149(w_021_149, w_014_403, w_005_960);
  not1 I021_150(w_021_150, w_011_357);
  not1 I021_151(w_021_151, w_010_155);
  nand2 I021_153(w_021_153, w_012_281, w_010_234);
  or2  I021_154(w_021_154, w_010_029, w_001_513);
  or2  I021_155(w_021_155, w_005_548, w_020_1194);
  not1 I021_156(w_021_156, w_008_168);
  and2 I021_157(w_021_157, w_018_209, w_007_1211);
  or2  I021_158(w_021_158, w_019_470, w_003_000);
  and2 I021_159(w_021_159, w_002_396, w_006_235);
  nand2 I021_161(w_021_161, w_011_816, w_008_612);
  and2 I021_162(w_021_162, w_007_182, w_008_526);
  nand2 I021_163(w_021_163, w_006_267, w_012_375);
  nand2 I021_166(w_021_166, w_015_106, w_014_005);
  nand2 I021_167(w_021_167, w_002_200, w_001_742);
  and2 I021_169(w_021_169, w_004_1402, w_016_011);
  or2  I021_171(w_021_171, w_013_325, w_016_035);
  not1 I021_172(w_021_172, w_017_040);
  not1 I021_174(w_021_174, w_001_1599);
  and2 I021_177(w_021_177, w_006_093, w_018_104);
  not1 I021_179(w_021_179, w_009_070);
  or2  I021_180(w_021_180, w_017_1092, w_002_137);
  or2  I021_182(w_021_182, w_001_193, w_006_076);
  nand2 I021_184(w_021_184, w_009_067, w_004_1686);
  not1 I021_185(w_021_185, w_013_025);
  not1 I021_186(w_021_186, w_005_535);
  not1 I021_187(w_021_187, w_017_1924);
  or2  I021_189(w_021_189, w_006_310, w_019_161);
  or2  I021_191(w_021_191, w_017_244, w_000_988);
  or2  I021_193(w_021_193, w_015_184, w_017_1374);
  and2 I021_194(w_021_194, w_002_018, w_019_701);
  and2 I021_195(w_021_195, w_016_004, w_000_335);
  and2 I021_198(w_021_198, w_012_402, w_009_035);
  nand2 I021_199(w_021_199, w_012_399, w_015_190);
  not1 I021_201(w_021_201, w_015_086);
  or2  I021_202(w_021_202, w_016_037, w_001_1383);
  or2  I021_203(w_021_203, w_014_722, w_011_589);
  or2  I021_204(w_021_204, w_003_196, w_001_010);
  nand2 I021_205(w_021_205, w_008_519, w_001_877);
  nand2 I021_207(w_021_207, w_009_007, w_015_146);
  or2  I021_208(w_021_208, w_009_066, w_004_1693);
  nand2 I021_210(w_021_210, w_000_1060, w_011_161);
  and2 I021_211(w_021_211, w_011_213, w_017_1218);
  and2 I021_212(w_021_212, w_016_017, w_020_614);
  nand2 I021_214(w_021_214, w_019_329, w_001_1200);
  and2 I021_216(w_021_216, w_002_408, w_010_124);
  or2  I021_218(w_021_218, w_018_282, w_013_134);
  and2 I021_220(w_021_220, w_004_1051, w_005_860);
  nand2 I021_221(w_021_221, w_002_514, w_000_608);
  and2 I021_223(w_021_223, w_002_405, w_016_006);
  or2  I021_224(w_021_224, w_014_051, w_013_016);
  not1 I021_225(w_021_225, w_005_251);
  or2  I021_226(w_021_226, w_014_143, w_000_1020);
  not1 I021_227(w_021_227, w_005_232);
  not1 I021_228(w_021_228, w_005_259);
  not1 I021_229(w_021_229, w_010_239);
  and2 I021_231(w_021_231, w_016_028, w_006_169);
  nand2 I021_232(w_021_232, w_014_032, w_001_1629);
  not1 I021_233(w_021_233, w_018_011);
  and2 I021_234(w_021_234, w_013_296, w_010_221);
  or2  I021_235(w_021_235, w_011_414, w_011_631);
  and2 I021_236(w_021_236, w_019_106, w_007_149);
  and2 I021_237(w_021_237, w_001_710, w_010_029);
  or2  I021_238(w_021_238, w_017_417, w_003_151);
  or2  I021_239(w_021_239, w_002_592, w_012_219);
  not1 I021_240(w_021_240, w_003_232);
  nand2 I021_241(w_021_241, w_013_328, w_014_696);
  not1 I021_242(w_021_242, w_003_083);
  or2  I021_244(w_021_244, w_013_091, w_003_269);
  and2 I021_245(w_021_245, w_020_286, w_000_1544);
  nand2 I021_246(w_021_246, w_002_488, w_006_277);
  not1 I021_248(w_021_248, w_016_002);
  or2  I021_249(w_021_249, w_017_1308, w_012_000);
  or2  I021_250(w_021_250, w_003_065, w_019_615);
  and2 I021_251(w_021_251, w_000_1585, w_001_1345);
  not1 I021_253(w_021_253, w_002_446);
  or2  I021_254(w_021_254, w_010_308, w_009_004);
  not1 I021_255(w_021_255, w_003_173);
  nand2 I021_256(w_021_256, w_020_527, w_008_222);
  nand2 I021_257(w_021_257, w_012_259, w_017_366);
  nand2 I021_258(w_021_258, w_017_303, w_004_575);
  not1 I021_259(w_021_259, w_004_1817);
  and2 I021_260(w_021_260, w_006_056, w_002_240);
  or2  I021_261(w_021_261, w_011_016, w_000_383);
  nand2 I021_262(w_021_262, w_003_236, w_006_273);
  not1 I021_263(w_021_263, w_015_224);
  not1 I021_264(w_021_264, w_006_127);
  and2 I021_265(w_021_265, w_010_235, w_017_805);
  nand2 I021_266(w_021_266, w_010_420, w_011_715);
  and2 I021_268(w_021_268, w_008_751, w_003_129);
  nand2 I021_269(w_021_269, w_004_318, w_017_1718);
  and2 I021_270(w_021_270, w_009_038, w_013_180);
  or2  I021_271(w_021_271, w_015_244, w_000_1820);
  nand2 I021_272(w_021_272, w_005_1602, w_011_496);
  or2  I021_273(w_021_273, w_008_126, w_011_640);
  and2 I021_274(w_021_274, w_014_163, w_010_109);
  and2 I021_275(w_021_275, w_019_246, w_018_090);
  and2 I021_276(w_021_276, w_005_298, w_003_197);
  not1 I021_277(w_021_277, w_001_412);
  and2 I022_000(w_022_000, w_006_095, w_000_186);
  or2  I022_001(w_022_001, w_004_1739, w_006_060);
  nand2 I022_002(w_022_002, w_012_316, w_002_593);
  or2  I022_003(w_022_003, w_000_218, w_003_076);
  and2 I022_004(w_022_004, w_019_252, w_017_677);
  nand2 I022_005(w_022_005, w_007_187, w_019_888);
  and2 I022_007(w_022_007, w_003_212, w_013_313);
  or2  I022_008(w_022_008, w_005_1439, w_019_342);
  or2  I022_009(w_022_009, w_012_233, w_013_243);
  or2  I022_010(w_022_010, w_001_292, w_006_215);
  nand2 I022_011(w_022_011, w_002_230, w_002_363);
  or2  I022_012(w_022_012, w_011_217, w_004_819);
  or2  I022_013(w_022_013, w_020_030, w_016_016);
  and2 I022_015(w_022_015, w_012_195, w_001_543);
  not1 I022_016(w_022_016, w_016_011);
  or2  I022_018(w_022_018, w_003_140, w_016_008);
  nand2 I022_023(w_022_023, w_014_370, w_006_058);
  or2  I022_025(w_022_025, w_007_118, w_020_612);
  and2 I022_026(w_022_026, w_017_1067, w_012_508);
  not1 I022_027(w_022_027, w_009_074);
  and2 I022_028(w_022_028, w_020_549, w_017_1207);
  nand2 I022_029(w_022_029, w_006_267, w_008_685);
  or2  I022_030(w_022_030, w_012_316, w_003_191);
  and2 I022_031(w_022_031, w_007_225, w_004_1268);
  and2 I022_032(w_022_032, w_000_1507, w_000_979);
  nand2 I022_033(w_022_033, w_010_155, w_011_666);
  not1 I022_036(w_022_036, w_019_507);
  not1 I022_037(w_022_037, w_020_151);
  nand2 I022_038(w_022_038, w_005_001, w_011_213);
  or2  I022_039(w_022_039, w_011_837, w_013_258);
  nand2 I022_041(w_022_041, w_016_024, w_009_044);
  nand2 I022_042(w_022_042, w_020_808, w_003_313);
  not1 I022_043(w_022_043, w_020_593);
  not1 I022_045(w_022_045, w_020_312);
  nand2 I022_046(w_022_046, w_007_033, w_002_291);
  or2  I022_047(w_022_047, w_002_331, w_010_250);
  nand2 I022_051(w_022_051, w_006_206, w_014_417);
  not1 I022_053(w_022_053, w_008_470);
  not1 I022_054(w_022_054, w_001_1266);
  nand2 I022_055(w_022_055, w_020_182, w_000_1502);
  nand2 I022_056(w_022_056, w_002_302, w_010_256);
  not1 I022_057(w_022_057, w_005_444);
  not1 I022_058(w_022_058, w_002_003);
  and2 I022_059(w_022_059, w_019_507, w_001_473);
  and2 I022_060(w_022_060, w_021_099, w_017_1947);
  not1 I022_061(w_022_061, w_013_245);
  or2  I022_062(w_022_062, w_007_1141, w_004_704);
  not1 I022_064(w_022_064, w_001_601);
  and2 I022_066(w_022_066, w_012_594, w_011_877);
  not1 I022_067(w_022_067, w_010_417);
  or2  I022_068(w_022_068, w_006_191, w_018_226);
  and2 I022_069(w_022_069, w_003_174, w_012_146);
  not1 I022_070(w_022_070, w_021_042);
  or2  I022_072(w_022_072, w_021_263, w_011_123);
  nand2 I022_074(w_022_074, w_017_1008, w_014_076);
  or2  I022_075(w_022_075, w_018_192, w_021_095);
  nand2 I022_076(w_022_076, w_001_1508, w_012_067);
  and2 I022_078(w_022_078, w_001_157, w_011_678);
  not1 I022_079(w_022_079, w_021_246);
  or2  I022_081(w_022_081, w_016_034, w_011_328);
  not1 I022_083(w_022_083, w_014_427);
  and2 I022_084(w_022_084, w_001_1461, w_017_1060);
  or2  I022_085(w_022_085, w_018_085, w_008_125);
  or2  I022_088(w_022_088, w_000_440, w_009_099);
  nand2 I022_089(w_022_089, w_001_000, w_018_045);
  or2  I022_090(w_022_090, w_002_511, w_016_034);
  and2 I022_093(w_022_093, w_019_234, w_017_748);
  nand2 I022_094(w_022_094, w_013_282, w_018_078);
  or2  I022_096(w_022_096, w_009_032, w_006_196);
  and2 I022_097(w_022_097, w_017_891, w_004_058);
  or2  I022_098(w_022_098, w_012_097, w_011_504);
  and2 I022_099(w_022_099, w_003_264, w_015_019);
  and2 I022_101(w_022_101, w_015_204, w_008_447);
  or2  I022_103(w_022_103, w_015_038, w_010_226);
  or2  I022_104(w_022_104, w_020_796, w_000_191);
  and2 I022_105(w_022_105, w_002_354, w_010_073);
  not1 I022_107(w_022_107, w_004_1414);
  and2 I022_108(w_022_108, w_012_525, w_020_029);
  not1 I022_109(w_022_109, w_001_170);
  nand2 I022_111(w_022_111, w_010_035, w_000_1449);
  nand2 I022_113(w_022_113, w_010_204, w_006_123);
  and2 I022_114(w_022_114, w_008_225, w_017_1646);
  or2  I022_116(w_022_116, w_014_223, w_006_199);
  or2  I022_118(w_022_118, w_004_217, w_013_199);
  and2 I022_120(w_022_120, w_013_040, w_016_010);
  and2 I022_122(w_022_122, w_008_698, w_019_294);
  not1 I022_123(w_022_123, w_001_970);
  and2 I022_128(w_022_128, w_008_624, w_015_100);
  and2 I022_129(w_022_129, w_002_251, w_005_695);
  not1 I022_131(w_022_131, w_016_000);
  or2  I022_132(w_022_132, w_001_1509, w_014_483);
  not1 I022_133(w_022_133, w_009_110);
  not1 I022_135(w_022_135, w_021_229);
  nand2 I022_136(w_022_136, w_005_1597, w_019_273);
  not1 I022_137(w_022_137, w_020_152);
  or2  I022_139(w_022_139, w_008_343, w_005_1491);
  and2 I022_140(w_022_140, w_004_1437, w_021_076);
  and2 I022_141(w_022_141, w_014_662, w_007_269);
  and2 I022_142(w_022_142, w_006_155, w_010_330);
  and2 I022_143(w_022_143, w_005_967, w_021_238);
  not1 I022_144(w_022_144, w_004_478);
  and2 I022_146(w_022_146, w_008_394, w_000_014);
  or2  I022_148(w_022_148, w_004_1206, w_020_439);
  or2  I022_149(w_022_149, w_006_283, w_020_598);
  not1 I022_150(w_022_150, w_019_1019);
  not1 I022_152(w_022_152, w_018_216);
  not1 I022_153(w_022_153, w_005_042);
  nand2 I022_155(w_022_155, w_010_264, w_008_738);
  or2  I022_156(w_022_156, w_020_976, w_019_860);
  and2 I022_159(w_022_159, w_000_1935, w_016_003);
  or2  I022_161(w_022_161, w_017_1246, w_004_1546);
  nand2 I022_163(w_022_163, w_008_308, w_011_100);
  or2  I022_166(w_022_166, w_011_700, w_009_048);
  or2  I022_168(w_022_168, w_019_866, w_006_238);
  nand2 I022_169(w_022_169, w_019_278, w_012_426);
  and2 I022_171(w_022_171, w_021_078, w_013_271);
  not1 I022_172(w_022_172, w_006_297);
  nand2 I022_173(w_022_173, w_016_037, w_015_044);
  not1 I022_175(w_022_175, w_010_307);
  nand2 I022_177(w_022_177, w_012_227, w_003_286);
  not1 I022_178(w_022_178, w_012_343);
  and2 I022_179(w_022_179, w_008_851, w_021_018);
  not1 I022_181(w_022_181, w_015_170);
  not1 I022_182(w_022_182, w_009_102);
  not1 I022_184(w_022_184, w_002_239);
  not1 I022_185(w_022_185, w_006_329);
  or2  I022_186(w_022_186, w_010_356, w_014_470);
  or2  I022_188(w_022_188, w_006_276, w_017_203);
  and2 I022_194(w_022_194, w_005_1569, w_016_013);
  and2 I022_195(w_022_195, w_016_015, w_021_270);
  not1 I022_196(w_022_196, w_000_668);
  and2 I022_197(w_022_197, w_011_267, w_012_640);
  and2 I022_200(w_022_200, w_001_1228, w_002_286);
  and2 I022_201(w_022_201, w_005_801, w_004_907);
  or2  I022_202(w_022_202, w_019_404, w_018_065);
  not1 I022_203(w_022_203, w_018_167);
  not1 I022_204(w_022_204, w_007_803);
  not1 I022_206(w_022_206, w_002_442);
  not1 I022_208(w_022_208, w_013_299);
  nand2 I022_210(w_022_210, w_001_083, w_008_501);
  or2  I022_212(w_022_212, w_005_237, w_016_038);
  or2  I022_213(w_022_213, w_021_104, w_014_523);
  and2 I022_217(w_022_217, w_005_232, w_012_649);
  not1 I022_219(w_022_219, w_001_964);
  or2  I022_222(w_022_222, w_010_359, w_009_054);
  or2  I022_223(w_022_223, w_006_004, w_003_021);
  or2  I022_224(w_022_224, w_006_248, w_013_009);
  not1 I022_225(w_022_225, w_004_326);
  nand2 I022_227(w_022_227, w_001_1672, w_021_045);
  or2  I022_230(w_022_230, w_009_002, w_014_653);
  nand2 I022_231(w_022_231, w_019_085, w_014_032);
  nand2 I022_232(w_022_232, w_018_022, w_019_025);
  nand2 I022_233(w_022_233, w_005_1026, w_006_161);
  nand2 I022_234(w_022_234, w_005_1384, w_001_216);
  and2 I022_235(w_022_235, w_018_163, w_003_011);
  and2 I022_236(w_022_236, w_014_755, w_008_425);
  and2 I022_238(w_022_238, w_005_1281, w_007_360);
  and2 I022_244(w_022_244, w_017_1014, w_004_1622);
  and2 I022_246(w_022_246, w_005_1105, w_012_375);
  not1 I022_248(w_022_248, w_017_1729);
  nand2 I022_249(w_022_249, w_001_602, w_019_028);
  not1 I022_251(w_022_251, w_001_1628);
  not1 I022_254(w_022_254, w_015_191);
  or2  I022_262(w_022_262, w_018_211, w_012_326);
  nand2 I022_265(w_022_265, w_009_039, w_016_024);
  or2  I022_266(w_022_266, w_002_010, w_013_305);
  not1 I022_267(w_022_267, w_003_107);
  nand2 I022_268(w_022_268, w_009_011, w_011_791);
  or2  I022_275(w_022_275, w_012_413, w_017_691);
  or2  I022_277(w_022_277, w_018_257, w_007_1084);
  and2 I022_278(w_022_278, w_013_183, w_007_592);
  or2  I022_279(w_022_279, w_012_076, w_019_145);
  or2  I022_280(w_022_280, w_015_187, w_010_400);
  nand2 I022_281(w_022_281, w_017_088, w_004_1348);
  and2 I022_283(w_022_283, w_005_317, w_006_070);
  nand2 I022_286(w_022_286, w_021_202, w_008_584);
  and2 I022_287(w_022_287, w_018_135, w_003_078);
  or2  I022_289(w_022_289, w_003_138, w_007_1208);
  nand2 I022_290(w_022_290, w_014_662, w_003_255);
  or2  I022_293(w_022_293, w_004_703, w_001_1271);
  or2  I022_294(w_022_294, w_013_163, w_001_644);
  and2 I022_295(w_022_295, w_005_1189, w_004_950);
  or2  I022_296(w_022_296, w_021_072, w_018_049);
  nand2 I022_297(w_022_297, w_016_023, w_012_215);
  not1 I022_298(w_022_298, w_004_049);
  nand2 I022_300(w_022_300, w_012_269, w_006_224);
  not1 I022_302(w_022_302, w_009_039);
  nand2 I022_304(w_022_304, w_012_181, w_003_047);
  nand2 I022_305(w_022_305, w_005_049, w_018_018);
  or2  I022_306(w_022_306, w_007_997, w_000_1806);
  nand2 I022_307(w_022_307, w_004_1406, w_014_599);
  not1 I022_308(w_022_308, w_017_088);
  and2 I022_309(w_022_309, w_004_047, w_020_244);
  not1 I022_310(w_022_310, w_017_1348);
  or2  I022_311(w_022_311, w_007_865, w_017_1071);
  and2 I022_312(w_022_312, w_020_1120, w_000_718);
  nand2 I022_316(w_022_316, w_006_261, w_019_294);
  and2 I022_320(w_022_320, w_005_1624, w_009_053);
  nand2 I022_321(w_022_321, w_010_371, w_009_050);
  and2 I022_322(w_022_322, w_003_103, w_003_044);
  not1 I022_323(w_022_323, w_008_078);
  and2 I022_324(w_022_324, w_004_312, w_002_176);
  or2  I022_325(w_022_325, w_008_225, w_018_197);
  or2  I022_327(w_022_327, w_009_041, w_002_283);
  or2  I022_329(w_022_329, w_013_231, w_001_233);
  and2 I022_331(w_022_331, w_007_1592, w_020_673);
  and2 I022_332(w_022_332, w_014_218, w_020_676);
  or2  I022_335(w_022_335, w_011_193, w_018_091);
  nand2 I022_338(w_022_338, w_001_345, w_009_059);
  nand2 I022_339(w_022_339, w_005_570, w_001_849);
  nand2 I022_340(w_022_340, w_007_1366, w_009_042);
  or2  I022_341(w_022_341, w_021_236, w_007_656);
  nand2 I022_342(w_022_342, w_001_514, w_007_583);
  or2  I022_343(w_022_343, w_002_289, w_003_257);
  or2  I022_344(w_022_344, w_004_1362, w_014_613);
  not1 I022_346(w_022_346, w_015_230);
  and2 I022_347(w_022_347, w_000_721, w_010_270);
  nand2 I022_348(w_022_348, w_015_229, w_004_1320);
  or2  I022_349(w_022_349, w_009_032, w_020_951);
  or2  I022_353(w_022_353, w_021_174, w_007_253);
  nand2 I022_354(w_022_354, w_015_120, w_012_188);
  or2  I022_356(w_022_356, w_003_153, w_008_043);
  nand2 I022_362(w_022_362, w_004_074, w_012_488);
  or2  I022_365(w_022_365, w_018_056, w_021_101);
  not1 I022_367(w_022_367, w_006_057);
  or2  I022_368(w_022_368, w_004_1665, w_012_217);
  or2  I022_369(w_022_369, w_014_315, w_015_036);
  not1 I022_370(w_022_370, w_006_266);
  not1 I022_371(w_022_371, w_000_289);
  nand2 I022_373(w_022_373, w_014_318, w_008_156);
  nand2 I022_374(w_022_374, w_011_805, w_003_005);
  and2 I022_376(w_022_376, w_009_043, w_017_1878);
  and2 I022_377(w_022_377, w_013_073, w_012_059);
  nand2 I022_381(w_022_381, w_003_101, w_016_026);
  nand2 I022_382(w_022_382, w_013_165, w_013_300);
  and2 I022_383(w_022_383, w_008_346, w_004_830);
  not1 I022_385(w_022_385, w_006_022);
  or2  I022_386(w_022_386, w_013_182, w_015_206);
  nand2 I022_388(w_022_388, w_019_450, w_014_112);
  and2 I022_390(w_022_390, w_018_202, w_008_481);
  or2  I022_391(w_022_391, w_017_1047, w_018_242);
  or2  I022_392(w_022_392, w_013_064, w_015_074);
  not1 I022_393(w_022_393, w_017_1419);
  nand2 I022_395(w_022_395, w_005_993, w_000_595);
  not1 I022_397(w_022_397, w_009_013);
  not1 I022_398(w_022_398, w_018_209);
  or2  I022_399(w_022_399, w_009_030, w_017_1026);
  nand2 I022_400(w_022_400, w_007_961, w_004_596);
  and2 I022_401(w_022_401, w_003_068, w_016_037);
  and2 I022_402(w_022_402, w_005_924, w_005_832);
  and2 I022_403(w_022_403, w_014_439, w_011_173);
  or2  I022_404(w_022_404, w_019_225, w_006_107);
  or2  I022_405(w_022_405, w_001_752, w_017_254);
  nand2 I022_407(w_022_407, w_019_467, w_013_162);
  and2 I022_408(w_022_408, w_005_439, w_020_404);
  nand2 I022_409(w_022_409, w_002_048, w_009_086);
  nand2 I022_410(w_022_410, w_019_1048, w_009_094);
  nand2 I022_412(w_022_412, w_014_721, w_021_033);
  nand2 I022_413(w_022_413, w_014_673, w_016_030);
  or2  I022_414(w_022_414, w_007_121, w_015_064);
  not1 I022_416(w_022_416, w_020_399);
  not1 I022_417(w_022_417, w_017_1074);
  nand2 I022_418(w_022_418, w_011_033, w_014_252);
  and2 I022_420(w_022_420, w_019_724, w_020_792);
  nand2 I022_428(w_022_428, w_021_208, w_020_114);
  nand2 I022_430(w_022_430, w_018_231, w_001_505);
  nand2 I022_439(w_022_441, w_010_322, w_022_440);
  not1 I022_440(w_022_442, w_022_441);
  nand2 I022_441(w_022_443, w_009_009, w_022_442);
  nand2 I022_442(w_022_444, w_022_443, w_003_271);
  not1 I022_443(w_022_445, w_022_444);
  nand2 I022_444(w_022_446, w_022_445, w_011_011);
  not1 I022_445(w_022_447, w_022_446);
  and2 I022_446(w_022_440, w_022_447, w_018_200);
  and2 I022_447(w_022_452, w_009_129, w_022_451);
  nand2 I022_448(w_022_453, w_013_302, w_022_452);
  and2 I022_449(w_022_454, w_010_135, w_022_453);
  or2  I022_450(w_022_455, w_022_454, w_003_289);
  and2 I022_451(w_022_456, w_022_455, w_017_1231);
  nand2 I022_452(w_022_457, w_011_256, w_022_456);
  or2  I022_453(w_022_458, w_003_319, w_022_457);
  nand2 I022_454(w_022_459, w_015_048, w_022_458);
  or2  I022_455(w_022_451, w_010_295, w_022_459);
  and2 I023_003(w_023_003, w_019_994, w_020_620);
  or2  I023_004(w_023_004, w_001_006, w_004_1631);
  nand2 I023_009(w_023_009, w_017_1822, w_007_609);
  and2 I023_010(w_023_010, w_021_022, w_009_083);
  or2  I023_012(w_023_012, w_020_687, w_005_1674);
  not1 I023_013(w_023_013, w_015_049);
  not1 I023_019(w_023_019, w_007_873);
  nand2 I023_020(w_023_020, w_018_147, w_017_1391);
  nand2 I023_023(w_023_023, w_004_534, w_007_255);
  not1 I023_026(w_023_026, w_007_509);
  and2 I023_029(w_023_029, w_004_583, w_012_209);
  nand2 I023_039(w_023_039, w_018_194, w_021_194);
  or2  I023_040(w_023_040, w_015_021, w_000_104);
  or2  I023_043(w_023_043, w_003_151, w_013_077);
  and2 I023_045(w_023_045, w_018_048, w_000_564);
  and2 I023_046(w_023_046, w_015_122, w_008_443);
  not1 I023_049(w_023_049, w_015_143);
  or2  I023_060(w_023_060, w_003_040, w_005_1348);
  not1 I023_061(w_023_061, w_018_271);
  or2  I023_062(w_023_062, w_020_1245, w_010_047);
  or2  I023_064(w_023_064, w_004_1288, w_004_997);
  nand2 I023_065(w_023_065, w_019_671, w_004_1795);
  not1 I023_066(w_023_066, w_004_1714);
  nand2 I023_070(w_023_070, w_002_398, w_020_007);
  or2  I023_071(w_023_071, w_018_279, w_008_767);
  and2 I023_072(w_023_072, w_006_226, w_021_105);
  nand2 I023_076(w_023_076, w_002_173, w_019_124);
  or2  I023_077(w_023_077, w_000_1147, w_008_456);
  nand2 I023_088(w_023_088, w_001_121, w_002_004);
  and2 I023_091(w_023_091, w_012_435, w_009_104);
  or2  I023_093(w_023_093, w_013_035, w_022_054);
  and2 I023_097(w_023_097, w_021_080, w_015_094);
  and2 I023_100(w_023_100, w_002_236, w_017_1310);
  not1 I023_101(w_023_101, w_016_002);
  nand2 I023_111(w_023_111, w_019_1073, w_016_004);
  nand2 I023_114(w_023_114, w_017_1135, w_005_256);
  and2 I023_117(w_023_117, w_005_109, w_002_042);
  and2 I023_123(w_023_123, w_003_276, w_018_061);
  and2 I023_126(w_023_126, w_007_306, w_013_032);
  not1 I023_135(w_023_135, w_018_071);
  not1 I023_136(w_023_136, w_004_288);
  and2 I023_142(w_023_142, w_015_282, w_022_090);
  not1 I023_147(w_023_147, w_007_251);
  nand2 I023_154(w_023_154, w_018_280, w_000_460);
  nand2 I023_156(w_023_156, w_010_081, w_003_184);
  nand2 I023_157(w_023_157, w_013_033, w_022_062);
  or2  I023_158(w_023_158, w_002_322, w_000_1758);
  not1 I023_161(w_023_161, w_017_1937);
  not1 I023_169(w_023_169, w_003_110);
  nand2 I023_176(w_023_176, w_005_309, w_012_198);
  nand2 I023_180(w_023_180, w_003_105, w_000_730);
  or2  I023_181(w_023_181, w_008_772, w_000_678);
  or2  I023_187(w_023_187, w_007_559, w_017_1372);
  not1 I023_190(w_023_190, w_017_1497);
  nand2 I023_191(w_023_191, w_010_115, w_009_072);
  or2  I023_198(w_023_198, w_012_297, w_002_509);
  nand2 I023_199(w_023_199, w_001_176, w_001_1037);
  nand2 I023_204(w_023_204, w_013_189, w_002_474);
  not1 I023_205(w_023_205, w_004_524);
  not1 I023_206(w_023_206, w_006_012);
  and2 I023_211(w_023_211, w_016_028, w_017_1402);
  and2 I023_212(w_023_212, w_014_256, w_018_087);
  not1 I023_213(w_023_213, w_018_271);
  not1 I023_216(w_023_216, w_018_227);
  nand2 I023_219(w_023_219, w_000_907, w_008_420);
  and2 I023_227(w_023_227, w_010_060, w_013_090);
  nand2 I023_232(w_023_232, w_010_188, w_015_258);
  and2 I023_235(w_023_235, w_020_107, w_020_210);
  nand2 I023_236(w_023_236, w_020_317, w_012_403);
  not1 I023_237(w_023_237, w_015_181);
  nand2 I023_238(w_023_238, w_010_282, w_012_529);
  or2  I023_243(w_023_243, w_016_012, w_010_221);
  nand2 I023_245(w_023_245, w_016_016, w_017_1422);
  nand2 I023_250(w_023_250, w_018_235, w_007_757);
  and2 I023_253(w_023_253, w_021_261, w_007_228);
  nand2 I023_255(w_023_255, w_008_266, w_006_118);
  and2 I023_256(w_023_256, w_002_359, w_011_309);
  or2  I023_257(w_023_257, w_018_019, w_006_246);
  nand2 I023_261(w_023_261, w_000_1161, w_022_181);
  nand2 I023_262(w_023_262, w_008_394, w_004_1773);
  and2 I023_265(w_023_265, w_021_260, w_018_262);
  not1 I023_266(w_023_266, w_015_049);
  nand2 I023_269(w_023_269, w_011_159, w_021_274);
  nand2 I023_277(w_023_277, w_002_223, w_009_050);
  or2  I023_278(w_023_278, w_008_608, w_021_093);
  nand2 I023_280(w_023_280, w_002_487, w_016_017);
  not1 I023_282(w_023_282, w_008_074);
  nand2 I023_283(w_023_283, w_002_198, w_011_067);
  or2  I023_289(w_023_289, w_005_1617, w_013_143);
  or2  I023_290(w_023_290, w_010_186, w_009_059);
  nand2 I023_291(w_023_291, w_000_537, w_009_024);
  nand2 I023_293(w_023_293, w_021_134, w_015_118);
  nand2 I023_294(w_023_294, w_005_1168, w_018_010);
  or2  I023_299(w_023_299, w_000_057, w_002_478);
  and2 I023_300(w_023_300, w_005_052, w_003_287);
  and2 I023_301(w_023_301, w_001_1115, w_018_011);
  nand2 I023_311(w_023_311, w_019_859, w_008_679);
  not1 I023_318(w_023_318, w_000_725);
  not1 I023_319(w_023_319, w_011_444);
  or2  I023_321(w_023_321, w_007_270, w_016_000);
  or2  I023_328(w_023_328, w_000_982, w_012_281);
  not1 I023_329(w_023_329, w_007_453);
  or2  I023_331(w_023_331, w_013_047, w_007_881);
  and2 I023_333(w_023_333, w_001_141, w_021_081);
  nand2 I023_334(w_023_334, w_000_1784, w_005_593);
  and2 I023_335(w_023_335, w_012_095, w_020_525);
  or2  I023_336(w_023_336, w_013_190, w_009_062);
  or2  I023_338(w_023_338, w_013_049, w_002_578);
  nand2 I023_339(w_023_339, w_021_033, w_016_015);
  not1 I023_342(w_023_342, w_009_101);
  and2 I023_345(w_023_345, w_008_438, w_001_569);
  and2 I023_347(w_023_347, w_005_272, w_012_401);
  nand2 I023_348(w_023_348, w_003_031, w_003_172);
  not1 I023_349(w_023_349, w_006_081);
  or2  I023_353(w_023_353, w_011_197, w_017_1284);
  and2 I023_355(w_023_355, w_005_1355, w_009_020);
  nand2 I023_357(w_023_357, w_020_039, w_021_082);
  nand2 I023_359(w_023_359, w_003_171, w_001_1606);
  or2  I023_364(w_023_364, w_012_436, w_021_261);
  or2  I023_367(w_023_367, w_002_229, w_019_411);
  not1 I023_379(w_023_379, w_007_360);
  not1 I023_380(w_023_380, w_007_439);
  or2  I023_412(w_023_412, w_006_162, w_016_032);
  or2  I023_414(w_023_414, w_009_092, w_011_086);
  or2  I023_447(w_023_447, w_022_113, w_003_279);
  or2  I023_448(w_023_448, w_007_137, w_003_026);
  or2  I023_449(w_023_449, w_015_124, w_018_003);
  or2  I023_450(w_023_450, w_007_048, w_016_009);
  and2 I023_459(w_023_459, w_002_054, w_012_594);
  and2 I023_474(w_023_474, w_022_305, w_001_1499);
  and2 I023_476(w_023_476, w_019_815, w_017_624);
  or2  I023_479(w_023_479, w_003_225, w_002_381);
  not1 I023_487(w_023_487, w_000_143);
  or2  I023_491(w_023_491, w_019_598, w_013_251);
  or2  I023_496(w_023_496, w_007_229, w_010_217);
  or2  I023_498(w_023_498, w_021_242, w_004_1851);
  or2  I023_502(w_023_502, w_016_004, w_002_099);
  and2 I023_514(w_023_514, w_017_508, w_013_141);
  and2 I023_515(w_023_515, w_006_250, w_019_647);
  or2  I023_527(w_023_527, w_014_059, w_011_803);
  nand2 I023_533(w_023_533, w_019_692, w_005_791);
  not1 I023_538(w_023_538, w_003_053);
  and2 I023_546(w_023_546, w_017_1639, w_021_180);
  nand2 I023_553(w_023_553, w_018_228, w_006_031);
  or2  I023_558(w_023_558, w_014_168, w_019_451);
  not1 I023_577(w_023_577, w_004_249);
  or2  I023_585(w_023_585, w_003_055, w_019_718);
  nand2 I023_589(w_023_589, w_002_569, w_020_867);
  and2 I023_596(w_023_596, w_004_418, w_003_275);
  or2  I023_614(w_023_614, w_002_211, w_021_006);
  or2  I023_622(w_023_622, w_019_726, w_002_564);
  and2 I023_624(w_023_624, w_013_235, w_010_106);
  and2 I023_625(w_023_625, w_010_299, w_005_962);
  or2  I023_632(w_023_632, w_006_224, w_016_005);
  or2  I023_635(w_023_635, w_009_099, w_001_837);
  or2  I023_640(w_023_640, w_019_219, w_016_018);
  and2 I023_642(w_023_642, w_011_548, w_019_377);
  not1 I023_646(w_023_646, w_022_152);
  nand2 I023_648(w_023_648, w_018_007, w_014_534);
  nand2 I023_650(w_023_650, w_018_115, w_002_138);
  or2  I023_654(w_023_654, w_000_416, w_001_677);
  or2  I023_656(w_023_656, w_016_017, w_011_643);
  not1 I023_666(w_023_666, w_017_1163);
  and2 I023_667(w_023_667, w_007_605, w_013_062);
  and2 I023_679(w_023_679, w_014_717, w_020_348);
  and2 I023_682(w_023_682, w_012_235, w_010_210);
  or2  I023_702(w_023_702, w_007_214, w_002_534);
  nand2 I023_708(w_023_708, w_000_073, w_015_093);
  or2  I023_710(w_023_710, w_018_121, w_006_071);
  and2 I023_718(w_023_718, w_008_027, w_014_500);
  not1 I023_720(w_023_720, w_001_023);
  not1 I023_726(w_023_726, w_011_152);
  not1 I023_732(w_023_732, w_017_1182);
  or2  I023_733(w_023_733, w_011_127, w_000_1046);
  or2  I023_736(w_023_736, w_020_517, w_008_712);
  nand2 I023_748(w_023_748, w_021_136, w_014_703);
  or2  I023_758(w_023_758, w_002_574, w_003_272);
  not1 I023_759(w_023_759, w_010_246);
  not1 I023_764(w_023_764, w_008_081);
  nand2 I023_769(w_023_769, w_017_218, w_006_033);
  and2 I023_775(w_023_775, w_022_146, w_007_1555);
  not1 I023_776(w_023_776, w_002_234);
  or2  I023_780(w_023_780, w_003_233, w_012_627);
  and2 I023_785(w_023_785, w_005_564, w_011_739);
  nand2 I023_787(w_023_787, w_022_194, w_013_225);
  and2 I023_791(w_023_791, w_011_584, w_018_218);
  or2  I023_811(w_023_811, w_017_303, w_002_297);
  and2 I023_818(w_023_818, w_021_223, w_006_225);
  or2  I023_820(w_023_820, w_022_076, w_006_308);
  nand2 I023_822(w_023_822, w_020_265, w_003_107);
  and2 I023_824(w_023_824, w_011_815, w_016_000);
  or2  I023_826(w_023_826, w_018_144, w_009_098);
  and2 I023_829(w_023_829, w_011_491, w_001_813);
  and2 I023_834(w_023_834, w_002_174, w_008_721);
  or2  I023_836(w_023_836, w_003_161, w_001_010);
  or2  I023_848(w_023_848, w_016_013, w_017_1598);
  not1 I023_849(w_023_849, w_018_024);
  not1 I023_852(w_023_852, w_000_495);
  not1 I023_864(w_023_864, w_004_059);
  not1 I023_878(w_023_878, w_020_520);
  or2  I023_880(w_023_880, w_003_001, w_022_335);
  or2  I023_882(w_023_882, w_003_170, w_018_254);
  not1 I023_885(w_023_885, w_015_273);
  nand2 I023_902(w_023_902, w_019_001, w_011_839);
  and2 I023_903(w_023_903, w_017_1606, w_022_109);
  not1 I023_906(w_023_906, w_014_020);
  and2 I023_914(w_023_914, w_009_036, w_006_039);
  nand2 I023_915(w_023_915, w_021_128, w_005_279);
  not1 I023_921(w_023_921, w_009_055);
  not1 I023_929(w_023_929, w_001_1177);
  nand2 I023_934(w_023_934, w_002_477, w_012_514);
  not1 I023_937(w_023_937, w_017_450);
  nand2 I023_939(w_023_939, w_000_1912, w_005_168);
  not1 I023_956(w_023_956, w_013_097);
  or2  I023_969(w_023_969, w_008_078, w_013_168);
  and2 I023_974(w_023_974, w_021_136, w_012_268);
  nand2 I023_986(w_023_986, w_014_017, w_015_185);
  or2  I023_994(w_023_994, w_001_1423, w_022_178);
  nand2 I023_996(w_023_996, w_017_1655, w_020_929);
  not1 I023_1004(w_023_1004, w_015_073);
  not1 I023_1006(w_023_1006, w_018_131);
  or2  I023_1007(w_023_1007, w_009_006, w_015_049);
  and2 I023_1013(w_023_1013, w_018_168, w_012_097);
  or2  I023_1019(w_023_1019, w_004_592, w_021_137);
  or2  I023_1023(w_023_1023, w_020_1235, w_005_154);
  or2  I023_1026(w_023_1026, w_004_000, w_008_263);
  not1 I023_1031(w_023_1031, w_001_1413);
  nand2 I023_1037(w_023_1037, w_008_488, w_001_1077);
  not1 I023_1043(w_023_1043, w_022_016);
  nand2 I023_1046(w_023_1046, w_004_901, w_005_1668);
  not1 I023_1065(w_023_1065, w_010_037);
  not1 I023_1068(w_023_1068, w_006_109);
  or2  I023_1090(w_023_1090, w_010_067, w_001_659);
  nand2 I023_1098(w_023_1098, w_002_145, w_015_058);
  or2  I023_1105(w_023_1105, w_005_077, w_018_254);
  and2 I023_1114(w_023_1114, w_012_021, w_019_278);
  or2  I023_1115(w_023_1115, w_017_1079, w_018_104);
  or2  I023_1116(w_023_1116, w_012_193, w_022_120);
  not1 I023_1132(w_023_1132, w_011_042);
  or2  I023_1140(w_023_1140, w_016_020, w_004_1637);
  or2  I023_1141(w_023_1141, w_011_435, w_002_120);
  nand2 I023_1153(w_023_1153, w_017_777, w_001_815);
  not1 I023_1156(w_023_1156, w_015_274);
  nand2 I023_1163(w_023_1163, w_002_082, w_000_451);
  not1 I023_1166(w_023_1166, w_003_028);
  nand2 I023_1168(w_023_1168, w_012_143, w_011_572);
  and2 I023_1179(w_023_1179, w_001_820, w_011_137);
  nand2 I023_1180(w_023_1180, w_015_204, w_005_322);
  nand2 I023_1182(w_023_1182, w_012_351, w_017_998);
  not1 I023_1194(w_023_1194, w_021_050);
  nand2 I023_1196(w_023_1196, w_012_513, w_017_218);
  not1 I023_1199(w_023_1199, w_003_123);
  or2  I023_1200(w_023_1200, w_012_574, w_000_313);
  or2  I023_1208(w_023_1208, w_018_110, w_007_1397);
  or2  I023_1216(w_023_1216, w_001_313, w_004_1449);
  not1 I023_1218(w_023_1218, w_004_182);
  and2 I023_1219(w_023_1219, w_019_230, w_001_128);
  or2  I023_1225(w_023_1225, w_007_1487, w_006_061);
  not1 I023_1226(w_023_1226, w_001_232);
  or2  I023_1259(w_023_1259, w_013_332, w_017_1232);
  or2  I023_1262(w_023_1262, w_016_017, w_005_722);
  and2 I023_1265(w_023_1265, w_021_272, w_008_632);
  and2 I023_1266(w_023_1266, w_020_217, w_013_170);
  nand2 I023_1273(w_023_1273, w_015_135, w_005_199);
  nand2 I023_1275(w_023_1275, w_011_073, w_020_162);
  nand2 I023_1283(w_023_1283, w_019_643, w_018_269);
  or2  I023_1284(w_023_1284, w_021_180, w_006_186);
  nand2 I023_1292(w_023_1292, w_005_620, w_016_019);
  not1 I023_1294(w_023_1294, w_003_163);
  and2 I023_1298(w_023_1298, w_009_111, w_022_262);
  nand2 I023_1313(w_023_1313, w_022_064, w_015_094);
  not1 I023_1318(w_023_1318, w_005_886);
  nand2 I023_1327(w_023_1327, w_005_015, w_008_312);
  not1 I023_1336(w_023_1336, w_001_166);
  and2 I023_1348(w_023_1348, w_002_115, w_008_243);
  not1 I023_1357(w_023_1357, w_014_451);
  or2  I023_1363(w_023_1363, w_022_267, w_022_399);
  nand2 I023_1364(w_023_1364, w_017_428, w_007_391);
  or2  I023_1369(w_023_1369, w_020_946, w_009_104);
  or2  I023_1371(w_023_1371, w_019_183, w_006_298);
  and2 I023_1380(w_023_1380, w_015_031, w_022_096);
  not1 I023_1391(w_023_1391, w_016_015);
  nand2 I023_1396(w_023_1396, w_021_021, w_020_453);
  not1 I023_1398(w_023_1398, w_013_325);
  not1 I023_1410(w_023_1410, w_013_205);
  or2  I023_1412(w_023_1412, w_011_001, w_018_072);
  not1 I023_1421(w_023_1421, w_020_671);
  and2 I023_1431(w_023_1431, w_005_035, w_022_297);
  nand2 I023_1439(w_023_1439, w_004_1283, w_008_751);
  not1 I023_1452(w_023_1452, w_010_054);
  nand2 I023_1455(w_023_1455, w_021_019, w_009_058);
  or2  I023_1460(w_023_1460, w_017_393, w_011_622);
  and2 I023_1474(w_023_1474, w_020_869, w_022_185);
  and2 I023_1484(w_023_1484, w_003_013, w_007_351);
  and2 I023_1494(w_023_1494, w_021_187, w_008_163);
  not1 I023_1502(w_023_1502, w_019_287);
  or2  I023_1503(w_023_1503, w_003_264, w_004_1893);
  and2 I023_1507(w_023_1507, w_021_081, w_004_1016);
  not1 I023_1543(w_023_1543, w_009_081);
  or2  I023_1544(w_023_1544, w_002_481, w_022_377);
  or2  I023_1545(w_023_1545, w_015_133, w_010_226);
  and2 I023_1553(w_023_1553, w_013_177, w_013_031);
  not1 I023_1560(w_023_1560, w_006_279);
  not1 I023_1567(w_023_1567, w_017_921);
  nand2 I023_1569(w_023_1569, w_008_500, w_017_1778);
  nand2 I023_1572(w_023_1572, w_019_577, w_002_342);
  nand2 I023_1573(w_023_1573, w_006_105, w_020_1063);
  nand2 I023_1580(w_023_1580, w_003_195, w_015_039);
  and2 I023_1585(w_023_1585, w_010_306, w_018_190);
  nand2 I023_1594(w_023_1594, w_016_004, w_013_041);
  and2 I023_1595(w_023_1595, w_014_606, w_000_293);
  not1 I023_1596(w_023_1596, w_017_124);
  not1 I023_1598(w_023_1598, w_009_023);
  or2  I023_1604(w_023_1604, w_007_999, w_011_120);
  or2  I023_1607(w_023_1607, w_011_640, w_009_082);
  and2 I023_1608(w_023_1608, w_001_1299, w_009_084);
  nand2 I023_1612(w_023_1612, w_008_376, w_000_1154);
  or2  I024_000(w_024_000, w_020_517, w_007_084);
  and2 I024_002(w_024_002, w_009_012, w_000_279);
  or2  I024_003(w_024_003, w_002_458, w_009_039);
  and2 I024_004(w_024_004, w_001_793, w_008_294);
  not1 I024_009(w_024_009, w_004_1625);
  nand2 I024_011(w_024_011, w_005_179, w_008_605);
  nand2 I024_016(w_024_016, w_009_048, w_002_593);
  not1 I024_017(w_024_017, w_000_716);
  or2  I024_018(w_024_018, w_021_088, w_021_005);
  or2  I024_022(w_024_022, w_020_440, w_020_1085);
  or2  I024_028(w_024_028, w_003_317, w_014_191);
  and2 I024_029(w_024_029, w_010_099, w_019_025);
  and2 I024_031(w_024_031, w_000_1943, w_019_707);
  or2  I024_032(w_024_032, w_003_288, w_007_059);
  not1 I024_035(w_024_035, w_008_566);
  nand2 I024_038(w_024_038, w_017_478, w_004_364);
  nand2 I024_043(w_024_043, w_023_577, w_004_1025);
  nand2 I024_044(w_024_044, w_001_796, w_018_140);
  and2 I024_047(w_024_047, w_004_1616, w_022_132);
  not1 I024_054(w_024_054, w_000_1460);
  not1 I024_055(w_024_055, w_012_410);
  or2  I024_059(w_024_059, w_005_318, w_014_688);
  nand2 I024_061(w_024_061, w_014_277, w_003_298);
  nand2 I024_062(w_024_062, w_015_198, w_023_1046);
  not1 I024_064(w_024_064, w_007_987);
  and2 I024_065(w_024_065, w_016_005, w_001_1349);
  nand2 I024_066(w_024_066, w_007_869, w_007_215);
  nand2 I024_071(w_024_071, w_004_1216, w_008_157);
  nand2 I024_072(w_024_072, w_012_078, w_015_091);
  not1 I024_075(w_024_075, w_003_306);
  nand2 I024_077(w_024_077, w_023_1369, w_002_165);
  and2 I024_081(w_024_081, w_007_124, w_002_165);
  or2  I024_082(w_024_082, w_017_873, w_016_032);
  and2 I024_084(w_024_084, w_004_225, w_002_480);
  or2  I024_087(w_024_087, w_020_007, w_021_268);
  or2  I024_088(w_024_088, w_018_221, w_002_076);
  nand2 I024_089(w_024_089, w_019_365, w_020_597);
  nand2 I024_091(w_024_091, w_015_238, w_007_532);
  not1 I024_092(w_024_092, w_012_569);
  and2 I024_095(w_024_095, w_016_008, w_002_154);
  and2 I024_098(w_024_098, w_019_152, w_003_200);
  not1 I024_103(w_024_103, w_019_1059);
  not1 I024_107(w_024_107, w_012_188);
  nand2 I024_111(w_024_111, w_001_1412, w_003_207);
  not1 I024_114(w_024_114, w_014_545);
  not1 I024_120(w_024_120, w_020_032);
  and2 I024_121(w_024_121, w_003_044, w_017_1710);
  nand2 I024_125(w_024_125, w_012_164, w_009_088);
  not1 I024_126(w_024_126, w_023_070);
  and2 I024_127(w_024_127, w_005_236, w_020_1176);
  or2  I024_132(w_024_132, w_008_374, w_009_024);
  not1 I024_134(w_024_134, w_011_115);
  or2  I024_143(w_024_143, w_019_595, w_001_1656);
  nand2 I024_145(w_024_145, w_015_251, w_003_236);
  nand2 I024_146(w_024_146, w_001_702, w_020_350);
  and2 I024_148(w_024_148, w_003_106, w_010_302);
  or2  I024_153(w_024_153, w_007_1189, w_023_1284);
  and2 I024_163(w_024_163, w_017_1457, w_008_521);
  and2 I024_164(w_024_164, w_004_935, w_004_1123);
  nand2 I024_165(w_024_165, w_012_295, w_023_448);
  not1 I024_166(w_024_166, w_021_085);
  or2  I024_168(w_024_168, w_003_003, w_019_1022);
  or2  I024_173(w_024_173, w_000_400, w_007_057);
  not1 I024_177(w_024_177, w_007_039);
  not1 I024_178(w_024_178, w_008_314);
  nand2 I024_179(w_024_179, w_020_510, w_001_895);
  and2 I024_182(w_024_182, w_007_187, w_021_064);
  not1 I024_186(w_024_186, w_009_081);
  or2  I024_189(w_024_189, w_019_842, w_014_506);
  and2 I024_194(w_024_194, w_021_035, w_009_001);
  and2 I024_195(w_024_195, w_021_134, w_001_031);
  or2  I024_197(w_024_197, w_013_321, w_010_139);
  nand2 I024_199(w_024_199, w_007_1522, w_006_215);
  and2 I024_200(w_024_200, w_002_211, w_012_091);
  not1 I024_201(w_024_201, w_021_000);
  not1 I024_208(w_024_208, w_010_109);
  and2 I024_211(w_024_211, w_023_632, w_019_643);
  not1 I024_212(w_024_212, w_023_311);
  not1 I024_217(w_024_217, w_001_661);
  nand2 I024_218(w_024_218, w_009_035, w_020_138);
  not1 I024_220(w_024_220, w_003_212);
  and2 I024_221(w_024_221, w_010_041, w_001_231);
  or2  I024_222(w_024_222, w_022_002, w_020_559);
  or2  I024_243(w_024_243, w_019_220, w_018_244);
  not1 I024_245(w_024_245, w_007_1248);
  nand2 I024_247(w_024_247, w_012_237, w_008_165);
  not1 I024_250(w_024_250, w_019_756);
  and2 I024_252(w_024_252, w_014_147, w_016_005);
  not1 I024_260(w_024_260, w_004_788);
  nand2 I024_262(w_024_262, w_023_181, w_000_1579);
  or2  I024_263(w_024_263, w_006_251, w_006_276);
  and2 I024_265(w_024_265, w_006_187, w_001_1121);
  and2 I024_269(w_024_269, w_009_049, w_007_176);
  nand2 I024_274(w_024_274, w_002_522, w_008_412);
  nand2 I024_277(w_024_277, w_022_385, w_003_115);
  not1 I024_282(w_024_282, w_007_272);
  or2  I024_284(w_024_284, w_010_177, w_012_157);
  nand2 I024_285(w_024_285, w_004_417, w_006_150);
  not1 I024_288(w_024_288, w_018_263);
  or2  I024_289(w_024_289, w_003_229, w_017_1059);
  nand2 I024_290(w_024_290, w_002_141, w_012_276);
  nand2 I024_292(w_024_292, w_011_547, w_011_791);
  nand2 I024_293(w_024_293, w_015_093, w_002_311);
  or2  I024_297(w_024_297, w_003_106, w_022_116);
  and2 I024_299(w_024_299, w_019_596, w_011_794);
  or2  I024_301(w_024_301, w_006_208, w_023_849);
  or2  I024_303(w_024_303, w_017_300, w_007_580);
  not1 I024_304(w_024_304, w_021_214);
  or2  I024_308(w_024_308, w_002_240, w_012_628);
  and2 I024_309(w_024_309, w_014_138, w_013_295);
  not1 I024_310(w_024_310, w_012_559);
  and2 I024_311(w_024_311, w_010_275, w_015_222);
  and2 I024_313(w_024_313, w_017_1607, w_014_375);
  or2  I024_316(w_024_316, w_000_1090, w_023_245);
  or2  I024_318(w_024_318, w_019_113, w_014_005);
  or2  I024_323(w_024_323, w_021_027, w_004_922);
  and2 I024_335(w_024_335, w_011_157, w_006_035);
  or2  I024_336(w_024_336, w_000_391, w_013_297);
  and2 I024_337(w_024_337, w_018_030, w_005_1593);
  and2 I024_342(w_024_342, w_019_978, w_009_059);
  not1 I024_345(w_024_345, w_008_554);
  not1 I024_346(w_024_346, w_011_694);
  or2  I024_347(w_024_347, w_014_556, w_019_778);
  and2 I024_348(w_024_348, w_014_365, w_020_1021);
  or2  I024_349(w_024_349, w_015_235, w_011_263);
  or2  I024_351(w_024_351, w_010_239, w_000_083);
  and2 I024_355(w_024_355, w_000_388, w_018_152);
  and2 I024_366(w_024_366, w_020_448, w_006_155);
  and2 I024_380(w_024_380, w_009_005, w_022_204);
  or2  I024_403(w_024_403, w_003_013, w_020_252);
  nand2 I024_415(w_024_415, w_014_326, w_022_105);
  or2  I024_425(w_024_425, w_018_223, w_009_012);
  and2 I024_430(w_024_430, w_021_214, w_006_234);
  and2 I024_435(w_024_435, w_014_745, w_002_194);
  not1 I024_439(w_024_439, w_005_1609);
  and2 I024_444(w_024_444, w_010_115, w_016_034);
  nand2 I024_453(w_024_453, w_012_547, w_010_328);
  or2  I024_460(w_024_460, w_020_611, w_023_093);
  and2 I024_462(w_024_462, w_020_045, w_020_096);
  and2 I024_468(w_024_468, w_021_122, w_016_014);
  not1 I024_471(w_024_471, w_007_763);
  not1 I024_473(w_024_473, w_018_197);
  and2 I024_480(w_024_480, w_005_1243, w_005_503);
  and2 I024_488(w_024_488, w_006_097, w_010_337);
  nand2 I024_503(w_024_503, w_009_095, w_015_187);
  nand2 I024_506(w_024_506, w_020_111, w_023_253);
  not1 I024_509(w_024_509, w_010_225);
  and2 I024_514(w_024_514, w_015_280, w_014_477);
  nand2 I024_524(w_024_524, w_018_136, w_017_1550);
  and2 I024_528(w_024_528, w_010_023, w_014_125);
  nand2 I024_533(w_024_533, w_008_564, w_012_407);
  nand2 I024_539(w_024_539, w_002_220, w_014_074);
  and2 I024_542(w_024_542, w_015_268, w_012_487);
  and2 I024_559(w_024_559, w_018_144, w_000_1772);
  or2  I024_563(w_024_563, w_022_416, w_004_1637);
  and2 I024_577(w_024_577, w_015_275, w_013_210);
  nand2 I024_585(w_024_585, w_014_319, w_017_102);
  or2  I024_593(w_024_593, w_022_267, w_014_158);
  and2 I024_596(w_024_596, w_018_078, w_001_1622);
  not1 I024_606(w_024_606, w_001_1687);
  nand2 I024_610(w_024_610, w_007_924, w_015_034);
  nand2 I024_616(w_024_616, w_001_569, w_010_086);
  or2  I024_617(w_024_617, w_018_135, w_022_007);
  not1 I024_621(w_024_621, w_008_132);
  or2  I024_647(w_024_647, w_017_1541, w_018_012);
  not1 I024_677(w_024_677, w_021_002);
  not1 I024_679(w_024_679, w_010_394);
  or2  I024_682(w_024_682, w_000_847, w_016_029);
  or2  I024_683(w_024_683, w_014_345, w_022_036);
  not1 I024_685(w_024_685, w_012_374);
  or2  I024_686(w_024_686, w_014_124, w_005_115);
  or2  I024_688(w_024_688, w_022_079, w_010_012);
  not1 I024_692(w_024_692, w_017_1935);
  or2  I024_700(w_024_700, w_003_152, w_014_070);
  and2 I024_723(w_024_723, w_012_277, w_009_045);
  or2  I024_735(w_024_735, w_005_1136, w_009_019);
  nand2 I024_736(w_024_736, w_018_006, w_011_244);
  nand2 I024_741(w_024_741, w_021_092, w_016_014);
  not1 I024_757(w_024_757, w_016_007);
  and2 I024_761(w_024_761, w_008_209, w_008_562);
  or2  I024_772(w_024_772, w_001_262, w_023_020);
  not1 I024_777(w_024_777, w_001_199);
  nand2 I024_778(w_024_778, w_006_074, w_015_011);
  or2  I024_781(w_024_781, w_013_014, w_010_038);
  nand2 I024_785(w_024_785, w_021_276, w_006_150);
  nand2 I024_790(w_024_790, w_021_023, w_000_907);
  not1 I024_791(w_024_791, w_007_1161);
  and2 I024_800(w_024_800, w_006_014, w_015_041);
  or2  I024_812(w_024_812, w_023_1168, w_002_494);
  or2  I024_823(w_024_823, w_016_012, w_012_404);
  not1 I024_827(w_024_827, w_011_104);
  nand2 I024_830(w_024_830, w_019_876, w_023_1543);
  and2 I024_840(w_024_840, w_017_1694, w_022_018);
  or2  I024_842(w_024_842, w_016_015, w_008_728);
  and2 I024_844(w_024_844, w_017_077, w_018_236);
  nand2 I024_857(w_024_857, w_013_103, w_009_027);
  not1 I024_869(w_024_869, w_000_1557);
  and2 I024_874(w_024_874, w_011_041, w_016_029);
  not1 I024_880(w_024_880, w_004_364);
  not1 I024_882(w_024_882, w_003_157);
  not1 I024_887(w_024_887, w_010_129);
  not1 I024_888(w_024_888, w_009_106);
  or2  I024_895(w_024_895, w_015_133, w_004_218);
  or2  I024_899(w_024_899, w_020_154, w_013_309);
  and2 I024_905(w_024_905, w_023_1006, w_022_148);
  and2 I024_915(w_024_915, w_023_769, w_023_934);
  not1 I024_917(w_024_917, w_011_244);
  or2  I024_918(w_024_918, w_000_010, w_006_035);
  not1 I024_924(w_024_924, w_015_131);
  nand2 I024_927(w_024_927, w_005_733, w_004_588);
  nand2 I024_929(w_024_929, w_022_287, w_021_128);
  and2 I024_933(w_024_933, w_017_985, w_004_558);
  not1 I024_934(w_024_934, w_008_633);
  or2  I024_939(w_024_939, w_014_078, w_005_143);
  nand2 I024_940(w_024_940, w_009_030, w_005_1561);
  or2  I024_944(w_024_944, w_005_1149, w_004_1189);
  nand2 I024_949(w_024_949, w_015_144, w_007_850);
  or2  I024_964(w_024_964, w_006_085, w_006_243);
  nand2 I024_965(w_024_965, w_012_268, w_012_328);
  and2 I024_972(w_024_972, w_002_247, w_012_546);
  not1 I024_976(w_024_976, w_018_125);
  nand2 I024_977(w_024_977, w_000_906, w_016_027);
  nand2 I024_986(w_024_986, w_021_080, w_010_284);
  not1 I024_995(w_024_995, w_021_259);
  and2 I024_998(w_024_998, w_005_1310, w_016_006);
  not1 I024_1001(w_024_1001, w_006_048);
  nand2 I024_1003(w_024_1003, w_019_782, w_002_401);
  not1 I024_1006(w_024_1006, w_017_1422);
  nand2 I024_1009(w_024_1009, w_016_001, w_017_846);
  nand2 I024_1010(w_024_1010, w_012_292, w_017_534);
  and2 I024_1032(w_024_1032, w_001_1319, w_015_131);
  nand2 I024_1050(w_024_1050, w_011_773, w_018_268);
  not1 I024_1053(w_024_1053, w_020_887);
  or2  I024_1055(w_024_1055, w_014_144, w_020_227);
  and2 I024_1059(w_024_1059, w_002_177, w_002_096);
  nand2 I024_1066(w_024_1066, w_018_194, w_010_040);
  nand2 I024_1076(w_024_1076, w_023_1364, w_020_1020);
  or2  I024_1079(w_024_1079, w_007_1459, w_011_406);
  nand2 I024_1085(w_024_1085, w_009_092, w_020_312);
  and2 I024_1089(w_024_1089, w_019_537, w_007_1157);
  and2 I024_1094(w_024_1094, w_004_809, w_000_1414);
  and2 I024_1098(w_024_1098, w_023_650, w_005_643);
  nand2 I024_1105(w_024_1105, w_012_660, w_010_124);
  not1 I024_1121(w_024_1121, w_011_042);
  nand2 I024_1133(w_024_1133, w_007_124, w_013_160);
  and2 I024_1137(w_024_1137, w_005_1187, w_010_375);
  not1 I024_1164(w_024_1164, w_013_275);
  or2  I024_1187(w_024_1187, w_011_147, w_001_345);
  not1 I024_1188(w_024_1188, w_003_014);
  nand2 I024_1190(w_024_1190, w_010_275, w_014_189);
  and2 I024_1193(w_024_1193, w_016_004, w_017_1924);
  and2 I024_1203(w_024_1203, w_002_002, w_012_050);
  and2 I024_1221(w_024_1221, w_022_152, w_013_144);
  nand2 I024_1225(w_024_1225, w_005_132, w_004_842);
  or2  I024_1226(w_024_1226, w_010_215, w_007_236);
  not1 I024_1230(w_024_1230, w_016_035);
  and2 I024_1235(w_024_1235, w_000_626, w_017_539);
  nand2 I024_1241(w_024_1241, w_016_034, w_011_360);
  or2  I024_1244(w_024_1244, w_018_211, w_019_463);
  nand2 I024_1248(w_024_1248, w_022_013, w_006_114);
  and2 I024_1250(w_024_1250, w_002_081, w_009_045);
  or2  I024_1261(w_024_1261, w_019_101, w_009_057);
  nand2 I024_1269(w_024_1269, w_010_033, w_021_135);
  or2  I024_1276(w_024_1276, w_003_093, w_012_452);
  or2  I024_1297(w_024_1297, w_015_137, w_022_343);
  and2 I024_1320(w_024_1320, w_021_136, w_002_359);
  nand2 I024_1327(w_024_1327, w_023_1585, w_000_1946);
  and2 I024_1341(w_024_1341, w_002_590, w_007_306);
  or2  I024_1362(w_024_1362, w_017_1792, w_009_072);
  and2 I024_1377(w_024_1377, w_004_056, w_012_261);
  or2  I024_1383(w_024_1383, w_011_698, w_001_031);
  not1 I024_1385(w_024_1385, w_018_038);
  nand2 I024_1393(w_024_1393, w_000_218, w_013_025);
  nand2 I024_1399(w_024_1399, w_000_626, w_023_311);
  nand2 I024_1401(w_024_1401, w_016_030, w_012_461);
  and2 I024_1404(w_024_1404, w_023_142, w_003_226);
  not1 I024_1408(w_024_1408, w_000_950);
  nand2 I024_1422(w_024_1422, w_003_003, w_014_218);
  not1 I024_1424(w_024_1424, w_017_468);
  not1 I024_1430(w_024_1430, w_000_225);
  and2 I024_1431(w_024_1431, w_017_694, w_001_1193);
  not1 I024_1438(w_024_1438, w_013_019);
  or2  I024_1465(w_024_1465, w_000_1306, w_015_036);
  and2 I024_1466(w_024_1466, w_004_1406, w_023_1391);
  or2  I024_1473(w_024_1473, w_005_1180, w_014_598);
  and2 I024_1478(w_024_1478, w_013_263, w_005_1173);
  not1 I024_1489(w_024_1489, w_019_702);
  nand2 I024_1495(w_024_1495, w_000_249, w_012_222);
  and2 I024_1498(w_024_1498, w_000_1342, w_011_185);
  or2  I024_1504(w_024_1504, w_017_1636, w_006_148);
  and2 I024_1522(w_024_1522, w_019_058, w_009_102);
  not1 I024_1523(w_024_1523, w_022_031);
  or2  I024_1539(w_024_1539, w_022_129, w_018_187);
  not1 I024_1544(w_024_1544, w_023_003);
  or2  I024_1545(w_024_1545, w_010_203, w_006_265);
  nand2 I024_1555(w_024_1555, w_000_1376, w_002_213);
  not1 I024_1557(w_024_1557, w_001_1067);
  and2 I024_1561(w_024_1561, w_010_414, w_012_319);
  not1 I024_1563(w_024_1563, w_010_002);
  or2  I024_1568(w_024_1568, w_014_508, w_001_885);
  nand2 I024_1569(w_024_1569, w_006_237, w_013_171);
  nand2 I024_1570(w_024_1570, w_023_1545, w_023_020);
  or2  I024_1572(w_024_1572, w_012_040, w_004_398);
  or2  I024_1576(w_024_1576, w_000_1356, w_010_315);
  nand2 I024_1579(w_024_1579, w_018_139, w_019_305);
  not1 I024_1583(w_024_1583, w_019_881);
  and2 I024_1590(w_024_1590, w_011_060, w_017_525);
  nand2 I024_1591(w_024_1591, w_023_091, w_000_629);
  nand2 I024_1607(w_024_1607, w_017_253, w_008_016);
  nand2 I024_1615(w_024_1615, w_002_558, w_006_293);
  nand2 I024_1617(w_024_1617, w_017_459, w_004_1236);
  nand2 I024_1622(w_024_1622, w_007_451, w_005_1652);
  or2  I024_1623(w_024_1623, w_002_463, w_016_034);
  and2 I024_1624(w_024_1624, w_012_476, w_008_125);
  not1 I024_1638(w_024_1638, w_013_179);
  or2  I024_1640(w_024_1640, w_005_208, w_013_055);
  nand2 I024_1642(w_024_1642, w_021_136, w_016_037);
  or2  I024_1645(w_024_1645, w_021_201, w_011_199);
  or2  I024_1649(w_024_1649, w_022_153, w_006_288);
  nand2 I025_000(w_025_000, w_017_133, w_015_274);
  or2  I025_006(w_025_006, w_019_593, w_012_018);
  not1 I025_007(w_025_007, w_007_1536);
  nand2 I025_008(w_025_008, w_007_329, w_019_691);
  nand2 I025_013(w_025_013, w_006_108, w_015_130);
  not1 I025_014(w_025_014, w_024_1430);
  or2  I025_015(w_025_015, w_006_111, w_009_000);
  nand2 I025_016(w_025_016, w_014_581, w_019_353);
  not1 I025_017(w_025_017, w_002_263);
  and2 I025_021(w_025_021, w_021_050, w_011_753);
  and2 I025_022(w_025_022, w_017_1216, w_008_577);
  nand2 I025_029(w_025_029, w_003_183, w_006_009);
  or2  I025_031(w_025_031, w_016_029, w_024_1495);
  or2  I025_032(w_025_032, w_001_242, w_007_597);
  and2 I025_034(w_025_034, w_017_087, w_018_155);
  nand2 I025_035(w_025_035, w_024_091, w_010_198);
  and2 I025_036(w_025_036, w_023_885, w_020_622);
  and2 I025_059(w_025_059, w_009_037, w_010_328);
  and2 I025_061(w_025_061, w_010_242, w_012_625);
  or2  I025_064(w_025_064, w_001_1323, w_010_346);
  not1 I025_070(w_025_070, w_002_394);
  or2  I025_080(w_025_080, w_024_077, w_002_150);
  and2 I025_081(w_025_081, w_022_103, w_012_338);
  nand2 I025_082(w_025_082, w_007_406, w_010_420);
  and2 I025_088(w_025_088, w_008_675, w_009_096);
  and2 I025_092(w_025_092, w_011_734, w_017_183);
  not1 I025_097(w_025_097, w_010_094);
  not1 I025_099(w_025_099, w_019_465);
  and2 I025_100(w_025_100, w_003_041, w_020_160);
  and2 I025_101(w_025_101, w_007_127, w_007_280);
  and2 I025_102(w_025_102, w_017_1140, w_006_204);
  or2  I025_106(w_025_106, w_001_200, w_001_621);
  nand2 I025_111(w_025_111, w_005_943, w_007_221);
  or2  I025_116(w_025_116, w_017_1633, w_017_044);
  not1 I025_119(w_025_119, w_016_030);
  nand2 I025_137(w_025_137, w_020_842, w_002_121);
  or2  I025_142(w_025_142, w_015_087, w_018_228);
  not1 I025_145(w_025_145, w_003_315);
  not1 I025_150(w_025_150, w_020_895);
  and2 I025_165(w_025_165, w_013_156, w_019_610);
  and2 I025_171(w_025_171, w_022_196, w_015_012);
  and2 I025_172(w_025_172, w_003_044, w_000_1591);
  nand2 I025_173(w_025_173, w_022_113, w_019_099);
  or2  I025_177(w_025_177, w_022_335, w_014_412);
  and2 I025_178(w_025_178, w_006_340, w_006_255);
  or2  I025_179(w_025_179, w_009_094, w_002_568);
  not1 I025_180(w_025_180, w_023_237);
  not1 I025_182(w_025_182, w_014_824);
  not1 I025_186(w_025_186, w_005_677);
  or2  I025_198(w_025_198, w_000_1947, w_015_016);
  or2  I025_202(w_025_202, w_022_046, w_009_067);
  nand2 I025_206(w_025_206, w_009_000, w_004_303);
  or2  I025_208(w_025_208, w_009_065, w_007_1276);
  not1 I025_209(w_025_209, w_006_055);
  nand2 I025_216(w_025_216, w_021_265, w_021_051);
  and2 I025_221(w_025_221, w_018_068, w_002_374);
  and2 I025_230(w_025_230, w_001_614, w_024_347);
  or2  I025_232(w_025_232, w_006_267, w_012_051);
  and2 I025_235(w_025_235, w_008_821, w_006_124);
  and2 I025_240(w_025_240, w_000_413, w_023_412);
  or2  I025_243(w_025_243, w_007_1442, w_016_012);
  and2 I025_244(w_025_244, w_004_1834, w_003_128);
  nand2 I025_247(w_025_247, w_000_1194, w_015_025);
  and2 I025_253(w_025_253, w_000_1240, w_011_063);
  not1 I025_255(w_025_255, w_008_152);
  or2  I025_259(w_025_259, w_014_604, w_008_750);
  or2  I025_262(w_025_262, w_008_574, w_008_787);
  or2  I025_267(w_025_267, w_001_790, w_023_589);
  or2  I025_287(w_025_287, w_018_187, w_020_870);
  and2 I025_289(w_025_289, w_016_032, w_006_305);
  or2  I025_290(w_025_290, w_022_428, w_014_384);
  and2 I025_298(w_025_298, w_015_214, w_015_210);
  and2 I025_300(w_025_300, w_020_603, w_024_514);
  not1 I025_307(w_025_307, w_011_159);
  nand2 I025_311(w_025_311, w_018_196, w_022_029);
  and2 I025_314(w_025_314, w_020_373, w_015_116);
  or2  I025_327(w_025_327, w_009_063, w_005_529);
  and2 I025_328(w_025_328, w_024_1523, w_008_014);
  nand2 I025_335(w_025_335, w_017_1224, w_022_225);
  or2  I025_337(w_025_337, w_013_257, w_003_040);
  not1 I025_342(w_025_342, w_007_1119);
  and2 I025_352(w_025_352, w_015_065, w_017_1416);
  and2 I025_355(w_025_355, w_001_712, w_003_203);
  and2 I025_358(w_025_358, w_002_331, w_016_031);
  nand2 I025_374(w_025_374, w_021_182, w_006_105);
  nand2 I025_377(w_025_377, w_010_064, w_020_892);
  nand2 I025_389(w_025_389, w_011_152, w_019_188);
  and2 I025_390(w_025_390, w_012_519, w_022_051);
  nand2 I025_396(w_025_396, w_005_255, w_012_559);
  not1 I025_414(w_025_414, w_013_108);
  or2  I025_416(w_025_416, w_019_844, w_004_1679);
  not1 I025_420(w_025_420, w_019_1007);
  and2 I025_422(w_025_422, w_022_185, w_014_529);
  nand2 I025_434(w_025_434, w_008_574, w_018_205);
  or2  I025_435(w_025_435, w_007_964, w_022_234);
  or2  I025_437(w_025_437, w_016_008, w_023_1474);
  nand2 I025_451(w_025_451, w_013_118, w_024_1422);
  or2  I025_455(w_025_455, w_004_1374, w_018_189);
  not1 I025_456(w_025_456, w_006_002);
  nand2 I025_458(w_025_458, w_022_027, w_023_1507);
  or2  I025_479(w_025_479, w_002_475, w_012_172);
  or2  I025_481(w_025_481, w_010_083, w_005_239);
  nand2 I025_491(w_025_491, w_016_027, w_017_990);
  not1 I025_492(w_025_492, w_020_521);
  or2  I025_502(w_025_502, w_004_1811, w_021_155);
  not1 I025_515(w_025_515, w_009_000);
  or2  I025_518(w_025_518, w_017_007, w_002_578);
  nand2 I025_521(w_025_521, w_015_052, w_018_127);
  or2  I025_527(w_025_527, w_024_1399, w_021_185);
  not1 I025_547(w_025_547, w_017_322);
  not1 I025_548(w_025_548, w_009_019);
  or2  I025_552(w_025_552, w_013_099, w_022_349);
  nand2 I025_553(w_025_553, w_011_692, w_000_590);
  not1 I025_556(w_025_556, w_021_048);
  nand2 I025_565(w_025_565, w_006_058, w_001_674);
  and2 I025_570(w_025_570, w_003_093, w_009_060);
  nand2 I025_573(w_025_573, w_010_184, w_013_033);
  and2 I025_579(w_025_579, w_008_413, w_024_995);
  nand2 I025_580(w_025_580, w_012_045, w_001_291);
  not1 I025_592(w_025_592, w_024_004);
  or2  I025_593(w_025_593, w_005_385, w_021_002);
  nand2 I025_596(w_025_596, w_002_022, w_007_244);
  not1 I025_601(w_025_601, w_000_162);
  not1 I025_604(w_025_604, w_022_322);
  nand2 I025_617(w_025_617, w_012_603, w_005_163);
  not1 I025_629(w_025_629, w_005_1057);
  or2  I025_630(w_025_630, w_011_368, w_004_1780);
  or2  I025_639(w_025_639, w_018_235, w_017_143);
  not1 I025_647(w_025_647, w_020_1139);
  nand2 I025_649(w_025_649, w_020_359, w_009_029);
  not1 I025_657(w_025_657, w_009_022);
  nand2 I025_661(w_025_661, w_006_264, w_003_013);
  or2  I025_668(w_025_668, w_002_579, w_006_009);
  and2 I025_679(w_025_679, w_013_122, w_024_1085);
  or2  I025_683(w_025_683, w_016_013, w_024_1341);
  and2 I025_688(w_025_688, w_010_059, w_020_487);
  not1 I025_695(w_025_695, w_004_1265);
  nand2 I025_697(w_025_697, w_001_1000, w_006_091);
  and2 I025_699(w_025_699, w_002_280, w_020_649);
  not1 I025_704(w_025_704, w_020_1163);
  not1 I025_705(w_025_705, w_010_408);
  not1 I025_707(w_025_707, w_013_323);
  not1 I025_711(w_025_711, w_022_321);
  and2 I025_712(w_025_712, w_016_017, w_022_061);
  and2 I025_718(w_025_718, w_003_104, w_007_298);
  and2 I025_719(w_025_719, w_005_1213, w_009_091);
  nand2 I025_725(w_025_725, w_024_1489, w_019_310);
  not1 I025_730(w_025_730, w_024_348);
  nand2 I025_734(w_025_734, w_009_044, w_022_392);
  nand2 I025_738(w_025_738, w_001_745, w_007_1065);
  or2  I025_739(w_025_739, w_000_1095, w_023_009);
  and2 I025_747(w_025_747, w_011_850, w_004_540);
  nand2 I025_759(w_025_759, w_003_203, w_017_1694);
  not1 I025_766(w_025_766, w_009_049);
  or2  I025_768(w_025_768, w_002_555, w_005_1027);
  and2 I025_775(w_025_775, w_020_875, w_020_116);
  nand2 I025_777(w_025_777, w_001_733, w_015_176);
  or2  I025_779(w_025_779, w_018_035, w_007_520);
  and2 I025_780(w_025_780, w_012_514, w_008_041);
  not1 I025_782(w_025_782, w_013_326);
  or2  I025_783(w_025_783, w_007_1250, w_024_533);
  and2 I025_788(w_025_788, w_021_073, w_006_009);
  and2 I025_795(w_025_795, w_009_051, w_018_249);
  nand2 I025_810(w_025_810, w_001_1563, w_011_196);
  or2  I025_815(w_025_815, w_007_1527, w_005_1059);
  nand2 I025_817(w_025_817, w_017_1133, w_007_623);
  or2  I025_823(w_025_823, w_013_170, w_003_025);
  or2  I025_824(w_025_824, w_020_441, w_013_003);
  not1 I025_825(w_025_825, w_021_210);
  nand2 I025_837(w_025_837, w_015_039, w_016_010);
  and2 I025_839(w_025_839, w_008_104, w_019_521);
  not1 I025_842(w_025_842, w_001_029);
  not1 I025_848(w_025_848, w_017_1552);
  and2 I025_877(w_025_877, w_004_1401, w_007_851);
  and2 I025_888(w_025_888, w_018_193, w_013_123);
  and2 I025_897(w_025_897, w_021_258, w_004_979);
  nand2 I025_911(w_025_911, w_009_065, w_012_447);
  or2  I025_913(w_025_913, w_010_303, w_018_184);
  or2  I025_914(w_025_914, w_001_1227, w_000_459);
  or2  I025_938(w_025_938, w_011_315, w_005_082);
  not1 I025_941(w_025_941, w_019_133);
  and2 I025_953(w_025_953, w_013_316, w_014_738);
  nand2 I025_959(w_025_959, w_009_008, w_022_060);
  not1 I025_961(w_025_961, w_009_017);
  not1 I025_976(w_025_976, w_024_366);
  or2  I025_982(w_025_982, w_023_1396, w_022_430);
  or2  I025_983(w_025_983, w_001_148, w_008_053);
  not1 I025_988(w_025_988, w_003_136);
  and2 I025_992(w_025_992, w_012_265, w_000_322);
  and2 I025_999(w_025_999, w_011_233, w_019_1084);
  and2 I025_1002(w_025_1002, w_017_1670, w_022_058);
  or2  I025_1004(w_025_1004, w_011_856, w_000_1347);
  nand2 I025_1006(w_025_1006, w_018_196, w_014_023);
  or2  I025_1007(w_025_1007, w_008_484, w_010_397);
  not1 I025_1025(w_025_1025, w_022_311);
  or2  I025_1028(w_025_1028, w_002_255, w_004_029);
  and2 I025_1036(w_025_1036, w_011_390, w_009_061);
  or2  I025_1037(w_025_1037, w_000_275, w_006_323);
  nand2 I025_1041(w_025_1041, w_005_206, w_018_157);
  nand2 I025_1042(w_025_1042, w_021_167, w_001_1260);
  or2  I025_1047(w_025_1047, w_014_729, w_006_189);
  nand2 I025_1048(w_025_1048, w_001_1661, w_004_598);
  not1 I025_1051(w_025_1051, w_010_217);
  not1 I025_1053(w_025_1053, w_002_135);
  or2  I025_1065(w_025_1065, w_013_304, w_011_227);
  not1 I025_1070(w_025_1070, w_011_785);
  not1 I025_1079(w_025_1079, w_010_188);
  and2 I025_1083(w_025_1083, w_014_161, w_021_130);
  not1 I025_1084(w_025_1084, w_018_124);
  and2 I025_1085(w_025_1085, w_009_031, w_020_696);
  and2 I025_1094(w_025_1094, w_005_240, w_017_373);
  not1 I025_1097(w_025_1097, w_017_396);
  nand2 I025_1120(w_025_1120, w_002_196, w_013_086);
  or2  I025_1124(w_025_1124, w_009_047, w_003_202);
  or2  I025_1125(w_025_1125, w_021_116, w_002_271);
  not1 I025_1126(w_025_1126, w_003_139);
  and2 I025_1134(w_025_1134, w_011_363, w_015_194);
  nand2 I025_1161(w_025_1161, w_002_587, w_000_1213);
  nand2 I025_1164(w_025_1164, w_011_230, w_009_095);
  or2  I025_1169(w_025_1169, w_007_660, w_015_101);
  or2  I025_1170(w_025_1170, w_000_1932, w_023_1585);
  and2 I025_1174(w_025_1174, w_018_108, w_009_098);
  not1 I025_1192(w_025_1192, w_022_043);
  nand2 I025_1211(w_025_1211, w_019_297, w_019_110);
  or2  I025_1222(w_025_1222, w_024_145, w_012_617);
  or2  I025_1241(w_025_1241, w_003_305, w_000_017);
  or2  I025_1242(w_025_1242, w_017_1672, w_016_027);
  or2  I025_1243(w_025_1243, w_002_123, w_015_103);
  or2  I025_1249(w_025_1249, w_019_775, w_012_659);
  or2  I025_1251(w_025_1251, w_007_288, w_008_534);
  and2 I025_1258(w_025_1258, w_005_124, w_019_682);
  or2  I025_1265(w_025_1265, w_005_025, w_003_239);
  nand2 I025_1273(w_025_1273, w_024_1076, w_021_034);
  or2  I025_1280(w_025_1280, w_001_720, w_019_402);
  and2 I025_1287(w_025_1287, w_011_460, w_005_655);
  nand2 I025_1295(w_025_1295, w_006_287, w_009_103);
  nand2 I025_1304(w_025_1304, w_011_037, w_019_527);
  nand2 I025_1309(w_025_1309, w_020_487, w_001_039);
  not1 I025_1317(w_025_1317, w_000_1223);
  nand2 I025_1321(w_025_1321, w_010_294, w_017_1913);
  nand2 I025_1338(w_025_1338, w_012_176, w_007_252);
  and2 I025_1341(w_025_1341, w_023_1598, w_013_036);
  and2 I025_1350(w_025_1350, w_004_537, w_003_044);
  nand2 I025_1351(w_025_1351, w_000_1717, w_012_161);
  not1 I025_1357(w_025_1357, w_010_128);
  nand2 I025_1374(w_025_1374, w_018_280, w_023_848);
  and2 I025_1375(w_025_1375, w_012_619, w_013_274);
  or2  I025_1379(w_025_1379, w_012_293, w_016_037);
  nand2 I025_1391(w_025_1391, w_004_588, w_006_008);
  or2  I025_1399(w_025_1399, w_005_223, w_022_386);
  nand2 I025_1401(w_025_1401, w_000_641, w_011_072);
  not1 I025_1406(w_025_1406, w_023_614);
  or2  I025_1407(w_025_1407, w_024_002, w_017_681);
  not1 I025_1408(w_025_1408, w_017_1322);
  or2  I025_1412(w_025_1412, w_007_210, w_003_038);
  or2  I025_1425(w_025_1425, w_024_103, w_019_257);
  or2  I025_1426(w_025_1426, w_011_469, w_024_1003);
  nand2 I025_1432(w_025_1432, w_007_380, w_021_225);
  nand2 I025_1433(w_025_1433, w_007_1209, w_020_677);
  nand2 I025_1434(w_025_1434, w_007_1103, w_023_558);
  not1 I025_1441(w_025_1441, w_016_018);
  not1 I025_1442(w_025_1442, w_021_254);
  nand2 I025_1452(w_025_1452, w_008_372, w_005_694);
  and2 I025_1456(w_025_1456, w_023_199, w_018_209);
  and2 I025_1469(w_025_1469, w_022_038, w_015_005);
  or2  I025_1472(w_025_1472, w_010_005, w_020_687);
  or2  I025_1476(w_025_1476, w_004_527, w_015_083);
  and2 I025_1483(w_025_1483, w_017_623, w_011_813);
  nand2 I025_1484(w_025_1484, w_010_169, w_001_103);
  or2  I025_1495(w_025_1495, w_021_211, w_011_119);
  and2 I025_1498(w_025_1498, w_022_310, w_010_012);
  not1 I025_1508(w_025_1508, w_023_347);
  and2 I025_1520(w_025_1520, w_011_425, w_009_050);
  nand2 I025_1524(w_025_1524, w_015_082, w_021_205);
  nand2 I025_1529(w_025_1529, w_013_288, w_011_543);
  or2  I025_1533(w_025_1533, w_006_224, w_014_263);
  nand2 I025_1537(w_025_1537, w_012_289, w_014_049);
  or2  I025_1538(w_025_1538, w_014_578, w_011_449);
  and2 I025_1540(w_025_1540, w_012_487, w_023_243);
  nand2 I025_1543(w_025_1543, w_003_011, w_012_076);
  and2 I025_1544(w_025_1544, w_018_028, w_023_262);
  or2  I025_1549(w_025_1549, w_012_006, w_007_449);
  not1 I025_1550(w_025_1550, w_020_720);
  nand2 I025_1564(w_025_1564, w_014_246, w_017_1206);
  not1 I025_1572(w_025_1572, w_001_562);
  or2  I025_1575(w_025_1575, w_000_1294, w_015_216);
  or2  I025_1597(w_025_1597, w_021_092, w_021_099);
  not1 I025_1611(w_025_1611, w_021_153);
  nand2 I025_1615(w_025_1615, w_014_159, w_001_1627);
  not1 I025_1622(w_025_1622, w_000_830);
  or2  I025_1626(w_025_1626, w_007_277, w_021_207);
  nand2 I025_1629(w_025_1629, w_004_003, w_019_106);
  nand2 I025_1633(w_025_1633, w_008_201, w_016_008);
  or2  I025_1651(w_025_1651, w_013_291, w_012_104);
  or2  I025_1655(w_025_1655, w_014_268, w_014_640);
  or2  I025_1661(w_025_1661, w_015_066, w_019_328);
  nand2 I025_1668(w_025_1668, w_007_1574, w_012_027);
  not1 I025_1671(w_025_1671, w_018_004);
  or2  I025_1674(w_025_1674, w_009_022, w_024_791);
  or2  I025_1675(w_025_1675, w_012_507, w_001_062);
  or2  I025_1678(w_025_1678, w_016_015, w_013_140);
  and2 I025_1698(w_025_1698, w_014_453, w_001_1172);
  not1 I025_1703(w_025_1703, w_014_092);
  or2  I026_001(w_026_001, w_020_239, w_025_1295);
  and2 I026_005(w_026_005, w_018_272, w_011_391);
  nand2 I026_007(w_026_007, w_023_213, w_015_154);
  or2  I026_010(w_026_010, w_025_244, w_004_248);
  or2  I026_011(w_026_011, w_020_332, w_007_378);
  nand2 I026_020(w_026_020, w_020_651, w_024_199);
  not1 I026_022(w_026_022, w_012_493);
  and2 I026_024(w_026_024, w_019_689, w_015_146);
  and2 I026_027(w_026_027, w_015_067, w_014_014);
  or2  I026_045(w_026_045, w_019_090, w_024_292);
  nand2 I026_048(w_026_048, w_005_488, w_021_257);
  nand2 I026_055(w_026_055, w_014_234, w_022_148);
  or2  I026_056(w_026_056, w_020_376, w_011_598);
  nand2 I026_058(w_026_058, w_009_016, w_017_1531);
  and2 I026_060(w_026_060, w_010_203, w_025_414);
  not1 I026_065(w_026_065, w_001_644);
  and2 I026_068(w_026_068, w_011_332, w_022_370);
  not1 I026_069(w_026_069, w_022_365);
  and2 I026_073(w_026_073, w_012_609, w_002_051);
  or2  I026_074(w_026_074, w_008_644, w_011_749);
  and2 I026_075(w_026_075, w_015_291, w_022_168);
  or2  I026_079(w_026_079, w_019_673, w_011_648);
  nand2 I026_090(w_026_090, w_017_472, w_022_037);
  nand2 I026_097(w_026_097, w_025_1434, w_013_228);
  or2  I026_099(w_026_099, w_015_194, w_025_422);
  and2 I026_103(w_026_103, w_010_133, w_012_571);
  and2 I026_106(w_026_106, w_005_333, w_012_486);
  not1 I026_108(w_026_108, w_018_078);
  and2 I026_110(w_026_110, w_025_661, w_014_540);
  and2 I026_117(w_026_117, w_011_536, w_023_342);
  nand2 I026_119(w_026_119, w_017_813, w_024_075);
  nand2 I026_123(w_026_123, w_011_209, w_014_270);
  not1 I026_125(w_026_125, w_002_411);
  or2  I026_127(w_026_127, w_009_035, w_012_258);
  and2 I026_134(w_026_134, w_023_321, w_013_184);
  nand2 I026_136(w_026_136, w_015_281, w_024_1248);
  or2  I026_144(w_026_144, w_021_151, w_015_201);
  and2 I026_148(w_026_148, w_024_430, w_020_674);
  or2  I026_152(w_026_152, w_025_604, w_011_081);
  not1 I026_153(w_026_153, w_019_1008);
  and2 I026_154(w_026_154, w_005_1522, w_019_633);
  and2 I026_155(w_026_155, w_013_254, w_005_021);
  nand2 I026_156(w_026_156, w_008_651, w_023_787);
  and2 I026_159(w_026_159, w_004_730, w_015_007);
  and2 I026_161(w_026_161, w_003_156, w_019_897);
  and2 I026_170(w_026_170, w_020_720, w_005_630);
  nand2 I026_172(w_026_172, w_022_295, w_000_1536);
  nand2 I026_175(w_026_175, w_003_169, w_016_020);
  not1 I026_189(w_026_189, w_023_1216);
  not1 I026_190(w_026_190, w_017_1301);
  nand2 I026_192(w_026_192, w_000_059, w_014_623);
  or2  I026_195(w_026_195, w_000_1193, w_012_224);
  nand2 I026_201(w_026_201, w_006_174, w_014_664);
  not1 I026_203(w_026_203, w_007_028);
  or2  I026_216(w_026_216, w_002_566, w_007_1042);
  nand2 I026_218(w_026_218, w_020_327, w_019_132);
  or2  I026_219(w_026_219, w_002_424, w_022_275);
  and2 I026_224(w_026_224, w_004_1344, w_022_026);
  not1 I026_227(w_026_227, w_017_045);
  nand2 I026_230(w_026_230, w_018_203, w_008_025);
  not1 I026_233(w_026_233, w_023_824);
  and2 I026_234(w_026_234, w_014_342, w_003_273);
  not1 I026_236(w_026_236, w_017_075);
  not1 I026_238(w_026_238, w_009_001);
  and2 I026_257(w_026_257, w_012_130, w_024_777);
  nand2 I026_258(w_026_258, w_020_1062, w_006_311);
  nand2 I026_262(w_026_262, w_012_478, w_003_109);
  not1 I026_265(w_026_265, w_008_253);
  nand2 I026_266(w_026_266, w_004_1053, w_025_1498);
  or2  I026_267(w_026_267, w_025_657, w_004_1502);
  not1 I026_268(w_026_268, w_003_296);
  nand2 I026_275(w_026_275, w_022_153, w_003_091);
  or2  I026_276(w_026_276, w_022_058, w_003_127);
  or2  I026_287(w_026_287, w_007_015, w_019_500);
  or2  I026_288(w_026_288, w_013_226, w_018_066);
  and2 I026_291(w_026_291, w_001_926, w_005_1147);
  nand2 I026_295(w_026_295, w_020_359, w_019_216);
  or2  I026_300(w_026_300, w_023_335, w_003_151);
  and2 I026_311(w_026_311, w_001_117, w_013_289);
  and2 I026_317(w_026_317, w_007_027, w_002_328);
  and2 I026_318(w_026_318, w_015_047, w_011_092);
  not1 I026_324(w_026_324, w_011_440);
  not1 I026_325(w_026_325, w_021_055);
  not1 I026_330(w_026_330, w_003_058);
  not1 I026_331(w_026_331, w_013_222);
  not1 I026_337(w_026_337, w_024_221);
  nand2 I026_341(w_026_341, w_022_128, w_003_281);
  or2  I026_345(w_026_345, w_006_180, w_006_218);
  and2 I026_352(w_026_352, w_013_236, w_021_096);
  nand2 I026_354(w_026_354, w_018_254, w_002_248);
  nand2 I026_360(w_026_360, w_016_015, w_004_909);
  not1 I026_366(w_026_366, w_012_445);
  and2 I026_374(w_026_374, w_017_1126, w_003_122);
  and2 I026_376(w_026_376, w_022_417, w_013_029);
  and2 I026_378(w_026_378, w_005_143, w_012_201);
  nand2 I026_379(w_026_379, w_008_297, w_012_470);
  nand2 I026_382(w_026_382, w_007_1003, w_009_049);
  and2 I026_388(w_026_388, w_017_457, w_002_163);
  nand2 I026_394(w_026_394, w_017_1818, w_005_752);
  or2  I026_396(w_026_396, w_021_149, w_025_502);
  nand2 I026_404(w_026_404, w_015_042, w_000_292);
  not1 I026_416(w_026_416, w_022_045);
  nand2 I026_419(w_026_419, w_007_946, w_016_018);
  and2 I026_423(w_026_423, w_005_046, w_025_451);
  or2  I026_431(w_026_431, w_017_106, w_012_292);
  not1 I026_435(w_026_435, w_010_114);
  not1 I026_439(w_026_439, w_014_123);
  not1 I026_440(w_026_440, w_018_225);
  nand2 I026_443(w_026_443, w_004_188, w_005_1620);
  not1 I026_446(w_026_446, w_014_518);
  nand2 I026_449(w_026_449, w_021_161, w_006_246);
  or2  I026_450(w_026_450, w_011_022, w_020_203);
  nand2 I026_451(w_026_451, w_004_1288, w_005_812);
  not1 I026_453(w_026_453, w_012_090);
  and2 I026_457(w_026_457, w_018_266, w_002_180);
  nand2 I026_466(w_026_466, w_006_078, w_015_162);
  nand2 I026_467(w_026_467, w_018_092, w_007_1343);
  or2  I026_468(w_026_468, w_018_253, w_010_037);
  not1 I026_480(w_026_480, w_005_377);
  and2 I026_481(w_026_481, w_008_211, w_009_024);
  and2 I026_491(w_026_491, w_013_119, w_001_362);
  nand2 I026_510(w_026_510, w_005_212, w_014_567);
  nand2 I026_515(w_026_515, w_003_173, w_005_228);
  and2 I026_521(w_026_521, w_011_762, w_012_400);
  nand2 I026_533(w_026_533, w_015_225, w_004_1329);
  not1 I026_545(w_026_545, w_008_758);
  or2  I026_567(w_026_567, w_015_189, w_023_154);
  and2 I026_570(w_026_570, w_018_263, w_001_512);
  nand2 I026_572(w_026_572, w_011_193, w_023_479);
  not1 I026_577(w_026_577, w_009_044);
  not1 I026_588(w_026_588, w_003_045);
  nand2 I026_595(w_026_595, w_012_232, w_019_401);
  or2  I026_597(w_026_597, w_003_224, w_009_059);
  or2  I026_601(w_026_601, w_005_485, w_014_453);
  and2 I026_602(w_026_602, w_007_1256, w_004_197);
  and2 I026_609(w_026_609, w_012_559, w_024_933);
  not1 I026_610(w_026_610, w_011_128);
  not1 I026_620(w_026_620, w_025_1661);
  and2 I026_622(w_026_622, w_003_309, w_011_009);
  or2  I026_639(w_026_639, w_004_449, w_022_300);
  and2 I026_650(w_026_650, w_011_444, w_012_026);
  nand2 I026_654(w_026_654, w_000_324, w_017_040);
  and2 I026_658(w_026_658, w_007_654, w_024_103);
  or2  I026_660(w_026_660, w_014_649, w_011_339);
  or2  I026_661(w_026_661, w_001_1044, w_022_402);
  nand2 I026_665(w_026_665, w_015_247, w_014_545);
  nand2 I026_666(w_026_666, w_023_380, w_008_096);
  and2 I026_671(w_026_671, w_009_043, w_001_806);
  nand2 I026_691(w_026_691, w_024_323, w_005_1337);
  and2 I026_695(w_026_695, w_003_096, w_004_322);
  nand2 I026_699(w_026_699, w_011_327, w_025_1484);
  or2  I026_717(w_026_717, w_008_663, w_019_419);
  or2  I026_723(w_026_723, w_007_1511, w_008_646);
  and2 I026_725(w_026_725, w_022_309, w_008_464);
  or2  I026_741(w_026_741, w_002_300, w_006_139);
  nand2 I026_750(w_026_750, w_015_150, w_020_941);
  not1 I026_751(w_026_751, w_018_134);
  nand2 I026_763(w_026_763, w_003_087, w_019_668);
  not1 I026_771(w_026_771, w_021_084);
  nand2 I026_772(w_026_772, w_012_409, w_016_018);
  and2 I026_777(w_026_777, w_017_1578, w_001_192);
  not1 I026_785(w_026_785, w_013_161);
  or2  I026_790(w_026_790, w_014_528, w_001_1467);
  or2  I026_797(w_026_797, w_005_1271, w_001_233);
  not1 I026_813(w_026_813, w_006_239);
  not1 I026_815(w_026_815, w_005_971);
  or2  I026_817(w_026_817, w_021_177, w_014_204);
  nand2 I026_820(w_026_820, w_009_083, w_014_607);
  and2 I026_830(w_026_830, w_017_007, w_024_682);
  not1 I026_838(w_026_838, w_009_029);
  and2 I026_843(w_026_843, w_015_205, w_009_044);
  nand2 I026_844(w_026_844, w_003_232, w_008_224);
  or2  I026_846(w_026_846, w_006_090, w_012_579);
  and2 I026_860(w_026_860, w_023_147, w_000_259);
  not1 I026_871(w_026_871, w_000_606);
  nand2 I026_874(w_026_874, w_014_654, w_013_148);
  or2  I026_879(w_026_879, w_025_013, w_013_169);
  or2  I026_882(w_026_882, w_004_314, w_000_902);
  or2  I026_884(w_026_884, w_003_259, w_013_131);
  nand2 I026_901(w_026_901, w_018_273, w_020_629);
  nand2 I026_905(w_026_905, w_009_009, w_003_302);
  not1 I026_909(w_026_909, w_021_045);
  nand2 I026_937(w_026_937, w_007_1443, w_016_036);
  nand2 I026_949(w_026_949, w_011_866, w_019_753);
  or2  I026_952(w_026_952, w_019_151, w_005_910);
  nand2 I026_955(w_026_955, w_021_255, w_019_205);
  not1 I026_984(w_026_984, w_006_131);
  and2 I026_987(w_026_987, w_002_163, w_017_029);
  or2  I026_991(w_026_991, w_021_241, w_005_386);
  and2 I026_993(w_026_993, w_025_1703, w_008_652);
  or2  I026_994(w_026_994, w_009_017, w_003_070);
  not1 I026_995(w_026_995, w_008_805);
  and2 I026_997(w_026_997, w_010_403, w_006_086);
  nand2 I026_998(w_026_998, w_021_009, w_017_1036);
  not1 I026_1002(w_026_1002, w_009_033);
  or2  I026_1006(w_026_1006, w_006_264, w_019_881);
  or2  I026_1008(w_026_1008, w_015_240, w_011_650);
  or2  I026_1012(w_026_1012, w_005_116, w_024_1607);
  or2  I026_1016(w_026_1016, w_022_374, w_009_058);
  not1 I026_1026(w_026_1026, w_016_017);
  or2  I026_1027(w_026_1027, w_002_212, w_018_190);
  and2 I026_1028(w_026_1028, w_000_1328, w_010_281);
  not1 I026_1029(w_026_1029, w_001_188);
  not1 I026_1031(w_026_1031, w_022_412);
  not1 I026_1035(w_026_1035, w_000_1625);
  not1 I026_1043(w_026_1043, w_013_004);
  nand2 I026_1044(w_026_1044, w_022_399, w_006_224);
  not1 I026_1048(w_026_1048, w_014_830);
  and2 I026_1070(w_026_1070, w_007_439, w_015_131);
  not1 I026_1071(w_026_1071, w_018_192);
  or2  I026_1072(w_026_1072, w_007_072, w_016_034);
  and2 I026_1080(w_026_1080, w_005_1603, w_025_953);
  and2 I026_1084(w_026_1084, w_011_527, w_023_283);
  or2  I026_1094(w_026_1094, w_021_013, w_005_029);
  not1 I026_1097(w_026_1097, w_007_1333);
  nand2 I026_1105(w_026_1105, w_025_1622, w_025_775);
  not1 I026_1107(w_026_1107, w_022_353);
  and2 I026_1109(w_026_1109, w_022_153, w_020_538);
  or2  I026_1111(w_026_1111, w_010_017, w_012_107);
  not1 I026_1112(w_026_1112, w_012_214);
  not1 I026_1113(w_026_1113, w_018_090);
  and2 I026_1116(w_026_1116, w_001_471, w_007_1555);
  not1 I026_1123(w_026_1123, w_020_476);
  or2  I026_1126(w_026_1126, w_007_1465, w_014_807);
  or2  I026_1135(w_026_1135, w_017_1828, w_009_099);
  and2 I026_1136(w_026_1136, w_015_120, w_023_1132);
  and2 I026_1155(w_026_1155, w_000_1806, w_025_1483);
  and2 I026_1158(w_026_1158, w_005_1478, w_016_010);
  and2 I026_1159(w_026_1159, w_022_376, w_016_006);
  nand2 I026_1169(w_026_1169, w_008_114, w_008_534);
  or2  I026_1177(w_026_1177, w_025_1065, w_023_1560);
  or2  I026_1178(w_026_1178, w_015_137, w_007_304);
  and2 I026_1182(w_026_1182, w_012_558, w_007_802);
  not1 I026_1186(w_026_1186, w_012_353);
  not1 I026_1201(w_026_1201, w_008_524);
  and2 I026_1202(w_026_1202, w_003_010, w_003_016);
  or2  I026_1221(w_026_1221, w_018_198, w_004_359);
  nand2 I026_1223(w_026_1223, w_016_009, w_009_018);
  or2  I026_1226(w_026_1226, w_006_193, w_015_070);
  and2 I026_1240(w_026_1240, w_008_310, w_021_028);
  nand2 I026_1243(w_026_1243, w_006_033, w_012_428);
  not1 I026_1244(w_026_1244, w_011_169);
  and2 I026_1253(w_026_1253, w_015_068, w_014_551);
  not1 I026_1257(w_026_1257, w_025_182);
  not1 I026_1260(w_026_1260, w_018_046);
  not1 I026_1268(w_026_1268, w_013_111);
  not1 I026_1274(w_026_1274, w_005_154);
  or2  I026_1277(w_026_1277, w_014_819, w_024_335);
  nand2 I026_1287(w_026_1287, w_019_524, w_014_398);
  nand2 I026_1289(w_026_1289, w_025_1097, w_015_073);
  not1 I026_1296(w_026_1296, w_000_998);
  nand2 I026_1297(w_026_1297, w_009_002, w_002_431);
  and2 I026_1304(w_026_1304, w_022_141, w_003_239);
  nand2 I026_1305(w_026_1305, w_011_314, w_020_315);
  or2  I026_1316(w_026_1316, w_025_116, w_023_720);
  nand2 I026_1325(w_026_1325, w_018_267, w_006_278);
  nand2 I026_1336(w_026_1336, w_007_111, w_006_278);
  or2  I026_1347(w_026_1347, w_017_675, w_013_124);
  nand2 I026_1356(w_026_1356, w_004_1875, w_011_584);
  nand2 I026_1357(w_026_1357, w_019_604, w_012_588);
  or2  I026_1359(w_026_1359, w_011_262, w_010_190);
  or2  I026_1365(w_026_1365, w_003_272, w_023_974);
  nand2 I026_1366(w_026_1366, w_009_092, w_000_1618);
  and2 I026_1371(w_026_1371, w_014_360, w_014_709);
  or2  I026_1376(w_026_1376, w_006_199, w_012_228);
  nand2 I026_1407(w_026_1407, w_022_302, w_004_445);
  nand2 I026_1415(w_026_1415, w_001_1671, w_000_1679);
  and2 I026_1418(w_026_1418, w_020_383, w_010_168);
  not1 I026_1424(w_026_1424, w_010_173);
  or2  I026_1427(w_026_1427, w_020_1189, w_000_1949);
  not1 I026_1429(w_026_1429, w_023_1369);
  not1 I026_1436(w_026_1436, w_012_022);
  nand2 I026_1443(w_026_1443, w_017_812, w_017_779);
  nand2 I026_1448(w_026_1448, w_018_160, w_001_379);
  or2  I026_1455(w_026_1455, w_015_069, w_021_048);
  not1 I026_1456(w_026_1456, w_000_466);
  or2  I026_1463(w_026_1463, w_025_1524, w_012_421);
  not1 I026_1467(w_026_1467, w_018_162);
  not1 I026_1470(w_026_1470, w_017_984);
  or2  I026_1483(w_026_1483, w_004_886, w_010_311);
  and2 I026_1489(w_026_1489, w_010_329, w_002_293);
  not1 I026_1491(w_026_1491, w_013_038);
  or2  I026_1507(w_026_1507, w_025_390, w_023_1200);
  not1 I026_1512(w_026_1512, w_025_186);
  nand2 I026_1520(w_026_1520, w_020_1043, w_022_231);
  and2 I027_001(w_027_001, w_012_040, w_005_1596);
  and2 I027_003(w_027_003, w_022_075, w_021_224);
  not1 I027_006(w_027_006, w_007_945);
  and2 I027_007(w_027_007, w_017_197, w_016_037);
  or2  I027_008(w_027_008, w_011_583, w_025_1433);
  or2  I027_011(w_027_011, w_025_647, w_019_476);
  nand2 I027_012(w_027_012, w_015_079, w_016_030);
  and2 I027_013(w_027_013, w_021_053, w_016_000);
  not1 I027_014(w_027_014, w_024_972);
  nand2 I027_016(w_027_016, w_007_524, w_023_1023);
  or2  I027_017(w_027_017, w_023_338, w_003_200);
  nand2 I027_018(w_027_018, w_022_298, w_015_119);
  and2 I027_019(w_027_019, w_020_498, w_012_428);
  not1 I027_028(w_027_028, w_021_000);
  nand2 I027_029(w_027_029, w_009_058, w_003_019);
  and2 I027_032(w_027_032, w_017_1020, w_024_346);
  not1 I027_033(w_027_033, w_006_334);
  nand2 I027_038(w_027_038, w_007_1562, w_020_663);
  and2 I027_040(w_027_040, w_012_288, w_015_043);
  not1 I027_041(w_027_041, w_022_280);
  not1 I027_043(w_027_043, w_011_743);
  nand2 I027_044(w_027_044, w_019_538, w_015_261);
  or2  I027_048(w_027_048, w_017_1430, w_019_296);
  or2  I027_052(w_027_052, w_017_956, w_016_024);
  not1 I027_054(w_027_054, w_010_303);
  nand2 I027_057(w_027_057, w_001_728, w_007_211);
  not1 I027_059(w_027_059, w_008_798);
  or2  I027_061(w_027_061, w_002_241, w_014_300);
  not1 I027_062(w_027_062, w_022_279);
  not1 I027_063(w_027_063, w_012_211);
  or2  I027_065(w_027_065, w_026_1112, w_025_1533);
  and2 I027_067(w_027_067, w_011_114, w_005_309);
  or2  I027_069(w_027_069, w_022_409, w_009_053);
  nand2 I027_074(w_027_074, w_004_1678, w_026_1135);
  nand2 I027_076(w_027_076, w_022_047, w_006_186);
  and2 I027_077(w_027_077, w_010_029, w_022_009);
  not1 I027_079(w_027_079, w_021_022);
  or2  I027_081(w_027_081, w_004_655, w_003_262);
  not1 I027_082(w_027_082, w_015_266);
  or2  I027_091(w_027_091, w_000_1231, w_025_007);
  nand2 I027_093(w_027_093, w_012_406, w_010_174);
  nand2 I027_097(w_027_097, w_026_189, w_016_028);
  not1 I027_102(w_027_102, w_001_110);
  and2 I027_105(w_027_105, w_010_295, w_018_244);
  and2 I027_107(w_027_107, w_006_330, w_008_772);
  or2  I027_108(w_027_108, w_005_1163, w_013_164);
  not1 I027_109(w_027_109, w_003_056);
  and2 I027_110(w_027_110, w_019_897, w_004_551);
  or2  I027_114(w_027_114, w_005_283, w_010_212);
  not1 I027_117(w_027_117, w_005_1646);
  and2 I027_120(w_027_120, w_009_110, w_020_573);
  or2  I027_122(w_027_122, w_017_1143, w_021_002);
  and2 I027_129(w_027_129, w_020_465, w_018_186);
  or2  I027_130(w_027_130, w_005_584, w_014_300);
  nand2 I027_132(w_027_132, w_021_171, w_008_399);
  or2  I027_143(w_027_143, w_012_659, w_022_108);
  and2 I027_144(w_027_144, w_001_308, w_019_836);
  nand2 I027_145(w_027_145, w_008_552, w_007_1120);
  nand2 I027_146(w_027_146, w_020_599, w_005_095);
  nand2 I027_147(w_027_147, w_009_053, w_023_682);
  not1 I027_149(w_027_149, w_017_089);
  or2  I027_150(w_027_150, w_001_1076, w_001_543);
  or2  I027_155(w_027_155, w_014_417, w_006_127);
  and2 I027_157(w_027_157, w_006_279, w_023_278);
  not1 I027_158(w_027_158, w_006_015);
  or2  I027_159(w_027_159, w_020_292, w_017_678);
  not1 I027_160(w_027_160, w_003_152);
  and2 I027_161(w_027_161, w_001_052, w_002_253);
  and2 I027_163(w_027_163, w_016_038, w_019_1037);
  and2 I027_167(w_027_167, w_005_1380, w_023_1572);
  or2  I027_172(w_027_172, w_023_921, w_020_685);
  or2  I027_174(w_027_174, w_019_918, w_011_810);
  or2  I027_175(w_027_175, w_007_298, w_010_246);
  nand2 I027_176(w_027_176, w_018_066, w_019_441);
  not1 I027_178(w_027_178, w_016_025);
  nand2 I027_180(w_027_180, w_019_1029, w_004_1404);
  or2  I027_182(w_027_182, w_002_032, w_016_033);
  or2  I027_183(w_027_183, w_024_503, w_008_435);
  nand2 I027_184(w_027_184, w_003_255, w_019_1017);
  nand2 I027_186(w_027_186, w_012_591, w_009_056);
  and2 I027_187(w_027_187, w_013_132, w_022_085);
  and2 I027_190(w_027_190, w_016_021, w_007_113);
  and2 I027_198(w_027_198, w_022_072, w_010_067);
  not1 I027_199(w_027_199, w_015_158);
  nand2 I027_201(w_027_201, w_013_113, w_024_425);
  not1 I027_203(w_027_203, w_024_917);
  not1 I027_204(w_027_204, w_023_1013);
  or2  I027_207(w_027_207, w_020_277, w_024_200);
  not1 I027_209(w_027_209, w_013_332);
  nand2 I027_210(w_027_210, w_017_229, w_013_013);
  nand2 I027_211(w_027_211, w_024_688, w_015_056);
  or2  I027_214(w_027_214, w_020_240, w_016_009);
  not1 I027_215(w_027_215, w_008_369);
  or2  I027_218(w_027_218, w_000_1248, w_017_352);
  not1 I027_219(w_027_219, w_004_642);
  nand2 I027_220(w_027_220, w_007_267, w_021_090);
  and2 I027_226(w_027_226, w_003_051, w_010_027);
  nand2 I027_229(w_027_229, w_016_005, w_017_933);
  nand2 I027_231(w_027_231, w_026_366, w_006_266);
  nand2 I027_236(w_027_236, w_003_018, w_026_468);
  or2  I027_237(w_027_237, w_023_135, w_016_037);
  nand2 I027_242(w_027_242, w_011_070, w_014_264);
  and2 I027_243(w_027_243, w_001_003, w_012_403);
  and2 I027_246(w_027_246, w_004_737, w_019_705);
  and2 I027_247(w_027_247, w_002_588, w_019_359);
  and2 I027_249(w_027_249, w_018_227, w_016_033);
  or2  I027_258(w_027_258, w_019_819, w_012_465);
  and2 I027_261(w_027_261, w_008_445, w_004_1330);
  and2 I027_272(w_027_272, w_012_394, w_008_125);
  or2  I027_276(w_027_276, w_003_176, w_002_344);
  and2 I027_277(w_027_277, w_005_344, w_005_208);
  nand2 I027_279(w_027_279, w_018_059, w_010_382);
  not1 I027_280(w_027_280, w_003_245);
  and2 I027_286(w_027_286, w_006_135, w_015_266);
  or2  I027_287(w_027_287, w_007_015, w_023_1380);
  or2  I027_288(w_027_288, w_007_1060, w_016_021);
  not1 I027_297(w_027_297, w_005_1047);
  not1 I027_301(w_027_301, w_024_563);
  or2  I027_303(w_027_303, w_014_672, w_013_316);
  and2 I027_308(w_027_308, w_002_011, w_026_639);
  and2 I027_318(w_027_318, w_011_485, w_003_067);
  nand2 I027_319(w_027_319, w_016_015, w_011_117);
  nand2 I027_322(w_027_322, w_005_1271, w_020_923);
  and2 I027_323(w_027_323, w_019_081, w_020_351);
  and2 I027_326(w_027_326, w_023_733, w_025_961);
  and2 I027_328(w_027_328, w_018_073, w_025_1241);
  nand2 I027_334(w_027_334, w_009_098, w_009_103);
  nand2 I027_335(w_027_335, w_002_238, w_022_093);
  or2  I027_344(w_027_344, w_019_360, w_005_926);
  nand2 I027_345(w_027_345, w_005_1430, w_018_031);
  nand2 I027_347(w_027_347, w_018_015, w_002_078);
  and2 I027_348(w_027_348, w_014_163, w_023_331);
  and2 I027_351(w_027_351, w_014_508, w_026_416);
  not1 I027_356(w_027_356, w_026_238);
  or2  I027_362(w_027_362, w_012_011, w_007_208);
  not1 I027_364(w_027_364, w_002_331);
  not1 I027_366(w_027_366, w_021_015);
  not1 I027_370(w_027_370, w_000_1795);
  not1 I027_371(w_027_371, w_007_026);
  and2 I027_374(w_027_374, w_009_095, w_014_106);
  nand2 I027_376(w_027_376, w_016_007, w_003_043);
  or2  I027_380(w_027_380, w_000_1802, w_018_089);
  not1 I027_383(w_027_383, w_014_290);
  nand2 I027_384(w_027_384, w_010_046, w_024_1226);
  nand2 I027_387(w_027_387, w_011_845, w_007_1615);
  nand2 I027_389(w_027_389, w_010_160, w_023_1116);
  or2  I027_393(w_027_393, w_005_303, w_016_030);
  or2  I027_394(w_027_394, w_001_1369, w_002_491);
  or2  I027_395(w_027_395, w_000_1527, w_011_568);
  not1 I027_396(w_027_396, w_022_331);
  not1 I027_397(w_027_397, w_020_746);
  nand2 I027_398(w_027_398, w_025_1036, w_021_107);
  and2 I027_403(w_027_403, w_003_306, w_005_1487);
  not1 I027_407(w_027_407, w_008_853);
  or2  I027_408(w_027_408, w_012_188, w_024_585);
  and2 I027_409(w_027_409, w_023_077, w_022_369);
  or2  I027_411(w_027_411, w_004_1265, w_022_098);
  nand2 I027_413(w_027_413, w_000_203, w_010_399);
  or2  I027_414(w_027_414, w_014_197, w_018_029);
  nand2 I027_417(w_027_417, w_004_235, w_010_158);
  nand2 I027_419(w_027_419, w_008_657, w_026_404);
  and2 I027_421(w_027_421, w_007_002, w_017_734);
  and2 I027_422(w_027_422, w_009_018, w_007_1036);
  and2 I027_427(w_027_427, w_026_695, w_004_871);
  and2 I027_429(w_027_429, w_021_094, w_008_207);
  nand2 I027_430(w_027_430, w_002_022, w_004_1887);
  and2 I027_436(w_027_436, w_023_791, w_010_136);
  nand2 I027_437(w_027_437, w_002_110, w_009_107);
  and2 I027_440(w_027_440, w_007_1459, w_011_304);
  or2  I027_443(w_027_443, w_005_876, w_002_535);
  not1 I027_444(w_027_444, w_011_338);
  and2 I027_447(w_027_447, w_006_127, w_021_069);
  or2  I027_451(w_027_451, w_002_434, w_007_891);
  nand2 I027_456(w_027_456, w_017_985, w_013_298);
  not1 I027_458(w_027_458, w_002_168);
  or2  I027_459(w_027_459, w_026_155, w_010_292);
  or2  I027_460(w_027_460, w_007_267, w_024_265);
  nand2 I027_461(w_027_461, w_002_290, w_002_006);
  and2 I027_465(w_027_465, w_018_018, w_017_057);
  nand2 I027_467(w_027_467, w_013_288, w_017_162);
  nand2 I027_469(w_027_469, w_006_277, w_016_038);
  nand2 I027_470(w_027_470, w_022_084, w_008_108);
  not1 I027_472(w_027_472, w_005_1077);
  or2  I027_475(w_027_475, w_003_042, w_021_261);
  not1 I027_476(w_027_476, w_017_624);
  nand2 I027_481(w_027_481, w_010_244, w_000_1760);
  nand2 I027_482(w_027_482, w_002_233, w_013_009);
  nand2 I027_493(w_027_493, w_009_057, w_025_000);
  not1 I027_496(w_027_496, w_014_262);
  nand2 I027_498(w_027_498, w_020_456, w_025_1006);
  not1 I027_507(w_027_507, w_005_159);
  or2  I027_509(w_027_509, w_021_214, w_001_629);
  not1 I027_512(w_027_512, w_009_076);
  or2  I027_513(w_027_513, w_020_204, w_000_1142);
  or2  I027_516(w_027_516, w_018_133, w_004_369);
  nand2 I027_521(w_027_521, w_007_364, w_021_015);
  not1 I027_523(w_027_523, w_024_403);
  or2  I027_524(w_027_524, w_001_597, w_019_656);
  or2  I027_529(w_027_529, w_019_290, w_025_810);
  nand2 I027_530(w_027_530, w_022_307, w_006_246);
  not1 I027_531(w_027_531, w_024_528);
  or2  I027_533(w_027_533, w_007_599, w_008_838);
  nand2 I027_536(w_027_536, w_003_280, w_019_655);
  and2 I027_543(w_027_543, w_004_1380, w_021_006);
  and2 I027_547(w_027_547, w_025_422, w_013_052);
  not1 I027_550(w_027_550, w_009_003);
  not1 I027_552(w_027_552, w_017_1327);
  and2 I027_553(w_027_553, w_018_261, w_020_880);
  not1 I027_556(w_027_556, w_005_057);
  and2 I027_558(w_027_558, w_007_1620, w_018_168);
  nand2 I027_560(w_027_560, w_020_527, w_008_551);
  and2 I027_563(w_027_563, w_014_561, w_003_076);
  and2 I027_564(w_027_564, w_002_057, w_004_041);
  nand2 I027_565(w_027_565, w_012_561, w_020_466);
  not1 I027_567(w_027_567, w_026_1080);
  and2 I027_571(w_027_571, w_010_008, w_009_086);
  and2 I027_572(w_027_572, w_002_353, w_007_034);
  and2 I027_574(w_027_574, w_004_1382, w_018_050);
  not1 I027_575(w_027_575, w_024_685);
  or2  I027_578(w_027_578, w_004_380, w_015_216);
  and2 I027_579(w_027_579, w_006_131, w_007_275);
  nand2 I027_580(w_027_580, w_016_020, w_004_852);
  nand2 I027_583(w_027_583, w_026_075, w_022_289);
  and2 I027_584(w_027_584, w_001_1651, w_015_060);
  nand2 I027_585(w_027_585, w_005_242, w_011_038);
  or2  I027_587(w_027_587, w_017_1910, w_020_551);
  or2  I027_588(w_027_588, w_014_713, w_018_175);
  or2  I027_590(w_027_590, w_003_181, w_026_1182);
  and2 I027_591(w_027_591, w_003_256, w_003_135);
  or2  I028_000(w_028_000, w_018_082, w_023_903);
  and2 I028_001(w_028_001, w_021_238, w_012_231);
  nand2 I028_002(w_028_002, w_022_201, w_018_265);
  nand2 I028_004(w_028_004, w_012_571, w_000_073);
  and2 I028_007(w_028_007, w_024_772, w_005_299);
  and2 I028_010(w_028_010, w_022_381, w_011_698);
  nand2 I028_018(w_028_018, w_013_191, w_019_204);
  nand2 I028_022(w_028_022, w_020_431, w_003_187);
  not1 I028_024(w_028_024, w_014_659);
  and2 I028_025(w_028_025, w_024_1230, w_025_070);
  not1 I028_026(w_028_026, w_017_1881);
  and2 I028_028(w_028_028, w_014_184, w_024_857);
  not1 I028_029(w_028_029, w_009_073);
  nand2 I028_035(w_028_035, w_027_443, w_009_061);
  and2 I028_038(w_028_038, w_000_081, w_004_1852);
  or2  I028_041(w_028_041, w_018_215, w_004_068);
  not1 I028_046(w_028_046, w_017_1322);
  and2 I028_049(w_028_049, w_019_023, w_004_1098);
  or2  I028_051(w_028_051, w_015_250, w_011_707);
  nand2 I028_054(w_028_054, w_027_187, w_009_035);
  not1 I028_056(w_028_056, w_018_195);
  nand2 I028_061(w_028_061, w_015_151, w_006_214);
  and2 I028_062(w_028_062, w_026_1109, w_002_288);
  not1 I028_064(w_028_064, w_007_241);
  or2  I028_066(w_028_066, w_022_027, w_025_1002);
  or2  I028_067(w_028_067, w_027_215, w_016_016);
  not1 I028_070(w_028_070, w_001_531);
  or2  I028_071(w_028_071, w_020_694, w_008_002);
  nand2 I028_076(w_028_076, w_012_141, w_001_817);
  and2 I028_077(w_028_077, w_018_012, w_005_1266);
  and2 I028_079(w_028_079, w_001_013, w_026_1226);
  or2  I028_082(w_028_082, w_016_025, w_022_018);
  and2 I028_083(w_028_083, w_023_039, w_006_072);
  or2  I028_084(w_028_084, w_014_091, w_006_232);
  and2 I028_087(w_028_087, w_026_117, w_013_036);
  nand2 I028_088(w_028_088, w_022_236, w_021_065);
  nand2 I028_092(w_028_092, w_007_1331, w_010_231);
  not1 I028_094(w_028_094, w_022_159);
  and2 I028_095(w_028_095, w_018_081, w_022_029);
  not1 I028_097(w_028_097, w_025_099);
  or2  I028_098(w_028_098, w_026_987, w_018_068);
  and2 I028_102(w_028_102, w_001_572, w_024_929);
  nand2 I028_106(w_028_106, w_002_523, w_011_133);
  nand2 I028_108(w_028_108, w_020_701, w_010_197);
  or2  I028_111(w_028_111, w_016_036, w_012_221);
  nand2 I028_112(w_028_112, w_007_903, w_015_105);
  or2  I028_114(w_028_114, w_022_097, w_026_597);
  and2 I028_116(w_028_116, w_005_1566, w_012_521);
  not1 I028_118(w_028_118, w_017_1242);
  not1 I028_119(w_028_119, w_024_146);
  or2  I028_120(w_028_120, w_001_518, w_011_132);
  and2 I028_124(w_028_124, w_025_1407, w_025_699);
  nand2 I028_126(w_028_126, w_016_038, w_014_648);
  not1 I028_130(w_028_130, w_027_567);
  nand2 I028_132(w_028_132, w_025_705, w_022_376);
  not1 I028_135(w_028_135, w_006_061);
  or2  I028_137(w_028_137, w_011_858, w_027_533);
  or2  I028_140(w_028_140, w_019_074, w_005_1165);
  or2  I028_145(w_028_145, w_018_022, w_004_030);
  nand2 I028_146(w_028_146, w_025_1243, w_012_504);
  or2  I028_149(w_028_149, w_016_023, w_013_179);
  nand2 I028_150(w_028_150, w_021_156, w_001_586);
  nand2 I028_152(w_028_152, w_001_673, w_023_710);
  not1 I028_155(w_028_155, w_015_045);
  not1 I028_157(w_028_157, w_021_266);
  or2  I028_158(w_028_158, w_012_042, w_020_112);
  or2  I028_159(w_028_159, w_022_347, w_013_024);
  nand2 I028_160(w_028_160, w_005_014, w_012_186);
  not1 I028_169(w_028_169, w_020_986);
  not1 I028_170(w_028_170, w_008_626);
  or2  I028_172(w_028_172, w_024_252, w_023_026);
  and2 I028_175(w_028_175, w_018_006, w_023_1455);
  nand2 I028_177(w_028_177, w_021_068, w_001_240);
  and2 I028_181(w_028_181, w_000_442, w_016_003);
  not1 I028_189(w_028_189, w_001_378);
  nand2 I028_191(w_028_191, w_007_264, w_001_1470);
  not1 I028_194(w_028_194, w_015_047);
  and2 I028_195(w_028_195, w_005_049, w_006_215);
  and2 I028_197(w_028_197, w_011_660, w_010_001);
  not1 I028_204(w_028_204, w_021_203);
  or2  I028_209(w_028_209, w_023_1218, w_016_007);
  and2 I028_217(w_028_217, w_027_396, w_005_534);
  or2  I028_219(w_028_219, w_006_175, w_001_809);
  or2  I028_223(w_028_223, w_021_085, w_013_000);
  and2 I028_231(w_028_231, w_003_058, w_005_802);
  or2  I028_236(w_028_236, w_012_025, w_014_588);
  or2  I028_237(w_028_237, w_007_726, w_021_256);
  or2  I028_243(w_028_243, w_022_404, w_023_198);
  not1 I028_244(w_028_244, w_014_092);
  not1 I028_247(w_028_247, w_018_273);
  and2 I028_251(w_028_251, w_024_976, w_020_401);
  not1 I028_253(w_028_253, w_025_006);
  and2 I028_256(w_028_256, w_006_274, w_007_851);
  and2 I028_257(w_028_257, w_017_551, w_004_933);
  nand2 I028_258(w_028_258, w_008_609, w_010_345);
  not1 I028_266(w_028_266, w_021_002);
  not1 I028_267(w_028_267, w_023_736);
  not1 I028_275(w_028_275, w_009_000);
  and2 I028_277(w_028_277, w_012_629, w_001_1485);
  and2 I028_279(w_028_279, w_011_250, w_023_1553);
  and2 I028_280(w_028_280, w_020_343, w_016_019);
  nand2 I028_285(w_028_285, w_012_632, w_011_800);
  not1 I028_287(w_028_287, w_027_323);
  and2 I028_292(w_028_292, w_008_111, w_004_588);
  and2 I028_298(w_028_298, w_019_339, w_008_515);
  nand2 I028_300(w_028_300, w_002_119, w_020_269);
  or2  I028_301(w_028_301, w_014_746, w_014_263);
  or2  I028_311(w_028_311, w_013_025, w_019_011);
  not1 I028_313(w_028_313, w_000_1379);
  nand2 I028_317(w_028_317, w_012_317, w_021_203);
  or2  I028_319(w_028_319, w_026_189, w_016_001);
  and2 I028_323(w_028_323, w_001_1425, w_017_1871);
  nand2 I028_325(w_028_325, w_013_119, w_018_274);
  and2 I028_335(w_028_335, w_026_1455, w_023_496);
  and2 I028_340(w_028_340, w_024_1190, w_005_543);
  not1 I028_342(w_028_342, w_016_003);
  and2 I028_346(w_028_346, w_015_124, w_002_583);
  or2  I028_353(w_028_353, w_019_671, w_007_199);
  or2  I028_355(w_028_355, w_025_777, w_019_406);
  not1 I028_365(w_028_365, w_023_914);
  not1 I028_373(w_028_373, w_016_002);
  or2  I028_380(w_028_380, w_009_053, w_009_093);
  or2  I028_381(w_028_381, w_007_399, w_018_089);
  or2  I028_384(w_028_384, w_009_052, w_018_018);
  or2  I028_397(w_028_397, w_019_232, w_000_1612);
  nand2 I028_399(w_028_399, w_025_1391, w_020_201);
  and2 I028_404(w_028_404, w_005_1141, w_012_390);
  or2  I028_409(w_028_409, w_002_235, w_000_1568);
  nand2 I028_414(w_028_414, w_003_073, w_000_476);
  and2 I028_418(w_028_418, w_005_154, w_019_627);
  and2 I028_420(w_028_420, w_006_322, w_025_034);
  nand2 I028_426(w_028_426, w_026_815, w_015_041);
  or2  I028_430(w_028_430, w_005_1143, w_004_1283);
  not1 I028_435(w_028_435, w_027_117);
  or2  I028_453(w_028_453, w_022_175, w_013_212);
  nand2 I028_454(w_028_454, w_012_390, w_014_195);
  or2  I028_461(w_028_461, w_000_401, w_001_093);
  or2  I028_463(w_028_463, w_008_281, w_019_526);
  or2  I028_465(w_028_465, w_013_133, w_024_682);
  or2  I028_469(w_028_469, w_013_051, w_006_289);
  or2  I028_470(w_028_470, w_009_048, w_007_546);
  nand2 I028_472(w_028_472, w_005_525, w_020_730);
  not1 I028_473(w_028_473, w_024_189);
  nand2 I028_479(w_028_479, w_026_572, w_020_544);
  or2  I028_480(w_028_480, w_010_069, w_017_142);
  and2 I028_485(w_028_485, w_001_805, w_003_135);
  or2  I028_491(w_028_491, w_015_022, w_005_780);
  nand2 I028_495(w_028_495, w_017_1269, w_025_839);
  or2  I028_513(w_028_513, w_000_1049, w_000_792);
  nand2 I028_516(w_028_516, w_010_077, w_024_1557);
  not1 I028_526(w_028_526, w_004_804);
  nand2 I028_528(w_028_528, w_020_473, w_010_177);
  and2 I028_529(w_028_529, w_024_621, w_011_263);
  or2  I028_530(w_028_530, w_016_001, w_000_735);
  nand2 I028_541(w_028_541, w_006_069, w_004_234);
  nand2 I028_546(w_028_546, w_010_124, w_023_1098);
  not1 I028_549(w_028_549, w_016_028);
  or2  I028_552(w_028_552, w_020_416, w_005_770);
  nand2 I028_553(w_028_553, w_027_158, w_022_197);
  not1 I028_557(w_028_557, w_022_026);
  not1 I028_565(w_028_565, w_022_283);
  nand2 I028_566(w_028_566, w_013_252, w_012_395);
  and2 I028_568(w_028_568, w_011_533, w_003_091);
  not1 I028_580(w_028_580, w_003_314);
  or2  I028_581(w_028_581, w_009_098, w_024_318);
  nand2 I028_583(w_028_583, w_009_078, w_015_178);
  nand2 I028_586(w_028_586, w_019_590, w_001_758);
  not1 I028_589(w_028_589, w_009_025);
  nand2 I028_592(w_028_592, w_006_074, w_010_046);
  or2  I028_595(w_028_595, w_006_054, w_011_659);
  or2  I028_610(w_028_610, w_025_180, w_026_152);
  not1 I028_619(w_028_619, w_002_196);
  not1 I028_622(w_028_622, w_013_023);
  and2 I028_623(w_028_623, w_001_1592, w_015_252);
  not1 I028_624(w_028_624, w_023_336);
  not1 I028_626(w_028_626, w_019_657);
  not1 I028_630(w_028_630, w_007_406);
  and2 I028_633(w_028_633, w_022_238, w_009_108);
  or2  I028_636(w_028_636, w_014_158, w_003_041);
  and2 I028_638(w_028_638, w_000_1033, w_006_103);
  not1 I028_639(w_028_639, w_007_1086);
  nand2 I028_641(w_028_641, w_008_160, w_006_007);
  or2  I028_647(w_028_647, w_025_100, w_024_577);
  not1 I028_648(w_028_648, w_003_041);
  not1 I028_653(w_028_653, w_018_039);
  not1 I028_655(w_028_655, w_018_156);
  and2 I028_664(w_028_664, w_018_219, w_021_237);
  and2 I028_666(w_028_666, w_019_617, w_007_289);
  or2  I028_668(w_028_668, w_014_019, w_007_130);
  nand2 I028_670(w_028_670, w_013_153, w_024_337);
  not1 I028_671(w_028_671, w_017_1058);
  not1 I028_674(w_028_674, w_009_108);
  not1 I028_678(w_028_678, w_013_150);
  and2 I028_680(w_028_680, w_006_086, w_012_350);
  nand2 I028_683(w_028_683, w_004_415, w_016_008);
  and2 I028_690(w_028_690, w_011_840, w_013_109);
  nand2 I028_698(w_028_698, w_022_004, w_024_927);
  and2 I028_704(w_028_704, w_023_1294, w_020_939);
  or2  I028_705(w_028_705, w_024_022, w_026_1356);
  or2  I028_706(w_028_706, w_019_843, w_010_211);
  or2  I028_714(w_028_714, w_016_009, w_018_044);
  or2  I028_716(w_028_716, w_020_314, w_022_089);
  not1 I028_719(w_028_719, w_011_522);
  or2  I028_721(w_028_721, w_006_128, w_005_433);
  not1 I028_722(w_028_722, w_022_178);
  not1 I028_725(w_028_725, w_002_402);
  not1 I028_727(w_028_727, w_008_201);
  nand2 I028_731(w_028_731, w_016_034, w_003_063);
  or2  I028_735(w_028_735, w_002_406, w_013_185);
  and2 I028_748(w_028_748, w_016_012, w_026_838);
  not1 I028_757(w_028_757, w_007_278);
  or2  I028_760(w_028_760, w_001_1520, w_012_409);
  nand2 I028_763(w_028_763, w_017_390, w_006_101);
  and2 I028_764(w_028_764, w_000_1463, w_023_072);
  or2  I028_766(w_028_766, w_026_134, w_006_227);
  not1 I028_767(w_028_767, w_018_261);
  or2  I028_768(w_028_768, w_026_515, w_002_467);
  or2  I028_777(w_028_777, w_024_506, w_010_263);
  not1 I028_780(w_028_780, w_024_1555);
  nand2 I028_783(w_028_783, w_000_1810, w_013_047);
  not1 I028_795(w_028_795, w_025_1375);
  and2 I028_798(w_028_798, w_019_486, w_000_570);
  or2  I028_801(w_028_801, w_026_1347, w_020_452);
  or2  I028_805(w_028_805, w_010_400, w_013_027);
  and2 I028_809(w_028_809, w_012_631, w_027_247);
  nand2 I028_813(w_028_813, w_025_515, w_003_280);
  or2  I028_814(w_028_814, w_023_515, w_011_077);
  nand2 I028_823(w_028_823, w_013_227, w_018_048);
  and2 I028_826(w_028_826, w_000_709, w_023_212);
  nand2 I028_829(w_028_829, w_023_353, w_018_077);
  nand2 I028_832(w_028_832, w_000_012, w_007_252);
  or2  I028_847(w_028_847, w_004_1255, w_023_1604);
  or2  I028_851(w_028_851, w_016_005, w_005_669);
  or2  I028_852(w_028_852, w_000_363, w_017_1753);
  or2  I028_853(w_028_853, w_006_313, w_016_037);
  nand2 I028_855(w_028_855, w_015_274, w_004_1364);
  nand2 I028_863(w_028_863, w_016_001, w_004_563);
  nand2 I028_866(w_028_866, w_027_062, w_016_025);
  nand2 I028_871(w_028_871, w_010_295, w_021_174);
  nand2 I028_873(w_028_873, w_013_078, w_011_498);
  and2 I028_874(w_028_874, w_026_658, w_025_1412);
  not1 I028_876(w_028_876, w_014_412);
  or2  I028_880(w_028_880, w_011_592, w_005_1297);
  not1 I028_889(w_028_889, w_013_188);
  or2  I028_907(w_028_907, w_001_341, w_014_018);
  nand2 I029_003(w_029_003, w_022_212, w_010_091);
  and2 I029_004(w_029_004, w_008_830, w_002_225);
  not1 I029_005(w_029_005, w_006_106);
  not1 I029_014(w_029_014, w_012_637);
  not1 I029_017(w_029_017, w_014_177);
  and2 I029_020(w_029_020, w_003_254, w_015_271);
  not1 I029_022(w_029_022, w_014_189);
  and2 I029_032(w_029_032, w_017_871, w_009_063);
  nand2 I029_033(w_029_033, w_014_512, w_002_572);
  or2  I029_036(w_029_036, w_024_029, w_028_832);
  not1 I029_039(w_029_039, w_006_180);
  nand2 I029_040(w_029_040, w_014_116, w_019_019);
  nand2 I029_042(w_029_042, w_026_1305, w_003_187);
  and2 I029_047(w_029_047, w_027_467, w_000_1121);
  and2 I029_051(w_029_051, w_025_734, w_002_137);
  not1 I029_053(w_029_053, w_010_354);
  not1 I029_061(w_029_061, w_017_929);
  not1 I029_070(w_029_070, w_008_088);
  not1 I029_072(w_029_072, w_022_025);
  nand2 I029_073(w_029_073, w_014_118, w_005_1602);
  nand2 I029_077(w_029_077, w_000_1232, w_003_129);
  and2 I029_083(w_029_083, w_008_428, w_018_004);
  not1 I029_084(w_029_084, w_008_425);
  or2  I029_085(w_029_085, w_017_1357, w_018_201);
  not1 I029_088(w_029_088, w_005_415);
  nand2 I029_090(w_029_090, w_000_778, w_011_381);
  or2  I029_092(w_029_092, w_017_253, w_002_374);
  nand2 I029_095(w_029_095, w_028_094, w_004_1848);
  or2  I029_098(w_029_098, w_021_157, w_022_031);
  nand2 I029_105(w_029_105, w_007_1117, w_021_151);
  not1 I029_106(w_029_106, w_018_147);
  not1 I029_110(w_029_110, w_013_205);
  not1 I029_113(w_029_113, w_003_092);
  or2  I029_119(w_029_119, w_007_883, w_006_328);
  and2 I029_125(w_029_125, w_010_222, w_006_127);
  or2  I029_129(w_029_129, w_017_977, w_011_504);
  and2 I029_130(w_029_130, w_002_130, w_024_1572);
  and2 I029_132(w_029_132, w_027_011, w_011_785);
  and2 I029_133(w_029_133, w_026_750, w_022_398);
  and2 I029_135(w_029_135, w_017_1612, w_004_566);
  and2 I029_136(w_029_136, w_000_687, w_012_413);
  not1 I029_142(w_029_142, w_016_029);
  nand2 I029_143(w_029_143, w_008_717, w_006_268);
  and2 I029_146(w_029_146, w_007_353, w_023_040);
  not1 I029_148(w_029_148, w_008_039);
  not1 I029_149(w_029_149, w_001_192);
  or2  I029_151(w_029_151, w_016_014, w_015_003);
  or2  I029_163(w_029_163, w_019_1060, w_010_021);
  and2 I029_164(w_029_164, w_008_279, w_005_1219);
  nand2 I029_165(w_029_165, w_011_328, w_021_077);
  not1 I029_166(w_029_166, w_002_193);
  not1 I029_178(w_029_178, w_004_1381);
  not1 I029_180(w_029_180, w_007_218);
  not1 I029_187(w_029_187, w_019_631);
  and2 I029_188(w_029_188, w_025_795, w_020_249);
  not1 I029_193(w_029_193, w_015_010);
  not1 I029_202(w_029_202, w_014_247);
  not1 I029_206(w_029_206, w_006_239);
  nand2 I029_210(w_029_210, w_013_106, w_023_498);
  nand2 I029_211(w_029_211, w_022_412, w_023_070);
  and2 I029_213(w_029_213, w_012_521, w_015_093);
  and2 I029_215(w_029_215, w_025_355, w_021_119);
  nand2 I029_220(w_029_220, w_017_730, w_020_939);
  and2 I029_227(w_029_227, w_028_150, w_021_233);
  not1 I029_233(w_029_233, w_011_822);
  not1 I029_242(w_029_242, w_021_273);
  and2 I029_243(w_029_243, w_007_055, w_010_184);
  nand2 I029_244(w_029_244, w_026_830, w_010_067);
  and2 I029_245(w_029_245, w_014_132, w_007_174);
  nand2 I029_250(w_029_250, w_020_388, w_013_314);
  and2 I029_251(w_029_251, w_002_308, w_014_059);
  or2  I029_256(w_029_256, w_009_031, w_011_051);
  or2  I029_258(w_029_258, w_026_1071, w_009_106);
  and2 I029_263(w_029_263, w_018_218, w_019_656);
  not1 I029_273(w_029_273, w_010_309);
  and2 I029_274(w_029_274, w_028_461, w_005_395);
  not1 I029_277(w_029_277, w_019_632);
  nand2 I029_281(w_029_281, w_026_457, w_026_376);
  or2  I029_283(w_029_283, w_016_002, w_019_150);
  nand2 I029_291(w_029_291, w_002_473, w_002_223);
  and2 I029_296(w_029_296, w_004_1239, w_017_003);
  not1 I029_300(w_029_300, w_028_353);
  or2  I029_305(w_029_305, w_024_1649, w_024_134);
  and2 I029_307(w_029_307, w_016_023, w_026_136);
  not1 I029_308(w_029_308, w_010_231);
  and2 I029_311(w_029_311, w_002_336, w_020_995);
  not1 I029_319(w_029_319, w_025_1304);
  not1 I029_328(w_029_328, w_000_1008);
  and2 I029_329(w_029_329, w_019_021, w_027_003);
  not1 I029_332(w_029_332, w_025_1495);
  or2  I029_347(w_029_347, w_004_1235, w_028_876);
  not1 I029_354(w_029_354, w_008_224);
  and2 I029_365(w_029_365, w_018_017, w_003_153);
  and2 I029_367(w_029_367, w_024_1642, w_004_1802);
  and2 I029_377(w_029_377, w_001_1548, w_005_602);
  and2 I029_383(w_029_383, w_024_016, w_010_004);
  nand2 I029_387(w_029_387, w_020_152, w_003_015);
  not1 I029_389(w_029_389, w_023_064);
  not1 I029_391(w_029_391, w_011_201);
  or2  I029_394(w_029_394, w_018_237, w_013_061);
  not1 I029_399(w_029_399, w_014_405);
  or2  I029_402(w_029_402, w_003_083, w_005_015);
  or2  I029_414(w_029_414, w_017_485, w_024_088);
  and2 I029_416(w_029_416, w_020_375, w_014_261);
  and2 I029_429(w_029_429, w_023_1065, w_005_070);
  nand2 I029_440(w_029_440, w_012_144, w_014_711);
  not1 I029_444(w_029_444, w_022_356);
  not1 I029_450(w_029_450, w_001_133);
  nand2 I029_453(w_029_453, w_004_015, w_027_102);
  nand2 I029_468(w_029_468, w_027_147, w_010_350);
  nand2 I029_470(w_029_470, w_019_917, w_014_387);
  not1 I029_471(w_029_471, w_000_1451);
  nand2 I029_474(w_029_474, w_004_843, w_024_882);
  or2  I029_475(w_029_475, w_001_303, w_009_088);
  nand2 I029_476(w_029_476, w_027_547, w_023_596);
  not1 I029_477(w_029_477, w_005_1513);
  nand2 I029_486(w_029_486, w_023_1196, w_010_347);
  not1 I029_490(w_029_490, w_028_705);
  nand2 I029_494(w_029_494, w_003_067, w_008_616);
  not1 I029_496(w_029_496, w_025_082);
  and2 I029_502(w_029_502, w_026_291, w_014_133);
  or2  I029_504(w_029_504, w_020_755, w_028_130);
  not1 I029_507(w_029_507, w_001_276);
  not1 I029_509(w_029_509, w_021_204);
  or2  I029_511(w_029_511, w_019_339, w_025_492);
  or2  I029_516(w_029_516, w_018_241, w_019_583);
  nand2 I029_524(w_029_524, w_004_449, w_009_019);
  or2  I029_529(w_029_529, w_007_980, w_011_206);
  and2 I029_532(w_029_532, w_014_662, w_006_050);
  nand2 I029_533(w_029_533, w_028_795, w_013_120);
  not1 I029_538(w_029_538, w_002_190);
  not1 I029_539(w_029_539, w_001_061);
  and2 I029_541(w_029_541, w_026_725, w_022_232);
  nand2 I029_547(w_029_547, w_013_177, w_021_186);
  or2  I029_548(w_029_548, w_011_051, w_017_821);
  nand2 I029_550(w_029_550, w_026_510, w_013_244);
  nand2 I029_552(w_029_552, w_019_092, w_011_325);
  nand2 I029_553(w_029_553, w_011_395, w_028_619);
  not1 I029_554(w_029_554, w_023_117);
  nand2 I029_557(w_029_557, w_024_596, w_024_179);
  nand2 I029_565(w_029_565, w_018_160, w_009_000);
  nand2 I029_567(w_029_567, w_007_027, w_005_390);
  or2  I029_568(w_029_568, w_005_1451, w_012_095);
  not1 I029_579(w_029_579, w_007_954);
  not1 I029_582(w_029_582, w_015_150);
  and2 I029_583(w_029_583, w_002_282, w_010_104);
  or2  I029_584(w_029_584, w_028_557, w_017_141);
  or2  I029_586(w_029_586, w_011_043, w_008_790);
  nand2 I029_589(w_029_589, w_015_172, w_004_910);
  or2  I029_594(w_029_594, w_018_028, w_028_866);
  nand2 I029_603(w_029_603, w_014_193, w_009_033);
  or2  I029_611(w_029_611, w_023_654, w_018_137);
  and2 I029_613(w_029_613, w_026_1044, w_024_111);
  or2  I029_614(w_029_614, w_016_035, w_014_211);
  not1 I029_615(w_029_615, w_027_571);
  not1 I029_622(w_029_622, w_002_164);
  and2 I029_626(w_029_626, w_001_799, w_028_768);
  nand2 I029_628(w_029_628, w_024_453, w_004_143);
  and2 I029_631(w_029_631, w_009_098, w_010_133);
  or2  I029_632(w_029_632, w_024_700, w_024_309);
  nand2 I029_637(w_029_637, w_013_002, w_006_294);
  nand2 I029_638(w_029_638, w_016_038, w_003_310);
  not1 I029_644(w_029_644, w_002_158);
  not1 I029_650(w_029_650, w_012_477);
  not1 I029_661(w_029_661, w_022_009);
  not1 I029_679(w_029_679, w_018_045);
  not1 I029_685(w_029_685, w_027_286);
  not1 I029_692(w_029_692, w_010_123);
  not1 I029_693(w_029_693, w_026_378);
  or2  I029_694(w_029_694, w_000_1682, w_006_107);
  and2 I029_709(w_029_709, w_022_200, w_002_192);
  not1 I029_715(w_029_715, w_024_089);
  nand2 I029_718(w_029_718, w_026_136, w_014_210);
  not1 I029_719(w_029_719, w_010_181);
  or2  I029_720(w_029_720, w_005_1418, w_020_1091);
  and2 I029_731(w_029_731, w_007_880, w_002_206);
  and2 I029_739(w_029_739, w_013_230, w_014_274);
  not1 I029_740(w_029_740, w_014_505);
  or2  I029_747(w_029_747, w_021_112, w_004_625);
  and2 I029_754(w_029_754, w_024_148, w_020_296);
  not1 I029_755(w_029_755, w_018_239);
  and2 I029_756(w_029_756, w_008_390, w_008_572);
  and2 I029_766(w_029_766, w_013_330, w_021_100);
  not1 I029_782(w_029_782, w_017_633);
  nand2 I029_792(w_029_792, w_016_004, w_019_894);
  nand2 I029_802(w_029_802, w_006_276, w_020_1072);
  not1 I029_810(w_029_810, w_025_455);
  not1 I029_836(w_029_836, w_005_477);
  not1 I029_837(w_029_837, w_003_032);
  or2  I029_849(w_029_849, w_026_123, w_022_398);
  not1 I029_856(w_029_856, w_022_265);
  or2  I029_887(w_029_887, w_008_373, w_010_131);
  and2 I029_892(w_029_892, w_014_569, w_016_011);
  and2 I029_899(w_029_899, w_013_280, w_015_112);
  nand2 I029_901(w_029_901, w_025_725, w_004_856);
  or2  I029_904(w_029_904, w_008_344, w_014_295);
  and2 I029_911(w_029_911, w_020_794, w_016_014);
  and2 I029_921(w_029_921, w_001_454, w_023_1031);
  or2  I029_934(w_029_934, w_005_228, w_002_573);
  or2  I029_935(w_029_935, w_005_591, w_025_142);
  or2  I029_943(w_029_943, w_014_529, w_028_041);
  not1 I029_945(w_029_945, w_026_577);
  and2 I029_962(w_029_962, w_026_1159, w_009_087);
  and2 I029_970(w_029_970, w_007_261, w_001_016);
  nand2 I029_976(w_029_976, w_012_073, w_028_323);
  or2  I029_982(w_029_982, w_016_004, w_004_834);
  and2 I029_985(w_029_985, w_003_241, w_000_1149);
  or2  I029_987(w_029_987, w_023_826, w_010_113);
  and2 I029_998(w_029_998, w_016_017, w_007_1477);
  nand2 I029_999(w_029_999, w_002_068, w_019_139);
  nand2 I029_1002(w_029_1002, w_003_089, w_009_057);
  or2  I029_1003(w_029_1003, w_025_1432, w_013_315);
  or2  I029_1005(w_029_1005, w_020_449, w_010_336);
  nand2 I029_1006(w_029_1006, w_007_421, w_015_023);
  not1 I029_1053(w_029_1053, w_020_494);
  not1 I029_1057(w_029_1057, w_002_290);
  and2 I029_1059(w_029_1059, w_024_1320, w_011_227);
  or2  I029_1074(w_029_1074, w_027_395, w_024_351);
  or2  I029_1077(w_029_1077, w_021_055, w_023_318);
  and2 I029_1087(w_029_1087, w_019_292, w_005_251);
  and2 I029_1091(w_029_1091, w_024_1401, w_016_011);
  or2  I029_1092(w_029_1092, w_003_036, w_020_1108);
  or2  I029_1106(w_029_1106, w_007_860, w_007_216);
  not1 I029_1109(w_029_1109, w_024_1557);
  nand2 I029_1118(w_029_1118, w_023_206, w_025_1025);
  or2  I029_1124(w_029_1124, w_018_105, w_015_126);
  or2  I029_1126(w_029_1126, w_020_404, w_016_007);
  nand2 I029_1127(w_029_1127, w_022_348, w_013_101);
  and2 I029_1129(w_029_1129, w_011_097, w_015_172);
  or2  I029_1135(w_029_1135, w_020_839, w_019_244);
  or2  I029_1141(w_029_1141, w_005_387, w_002_395);
  not1 I029_1142(w_029_1142, w_021_195);
  or2  I029_1155(w_029_1155, w_003_044, w_015_219);
  nand2 I029_1159(w_029_1159, w_012_570, w_013_105);
  or2  I029_1170(w_029_1170, w_007_1605, w_005_295);
  and2 I029_1171(w_029_1171, w_009_106, w_026_022);
  not1 I029_1172(w_029_1172, w_020_312);
  and2 I029_1176(w_029_1176, w_011_060, w_006_250);
  or2  I029_1193(w_029_1193, w_013_239, w_025_335);
  nand2 I029_1207(w_029_1207, w_014_251, w_013_332);
  nand2 I029_1210(w_029_1210, w_012_176, w_013_284);
  and2 I029_1236(w_029_1236, w_021_057, w_028_626);
  and2 I029_1240(w_029_1240, w_008_216, w_026_1424);
  and2 I029_1244(w_029_1244, w_011_619, w_021_088);
  not1 I029_1245(w_029_1245, w_015_264);
  nand2 I029_1272(w_029_1272, w_014_736, w_000_768);
  not1 I029_1276(w_029_1276, w_002_149);
  or2  I029_1281(w_029_1281, w_007_879, w_027_163);
  nand2 I029_1296(w_029_1296, w_025_327, w_007_640);
  nand2 I029_1328(w_029_1328, w_007_311, w_007_207);
  or2  I029_1337(w_029_1337, w_002_368, w_004_080);
  nand2 I030_000(w_030_000, w_026_005, w_005_893);
  and2 I030_003(w_030_003, w_027_231, w_022_093);
  not1 I030_007(w_030_007, w_024_1006);
  and2 I030_012(w_030_012, w_014_353, w_004_318);
  and2 I030_016(w_030_016, w_021_218, w_007_108);
  nand2 I030_017(w_030_017, w_010_253, w_019_340);
  nand2 I030_019(w_030_019, w_001_454, w_004_1135);
  not1 I030_020(w_030_020, w_006_007);
  not1 I030_025(w_030_025, w_012_177);
  nand2 I030_038(w_030_038, w_026_073, w_017_1126);
  and2 I030_042(w_030_042, w_000_197, w_029_429);
  or2  I030_048(w_030_048, w_002_586, w_016_011);
  not1 I030_050(w_030_050, w_021_077);
  nand2 I030_055(w_030_055, w_009_011, w_001_533);
  not1 I030_059(w_030_059, w_024_757);
  not1 I030_065(w_030_065, w_000_1103);
  not1 I030_067(w_030_067, w_002_005);
  nand2 I030_069(w_030_069, w_005_682, w_014_582);
  and2 I030_070(w_030_070, w_013_227, w_003_043);
  nand2 I030_071(w_030_071, w_013_134, w_027_272);
  and2 I030_072(w_030_072, w_028_002, w_029_329);
  nand2 I030_073(w_030_073, w_004_416, w_009_066);
  or2  I030_078(w_030_078, w_008_136, w_009_012);
  and2 I030_079(w_030_079, w_029_250, w_027_016);
  nand2 I030_082(w_030_082, w_005_1656, w_023_250);
  and2 I030_083(w_030_083, w_023_269, w_006_326);
  nand2 I030_098(w_030_098, w_023_1313, w_015_287);
  and2 I030_102(w_030_102, w_005_156, w_026_601);
  or2  I030_105(w_030_105, w_018_100, w_000_412);
  nand2 I030_110(w_030_110, w_002_289, w_001_1671);
  or2  I030_112(w_030_112, w_002_111, w_005_1213);
  not1 I030_124(w_030_124, w_012_191);
  not1 I030_126(w_030_126, w_009_006);
  nand2 I030_127(w_030_127, w_002_217, w_024_468);
  nand2 I030_134(w_030_134, w_006_086, w_026_287);
  nand2 I030_140(w_030_140, w_026_1436, w_003_204);
  nand2 I030_146(w_030_146, w_012_168, w_011_068);
  and2 I030_147(w_030_147, w_029_511, w_001_716);
  and2 I030_150(w_030_150, w_003_039, w_027_470);
  or2  I030_154(w_030_154, w_029_1003, w_005_202);
  or2  I030_159(w_030_159, w_018_086, w_006_248);
  nand2 I030_161(w_030_161, w_017_1005, w_021_233);
  not1 I030_167(w_030_167, w_026_994);
  nand2 I030_169(w_030_169, w_004_1091, w_005_285);
  and2 I030_170(w_030_170, w_006_191, w_000_1634);
  or2  I030_172(w_030_172, w_008_705, w_013_233);
  nand2 I030_173(w_030_173, w_019_882, w_013_143);
  or2  I030_174(w_030_174, w_009_038, w_024_165);
  and2 I030_175(w_030_175, w_009_011, w_023_656);
  not1 I030_179(w_030_179, w_007_228);
  nand2 I030_181(w_030_181, w_012_517, w_023_882);
  nand2 I030_182(w_030_182, w_010_251, w_020_123);
  or2  I030_183(w_030_183, w_026_602, w_021_240);
  or2  I030_184(w_030_184, w_010_119, w_000_682);
  not1 I030_185(w_030_185, w_022_304);
  nand2 I030_186(w_030_186, w_021_194, w_010_355);
  or2  I030_191(w_030_191, w_001_198, w_024_1623);
  and2 I030_196(w_030_196, w_003_163, w_022_310);
  not1 I030_206(w_030_206, w_018_232);
  and2 I030_207(w_030_207, w_029_740, w_008_502);
  and2 I030_208(w_030_208, w_000_1143, w_002_334);
  not1 I030_214(w_030_214, w_019_083);
  not1 I030_218(w_030_218, w_011_465);
  or2  I030_220(w_030_220, w_023_1348, w_029_583);
  nand2 I030_222(w_030_222, w_018_273, w_011_779);
  not1 I030_224(w_030_224, w_025_267);
  or2  I030_225(w_030_225, w_025_1273, w_010_013);
  not1 I030_227(w_030_227, w_028_342);
  nand2 I030_228(w_030_228, w_007_646, w_021_195);
  or2  I030_229(w_030_229, w_010_146, w_017_1365);
  and2 I030_239(w_030_239, w_015_008, w_007_216);
  or2  I030_240(w_030_240, w_027_563, w_001_506);
  nand2 I030_245(w_030_245, w_006_119, w_011_193);
  and2 I030_248(w_030_248, w_004_307, w_000_756);
  or2  I030_250(w_030_250, w_011_553, w_016_034);
  and2 I030_253(w_030_253, w_021_256, w_001_104);
  or2  I030_261(w_030_261, w_003_258, w_018_026);
  or2  I030_262(w_030_262, w_029_613, w_000_1054);
  nand2 I030_264(w_030_264, w_027_543, w_027_397);
  or2  I030_266(w_030_266, w_006_265, w_010_109);
  and2 I030_273(w_030_273, w_022_075, w_016_037);
  nand2 I030_302(w_030_302, w_014_070, w_029_709);
  nand2 I030_305(w_030_305, w_008_040, w_010_085);
  not1 I030_306(w_030_306, w_020_117);
  not1 I030_309(w_030_309, w_002_177);
  and2 I030_313(w_030_313, w_006_193, w_006_313);
  or2  I030_314(w_030_314, w_007_132, w_009_069);
  or2  I030_315(w_030_315, w_012_240, w_005_1119);
  or2  I030_317(w_030_317, w_013_252, w_008_108);
  nand2 I030_318(w_030_318, w_003_181, w_020_527);
  nand2 I030_334(w_030_334, w_012_482, w_028_624);
  or2  I030_339(w_030_339, w_006_001, w_010_024);
  and2 I030_344(w_030_344, w_014_333, w_008_622);
  or2  I030_345(w_030_345, w_018_171, w_001_1428);
  or2  I030_348(w_030_348, w_014_641, w_001_088);
  nand2 I030_349(w_030_349, w_009_059, w_005_425);
  nand2 I030_354(w_030_354, w_008_250, w_000_1474);
  and2 I030_362(w_030_362, w_001_326, w_015_171);
  nand2 I030_364(w_030_364, w_014_181, w_024_1241);
  not1 I030_368(w_030_368, w_003_078);
  not1 I030_380(w_030_380, w_009_073);
  not1 I030_382(w_030_382, w_005_1336);
  and2 I030_385(w_030_385, w_022_213, w_021_083);
  or2  I030_392(w_030_392, w_009_023, w_002_178);
  and2 I030_396(w_030_396, w_029_892, w_015_252);
  or2  I030_411(w_030_411, w_010_411, w_027_370);
  and2 I030_412(w_030_412, w_008_573, w_012_387);
  not1 I030_422(w_030_422, w_006_043);
  nand2 I030_424(w_030_424, w_017_647, w_004_926);
  or2  I030_426(w_030_426, w_021_189, w_019_586);
  not1 I030_430(w_030_430, w_026_491);
  or2  I030_434(w_030_434, w_001_310, w_029_1193);
  and2 I030_435(w_030_435, w_018_025, w_000_127);
  nand2 I030_444(w_030_444, w_005_1119, w_009_090);
  or2  I030_447(w_030_447, w_010_262, w_028_160);
  nand2 I030_454(w_030_454, w_017_1226, w_029_626);
  and2 I030_459(w_030_459, w_014_636, w_001_213);
  and2 I030_467(w_030_467, w_018_097, w_010_036);
  and2 I030_470(w_030_470, w_025_1379, w_017_1857);
  nand2 I030_471(w_030_471, w_003_271, w_025_518);
  or2  I030_477(w_030_477, w_027_014, w_019_141);
  not1 I030_491(w_030_491, w_025_768);
  nand2 I030_496(w_030_496, w_004_1595, w_000_717);
  nand2 I030_502(w_030_502, w_017_1469, w_024_1269);
  not1 I030_503(w_030_503, w_013_252);
  and2 I030_504(w_030_504, w_024_736, w_016_036);
  and2 I030_523(w_030_523, w_005_1045, w_022_210);
  not1 I030_525(w_030_525, w_013_160);
  or2  I030_533(w_030_533, w_008_788, w_022_012);
  and2 I030_534(w_030_534, w_016_003, w_021_276);
  not1 I030_542(w_030_542, w_001_715);
  or2  I030_548(w_030_548, w_019_024, w_002_175);
  nand2 I030_549(w_030_549, w_004_890, w_005_1501);
  or2  I030_557(w_030_557, w_002_348, w_029_486);
  nand2 I030_559(w_030_559, w_002_094, w_024_1327);
  and2 I030_561(w_030_561, w_013_136, w_005_1233);
  or2  I030_565(w_030_565, w_025_911, w_014_459);
  nand2 I030_570(w_030_570, w_022_369, w_021_150);
  not1 I030_571(w_030_571, w_000_1227);
  and2 I030_572(w_030_572, w_018_068, w_005_731);
  and2 I030_578(w_030_578, w_028_541, w_028_098);
  nand2 I030_591(w_030_591, w_019_491, w_013_171);
  nand2 I030_592(w_030_592, w_028_253, w_008_370);
  not1 I030_613(w_030_613, w_013_092);
  not1 I030_614(w_030_614, w_004_1466);
  not1 I030_615(w_030_615, w_002_022);
  or2  I030_620(w_030_620, w_011_028, w_014_703);
  not1 I030_623(w_030_623, w_025_695);
  and2 I030_625(w_030_625, w_007_151, w_017_1654);
  not1 I030_626(w_030_626, w_006_021);
  and2 I030_630(w_030_630, w_005_139, w_028_124);
  and2 I030_633(w_030_633, w_010_191, w_004_1413);
  not1 I030_634(w_030_634, w_005_668);
  not1 I030_635(w_030_635, w_011_328);
  or2  I030_636(w_030_636, w_013_151, w_012_195);
  and2 I030_638(w_030_638, w_019_123, w_024_1164);
  not1 I030_641(w_030_641, w_015_008);
  and2 I030_648(w_030_648, w_004_1423, w_006_256);
  and2 I030_653(w_030_653, w_029_073, w_002_114);
  nand2 I030_658(w_030_658, w_015_262, w_022_163);
  and2 I030_663(w_030_663, w_009_046, w_018_269);
  nand2 I030_664(w_030_664, w_013_057, w_019_202);
  and2 I030_667(w_030_667, w_001_1115, w_021_115);
  nand2 I030_670(w_030_670, w_025_817, w_015_200);
  or2  I030_677(w_030_677, w_011_597, w_021_089);
  not1 I030_679(w_030_679, w_014_420);
  and2 I030_695(w_030_695, w_025_1543, w_019_1031);
  nand2 I030_696(w_030_696, w_011_210, w_009_006);
  nand2 I030_699(w_030_699, w_003_130, w_017_982);
  nand2 I030_705(w_030_705, w_018_069, w_020_993);
  or2  I030_706(w_030_706, w_007_351, w_021_140);
  not1 I030_710(w_030_710, w_015_241);
  and2 I030_715(w_030_715, w_011_804, w_006_232);
  not1 I030_716(w_030_716, w_010_193);
  nand2 I030_723(w_030_723, w_012_512, w_005_576);
  not1 I030_727(w_030_727, w_000_638);
  nand2 I030_732(w_030_732, w_024_840, w_004_1552);
  and2 I030_737(w_030_737, w_029_584, w_003_050);
  or2  I030_742(w_030_742, w_007_1579, w_016_033);
  or2  I030_745(w_030_745, w_024_263, w_005_1034);
  not1 I030_747(w_030_747, w_006_185);
  and2 I030_753(w_030_753, w_000_1361, w_022_356);
  not1 I030_757(w_030_757, w_023_829);
  nand2 I030_766(w_030_766, w_011_631, w_019_212);
  not1 I030_767(w_030_767, w_009_032);
  or2  I030_769(w_030_769, w_004_1807, w_004_260);
  or2  I030_774(w_030_774, w_022_137, w_000_688);
  and2 I030_776(w_030_776, w_027_069, w_006_169);
  and2 I030_777(w_030_777, w_024_195, w_013_109);
  or2  I030_780(w_030_780, w_013_267, w_010_193);
  and2 I030_781(w_030_781, w_026_1491, w_029_084);
  and2 I030_783(w_030_783, w_001_1374, w_024_1404);
  or2  I030_789(w_030_789, w_021_271, w_022_371);
  nand2 I030_795(w_030_795, w_015_237, w_025_1085);
  not1 I030_799(w_030_799, w_006_105);
  nand2 I030_804(w_030_804, w_004_1206, w_028_244);
  and2 I030_811(w_030_811, w_010_078, w_018_052);
  or2  I030_816(w_030_816, w_009_067, w_020_811);
  nand2 I030_826(w_030_826, w_024_524, w_014_118);
  or2  I030_830(w_030_830, w_021_054, w_011_112);
  and2 I030_837(w_030_837, w_004_012, w_006_340);
  or2  I030_840(w_030_840, w_013_013, w_024_047);
  nand2 I030_845(w_030_845, w_017_773, w_029_1337);
  and2 I030_852(w_030_852, w_029_014, w_011_293);
  or2  I031_003(w_031_003, w_024_153, w_019_1085);
  and2 I031_004(w_031_004, w_012_223, w_026_382);
  or2  I031_012(w_031_012, w_024_311, w_009_016);
  not1 I031_016(w_031_016, w_018_102);
  or2  I031_021(w_031_021, w_003_040, w_018_050);
  and2 I031_027(w_031_027, w_006_068, w_020_460);
  nand2 I031_037(w_031_037, w_002_015, w_015_196);
  not1 I031_038(w_031_038, w_028_714);
  and2 I031_039(w_031_039, w_025_1441, w_000_708);
  not1 I031_040(w_031_040, w_020_1125);
  nand2 I031_050(w_031_050, w_021_122, w_015_047);
  not1 I031_051(w_031_051, w_023_1225);
  nand2 I031_052(w_031_052, w_028_325, w_002_468);
  or2  I031_054(w_031_054, w_021_244, w_010_207);
  and2 I031_057(w_031_057, w_012_416, w_013_209);
  not1 I031_061(w_031_061, w_004_1202);
  or2  I031_062(w_031_062, w_022_009, w_004_639);
  and2 I031_076(w_031_076, w_026_545, w_000_1396);
  not1 I031_078(w_031_078, w_017_1195);
  and2 I031_087(w_031_087, w_013_012, w_005_1562);
  or2  I031_091(w_031_091, w_017_1626, w_023_1502);
  or2  I031_092(w_031_092, w_020_323, w_026_419);
  not1 I031_100(w_031_100, w_006_124);
  nand2 I031_102(w_031_102, w_005_1094, w_002_363);
  or2  I031_111(w_031_111, w_022_129, w_003_198);
  nand2 I031_113(w_031_113, w_030_380, w_004_723);
  or2  I031_116(w_031_116, w_019_482, w_013_103);
  or2  I031_117(w_031_117, w_001_092, w_011_642);
  nand2 I031_123(w_031_123, w_014_686, w_000_1790);
  and2 I031_134(w_031_134, w_014_795, w_005_080);
  nand2 I031_136(w_031_136, w_010_244, w_003_081);
  not1 I031_137(w_031_137, w_004_836);
  and2 I031_145(w_031_145, w_000_534, w_027_048);
  and2 I031_150(w_031_150, w_019_962, w_006_011);
  or2  I031_152(w_031_152, w_029_490, w_023_758);
  or2  I031_153(w_031_153, w_024_905, w_021_207);
  and2 I031_159(w_031_159, w_008_773, w_006_141);
  or2  I031_184(w_031_184, w_026_1359, w_003_191);
  or2  I031_194(w_031_194, w_023_1068, w_000_1440);
  and2 I031_201(w_031_201, w_024_355, w_017_1557);
  or2  I031_210(w_031_210, w_008_646, w_003_025);
  or2  I031_217(w_031_217, w_020_717, w_012_173);
  or2  I031_226(w_031_226, w_015_062, w_013_291);
  and2 I031_228(w_031_228, w_015_015, w_009_045);
  nand2 I031_229(w_031_229, w_002_189, w_024_043);
  not1 I031_246(w_031_246, w_007_784);
  or2  I031_248(w_031_248, w_002_015, w_008_813);
  or2  I031_250(w_031_250, w_000_1046, w_001_1612);
  not1 I031_252(w_031_252, w_008_336);
  or2  I031_256(w_031_256, w_002_568, w_013_174);
  or2  I031_260(w_031_260, w_023_864, w_024_899);
  nand2 I031_265(w_031_265, w_003_191, w_002_107);
  not1 I031_270(w_031_270, w_015_008);
  nand2 I031_274(w_031_274, w_024_1404, w_002_074);
  nand2 I031_279(w_031_279, w_018_148, w_011_417);
  and2 I031_284(w_031_284, w_014_256, w_003_149);
  or2  I031_287(w_031_287, w_020_905, w_027_097);
  not1 I031_289(w_031_289, w_000_1241);
  or2  I031_292(w_031_292, w_030_102, w_010_093);
  or2  I031_296(w_031_296, w_025_145, w_019_797);
  not1 I031_300(w_031_300, w_013_017);
  or2  I031_306(w_031_306, w_000_1615, w_011_749);
  nand2 I031_308(w_031_308, w_002_138, w_029_210);
  not1 I031_312(w_031_312, w_023_190);
  or2  I031_315(w_031_315, w_019_032, w_002_435);
  not1 I031_330(w_031_330, w_028_159);
  nand2 I031_333(w_031_333, w_019_202, w_011_433);
  or2  I031_337(w_031_337, w_029_377, w_005_070);
  and2 I031_340(w_031_340, w_012_193, w_025_014);
  or2  I031_341(w_031_341, w_025_1401, w_028_135);
  or2  I031_343(w_031_343, w_021_065, w_030_534);
  and2 I031_349(w_031_349, w_017_781, w_018_005);
  and2 I031_350(w_031_350, w_015_212, w_014_629);
  and2 I031_351(w_031_351, w_003_032, w_017_1575);
  or2  I031_356(w_031_356, w_006_231, w_007_1565);
  and2 I031_357(w_031_357, w_008_495, w_017_841);
  not1 I031_359(w_031_359, w_018_255);
  not1 I031_366(w_031_366, w_008_438);
  nand2 I031_370(w_031_370, w_025_1007, w_022_304);
  not1 I031_378(w_031_378, w_003_125);
  not1 I031_384(w_031_384, w_012_510);
  not1 I031_385(w_031_385, w_020_764);
  nand2 I031_387(w_031_387, w_013_089, w_005_1152);
  nand2 I031_389(w_031_389, w_002_226, w_026_751);
  and2 I031_394(w_031_394, w_017_1768, w_022_306);
  or2  I031_395(w_031_395, w_023_261, w_024_1010);
  or2  I031_398(w_031_398, w_030_710, w_008_799);
  or2  I031_404(w_031_404, w_014_437, w_020_493);
  not1 I031_409(w_031_409, w_004_562);
  not1 I031_422(w_031_422, w_002_444);
  or2  I031_425(w_031_425, w_012_252, w_016_011);
  or2  I031_429(w_031_429, w_027_236, w_007_907);
  or2  I031_449(w_031_449, w_020_007, w_002_429);
  or2  I031_456(w_031_456, w_002_183, w_012_573);
  and2 I031_457(w_031_457, w_010_321, w_008_743);
  not1 I031_465(w_031_465, w_012_364);
  or2  I031_468(w_031_468, w_013_307, w_000_1629);
  nand2 I031_476(w_031_476, w_022_376, w_020_1198);
  nand2 I031_480(w_031_480, w_006_303, w_015_125);
  and2 I031_485(w_031_485, w_007_816, w_029_211);
  nand2 I031_492(w_031_492, w_021_101, w_025_179);
  not1 I031_495(w_031_495, w_000_421);
  and2 I031_500(w_031_500, w_001_1561, w_002_374);
  nand2 I031_502(w_031_502, w_016_020, w_019_259);
  and2 I031_509(w_031_509, w_024_277, w_003_120);
  and2 I031_510(w_031_510, w_014_376, w_008_569);
  nand2 I031_511(w_031_511, w_008_656, w_009_064);
  nand2 I031_513(w_031_513, w_007_205, w_018_143);
  or2  I031_515(w_031_515, w_030_179, w_029_143);
  not1 I031_517(w_031_517, w_016_004);
  or2  I031_521(w_031_521, w_008_817, w_023_293);
  or2  I031_529(w_031_529, w_000_695, w_017_479);
  nand2 I031_536(w_031_536, w_027_130, w_001_054);
  or2  I031_546(w_031_546, w_016_024, w_012_581);
  nand2 I031_564(w_031_564, w_013_132, w_022_083);
  nand2 I031_575(w_031_575, w_010_381, w_022_340);
  or2  I031_576(w_031_576, w_019_507, w_010_150);
  not1 I031_587(w_031_587, w_004_179);
  nand2 I031_594(w_031_594, w_025_1120, w_006_149);
  nand2 I031_597(w_031_597, w_019_1097, w_025_1472);
  or2  I031_609(w_031_609, w_014_477, w_022_137);
  and2 I031_610(w_031_610, w_023_1336, w_026_1201);
  not1 I031_611(w_031_611, w_019_494);
  not1 I031_617(w_031_617, w_010_051);
  nand2 I031_619(w_031_619, w_026_884, w_008_544);
  and2 I031_620(w_031_620, w_026_439, w_006_070);
  not1 I031_625(w_031_625, w_030_020);
  not1 I031_631(w_031_631, w_030_776);
  nand2 I031_634(w_031_634, w_007_1279, w_003_262);
  nand2 I031_635(w_031_635, w_004_1458, w_015_246);
  and2 I031_643(w_031_643, w_011_817, w_019_898);
  or2  I031_645(w_031_645, w_020_490, w_010_371);
  and2 I031_647(w_031_647, w_028_581, w_006_101);
  not1 I031_658(w_031_658, w_030_447);
  and2 I031_662(w_031_662, w_003_110, w_025_416);
  nand2 I031_674(w_031_674, w_005_611, w_020_196);
  or2  I031_676(w_031_676, w_002_549, w_029_305);
  not1 I031_684(w_031_684, w_005_949);
  and2 I031_697(w_031_697, w_000_1018, w_021_058);
  nand2 I031_704(w_031_704, w_026_453, w_003_248);
  nand2 I031_712(w_031_712, w_004_008, w_016_024);
  and2 I031_713(w_031_713, w_003_194, w_014_242);
  nand2 I031_715(w_031_715, w_010_394, w_015_089);
  nand2 I031_718(w_031_718, w_003_038, w_011_365);
  or2  I031_724(w_031_724, w_021_025, w_001_113);
  nand2 I031_726(w_031_726, w_008_426, w_019_627);
  and2 I031_733(w_031_733, w_023_1580, w_029_586);
  not1 I031_743(w_031_743, w_023_282);
  and2 I031_744(w_031_744, w_022_244, w_023_219);
  not1 I031_750(w_031_750, w_018_178);
  not1 I031_752(w_031_752, w_020_905);
  nand2 I031_753(w_031_753, w_019_547, w_011_611);
  nand2 I031_762(w_031_762, w_008_317, w_027_110);
  or2  I031_766(w_031_766, w_010_245, w_007_964);
  and2 I031_770(w_031_770, w_022_321, w_017_1128);
  not1 I031_777(w_031_777, w_005_1075);
  or2  I031_778(w_031_778, w_015_275, w_013_234);
  nand2 I031_781(w_031_781, w_004_840, w_026_1116);
  or2  I031_786(w_031_786, w_024_071, w_020_766);
  or2  I031_789(w_031_789, w_003_018, w_016_032);
  and2 I031_814(w_031_814, w_028_630, w_012_133);
  or2  I031_815(w_031_815, w_013_280, w_000_235);
  not1 I031_819(w_031_819, w_004_1127);
  and2 I031_820(w_031_820, w_027_161, w_021_046);
  and2 I031_825(w_031_825, w_021_193, w_014_226);
  or2  I031_827(w_031_827, w_027_521, w_009_018);
  or2  I031_828(w_031_828, w_016_005, w_019_288);
  or2  I031_842(w_031_842, w_014_178, w_025_287);
  or2  I031_847(w_031_847, w_018_250, w_010_405);
  or2  I031_848(w_031_848, w_023_646, w_026_1027);
  nand2 I031_852(w_031_852, w_022_290, w_025_1655);
  nand2 I031_853(w_031_853, w_024_011, w_000_1712);
  not1 I031_861(w_031_861, w_017_1049);
  nand2 I031_864(w_031_864, w_013_150, w_019_675);
  or2  I031_874(w_031_874, w_022_374, w_027_242);
  and2 I031_917(w_031_917, w_004_1840, w_018_206);
  nand2 I031_925(w_031_925, w_004_1760, w_016_029);
  not1 I031_934(w_031_934, w_001_034);
  or2  I031_937(w_031_937, w_011_247, w_000_1870);
  or2  I031_949(w_031_949, w_000_1231, w_022_265);
  or2  I031_963(w_031_963, w_025_008, w_020_1030);
  not1 I031_974(w_031_974, w_003_074);
  nand2 I031_981(w_031_981, w_002_109, w_017_1325);
  or2  I031_983(w_031_983, w_021_269, w_005_1304);
  not1 I031_985(w_031_985, w_029_1005);
  and2 I031_988(w_031_988, w_019_526, w_015_105);
  or2  I031_990(w_031_990, w_010_082, w_013_043);
  or2  I031_1001(w_031_1001, w_001_535, w_020_191);
  and2 I031_1006(w_031_1006, w_011_881, w_014_065);
  and2 I031_1019(w_031_1019, w_001_761, w_000_1460);
  nand2 I031_1021(w_031_1021, w_029_1296, w_013_024);
  or2  I031_1025(w_031_1025, w_003_114, w_013_070);
  nand2 I031_1026(w_031_1026, w_012_563, w_030_777);
  not1 I031_1027(w_031_1027, w_023_294);
  and2 I031_1037(w_031_1037, w_003_040, w_017_1071);
  not1 I031_1045(w_031_1045, w_027_516);
  not1 I031_1052(w_031_1052, w_000_1734);
  or2  I031_1054(w_031_1054, w_002_096, w_001_565);
  or2  I031_1065(w_031_1065, w_025_1357, w_008_706);
  and2 I031_1109(w_031_1109, w_009_009, w_001_1482);
  or2  I031_1110(w_031_1110, w_007_434, w_024_120);
  and2 I031_1126(w_031_1126, w_004_1696, w_018_011);
  nand2 I031_1129(w_031_1129, w_020_289, w_002_150);
  nand2 I031_1130(w_031_1130, w_016_019, w_019_834);
  or2  I032_000(w_032_000, w_005_307, w_004_981);
  not1 I032_001(w_032_001, w_012_250);
  nand2 I032_002(w_032_002, w_024_1473, w_006_322);
  and2 I032_003(w_032_003, w_027_061, w_009_077);
  and2 I032_004(w_032_004, w_031_340, w_011_151);
  nand2 I032_005(w_032_005, w_030_184, w_004_1188);
  not1 I032_009(w_032_009, w_009_091);
  and2 I032_011(w_032_011, w_003_152, w_007_1281);
  and2 I032_012(w_032_012, w_011_469, w_006_195);
  nand2 I032_013(w_032_013, w_008_269, w_015_173);
  not1 I032_015(w_032_015, w_002_205);
  not1 I032_018(w_032_018, w_003_071);
  or2  I032_019(w_032_019, w_005_1035, w_028_106);
  or2  I032_020(w_032_020, w_023_1502, w_026_119);
  or2  I032_021(w_032_021, w_009_016, w_003_188);
  nand2 I032_023(w_032_023, w_018_048, w_015_041);
  and2 I032_025(w_032_025, w_019_423, w_025_1544);
  and2 I032_026(w_032_026, w_021_002, w_001_1037);
  and2 I032_027(w_032_027, w_027_564, w_014_149);
  and2 I032_028(w_032_028, w_017_1633, w_025_1028);
  and2 I032_029(w_032_029, w_000_1206, w_020_519);
  not1 I032_030(w_032_030, w_003_161);
  and2 I032_031(w_032_031, w_019_014, w_024_084);
  nand2 I032_032(w_032_032, w_017_1630, w_019_090);
  not1 I032_035(w_032_035, w_021_255);
  nand2 I032_036(w_032_036, w_021_091, w_007_1495);
  not1 I032_037(w_032_037, w_010_328);
  not1 I032_038(w_032_038, w_029_694);
  nand2 I032_039(w_032_039, w_003_265, w_024_785);
  nand2 I032_042(w_032_042, w_018_129, w_012_503);
  nand2 I032_043(w_032_043, w_001_947, w_022_385);
  nand2 I032_045(w_032_045, w_022_388, w_000_1071);
  nand2 I032_046(w_032_046, w_029_476, w_005_974);
  or2  I032_048(w_032_048, w_026_741, w_021_053);
  nand2 I032_050(w_032_050, w_007_1355, w_008_712);
  and2 I032_051(w_032_051, w_024_823, w_019_081);
  or2  I032_052(w_032_052, w_019_253, w_012_052);
  and2 I032_053(w_032_053, w_018_046, w_014_266);
  or2  I032_054(w_032_054, w_011_645, w_018_080);
  not1 I032_056(w_032_056, w_005_1109);
  not1 I032_057(w_032_057, w_012_464);
  not1 I032_058(w_032_058, w_021_212);
  not1 I032_059(w_032_059, w_028_735);
  nand2 I032_061(w_032_061, w_006_035, w_002_176);
  nand2 I032_065(w_032_065, w_009_039, w_024_800);
  and2 I032_066(w_032_066, w_004_014, w_024_274);
  nand2 I032_067(w_032_067, w_029_1207, w_006_135);
  not1 I032_068(w_032_068, w_012_554);
  and2 I032_069(w_032_069, w_001_064, w_012_469);
  not1 I032_072(w_032_072, w_003_093);
  nand2 I032_073(w_032_073, w_008_748, w_027_572);
  or2  I032_075(w_032_075, w_010_123, w_026_1035);
  or2  I032_077(w_032_077, w_007_368, w_017_875);
  not1 I032_080(w_032_080, w_028_855);
  or2  I032_081(w_032_081, w_021_245, w_023_733);
  or2  I032_084(w_032_084, w_009_069, w_024_1089);
  or2  I032_086(w_032_086, w_020_385, w_022_344);
  nand2 I032_087(w_032_087, w_018_079, w_029_583);
  nand2 I032_089(w_032_089, w_013_209, w_030_126);
  or2  I032_090(w_032_090, w_015_057, w_030_227);
  and2 I032_091(w_032_091, w_021_126, w_004_1401);
  or2  I032_092(w_032_092, w_025_1406, w_007_543);
  and2 I032_095(w_032_095, w_008_480, w_017_102);
  not1 I032_098(w_032_098, w_029_088);
  nand2 I032_099(w_032_099, w_023_1494, w_002_274);
  and2 I032_101(w_032_101, w_003_016, w_029_1142);
  and2 I032_102(w_032_102, w_005_300, w_018_245);
  or2  I032_103(w_032_103, w_028_435, w_007_1365);
  and2 I032_105(w_032_105, w_013_253, w_018_016);
  nand2 I032_106(w_032_106, w_019_560, w_003_080);
  not1 I032_108(w_032_108, w_002_468);
  not1 I032_111(w_032_111, w_015_110);
  not1 I032_112(w_032_112, w_028_277);
  not1 I032_116(w_032_116, w_018_165);
  not1 I032_118(w_032_118, w_008_578);
  or2  I032_119(w_032_119, w_024_121, w_009_093);
  nand2 I032_122(w_032_122, w_002_461, w_021_077);
  and2 I032_126(w_032_126, w_023_1313, w_001_1629);
  not1 I032_127(w_032_127, w_029_538);
  nand2 I032_130(w_032_130, w_013_304, w_027_175);
  not1 I032_131(w_032_131, w_006_193);
  not1 I032_132(w_032_132, w_010_413);
  not1 I032_134(w_032_134, w_017_950);
  nand2 I032_135(w_032_135, w_018_082, w_021_263);
  and2 I032_138(w_032_138, w_029_692, w_023_319);
  or2  I032_140(w_032_140, w_027_215, w_022_428);
  or2  I032_141(w_032_141, w_008_609, w_020_431);
  and2 I032_142(w_032_142, w_010_171, w_004_399);
  or2  I032_144(w_032_144, w_016_003, w_022_146);
  or2  I032_146(w_032_146, w_003_183, w_002_391);
  and2 I032_147(w_032_147, w_029_976, w_019_347);
  not1 I032_148(w_032_148, w_027_409);
  and2 I032_150(w_032_150, w_031_658, w_012_093);
  or2  I032_152(w_032_152, w_007_934, w_021_120);
  nand2 I032_153(w_032_153, w_024_201, w_002_063);
  and2 I032_154(w_032_154, w_031_502, w_027_279);
  and2 I032_155(w_032_155, w_022_249, w_018_063);
  not1 I032_156(w_032_156, w_015_169);
  nand2 I032_158(w_032_158, w_011_677, w_020_503);
  not1 I032_160(w_032_160, w_017_947);
  nand2 I032_163(w_032_163, w_006_310, w_022_033);
  not1 I032_164(w_032_164, w_017_1530);
  and2 I032_165(w_032_165, w_023_013, w_015_084);
  nand2 I032_167(w_032_167, w_011_374, w_016_035);
  and2 I032_169(w_032_169, w_004_881, w_016_003);
  nand2 I032_170(w_032_170, w_006_284, w_030_264);
  nand2 I032_173(w_032_173, w_014_492, w_030_134);
  nand2 I032_175(w_032_175, w_015_128, w_020_1095);
  and2 I032_176(w_032_176, w_025_328, w_004_1028);
  or2  I032_179(w_032_179, w_031_777, w_001_1645);
  or2  I032_180(w_032_180, w_031_715, w_023_348);
  and2 I032_182(w_032_182, w_000_1040, w_029_165);
  and2 I032_185(w_032_185, w_006_109, w_017_1271);
  not1 I032_187(w_032_187, w_026_949);
  not1 I032_190(w_032_190, w_003_035);
  or2  I032_193(w_032_193, w_003_298, w_002_084);
  or2  I032_194(w_032_194, w_021_169, w_008_574);
  or2  I032_195(w_032_195, w_029_583, w_013_223);
  nand2 I032_196(w_032_196, w_001_982, w_021_276);
  or2  I032_197(w_032_197, w_001_188, w_026_108);
  not1 I032_199(w_032_199, w_029_911);
  not1 I032_201(w_032_201, w_002_319);
  nand2 I032_202(w_032_202, w_000_1436, w_025_287);
  not1 I032_206(w_032_206, w_026_1240);
  not1 I032_208(w_032_208, w_019_778);
  and2 I032_210(w_032_210, w_028_097, w_006_074);
  nand2 I032_211(w_032_211, w_004_1089, w_001_1567);
  not1 I032_212(w_032_212, w_016_032);
  or2  I032_215(w_032_215, w_025_111, w_020_342);
  or2  I032_216(w_032_216, w_010_223, w_022_392);
  nand2 I032_218(w_032_218, w_010_417, w_029_039);
  not1 I032_222(w_032_222, w_006_170);
  and2 I032_223(w_032_223, w_016_028, w_006_182);
  not1 I032_224(w_032_224, w_025_221);
  and2 I032_225(w_032_225, w_014_437, w_007_1284);
  nand2 I032_227(w_032_227, w_027_013, w_006_322);
  or2  I032_231(w_032_231, w_001_1409, w_030_523);
  not1 I032_232(w_032_232, w_013_293);
  or2  I032_233(w_032_233, w_017_899, w_021_026);
  nand2 I032_234(w_032_234, w_017_595, w_009_027);
  nand2 I032_235(w_032_235, w_007_1478, w_012_271);
  nand2 I032_236(w_032_236, w_030_025, w_022_084);
  and2 I032_237(w_032_237, w_025_1629, w_001_1515);
  nand2 I032_239(w_032_239, w_002_060, w_011_835);
  nand2 I032_241(w_032_241, w_018_195, w_025_206);
  nand2 I032_244(w_032_244, w_011_243, w_013_044);
  or2  I033_001(w_033_001, w_030_634, w_014_309);
  not1 I033_004(w_033_004, w_014_313);
  and2 I033_012(w_033_012, w_018_066, w_030_571);
  and2 I033_016(w_033_016, w_021_063, w_010_238);
  not1 I033_018(w_033_018, w_006_095);
  not1 I033_022(w_033_022, w_017_1505);
  not1 I033_033(w_033_033, w_008_689);
  not1 I033_040(w_033_040, w_002_203);
  and2 I033_053(w_033_053, w_020_717, w_004_075);
  or2  I033_055(w_033_055, w_013_249, w_024_1431);
  and2 I033_058(w_033_058, w_023_300, w_010_021);
  and2 I033_064(w_033_064, w_013_135, w_007_238);
  nand2 I033_067(w_033_067, w_003_234, w_006_288);
  and2 I033_069(w_033_069, w_014_335, w_026_153);
  or2  I033_081(w_033_081, w_013_117, w_022_225);
  and2 I033_082(w_033_082, w_000_761, w_010_374);
  not1 I033_083(w_033_083, w_023_097);
  or2  I033_086(w_033_086, w_012_662, w_003_202);
  and2 I033_087(w_033_087, w_028_764, w_012_101);
  nand2 I033_090(w_033_090, w_023_180, w_023_527);
  nand2 I033_093(w_033_093, w_004_283, w_015_289);
  or2  I033_099(w_033_099, w_028_491, w_010_286);
  and2 I033_103(w_033_103, w_006_106, w_026_1448);
  nand2 I033_107(w_033_107, w_026_027, w_003_144);
  or2  I033_109(w_033_109, w_025_1476, w_002_489);
  not1 I033_112(w_033_112, w_003_173);
  not1 I033_113(w_033_113, w_004_167);
  or2  I033_114(w_033_114, w_030_072, w_001_1036);
  nand2 I033_115(w_033_115, w_022_235, w_031_1045);
  not1 I033_117(w_033_117, w_006_078);
  and2 I033_121(w_033_121, w_028_549, w_030_430);
  nand2 I033_123(w_033_123, w_007_1353, w_003_140);
  not1 I033_127(w_033_127, w_005_1494);
  and2 I033_137(w_033_137, w_020_456, w_026_1427);
  or2  I033_138(w_033_138, w_027_394, w_018_059);
  or2  I033_139(w_033_139, w_005_319, w_028_145);
  or2  I033_168(w_033_168, w_031_384, w_027_362);
  or2  I033_175(w_033_175, w_010_203, w_012_523);
  not1 I033_191(w_033_191, w_032_167);
  nand2 I033_195(w_033_195, w_015_140, w_008_222);
  and2 I033_210(w_033_210, w_027_082, w_031_265);
  and2 I033_218(w_033_218, w_014_288, w_019_040);
  nand2 I033_221(w_033_221, w_011_394, w_003_243);
  and2 I033_222(w_033_222, w_022_013, w_010_276);
  nand2 I033_232(w_033_232, w_026_572, w_028_146);
  not1 I033_234(w_033_234, w_025_596);
  or2  I033_244(w_033_244, w_007_208, w_008_819);
  or2  I033_245(w_033_245, w_024_964, w_015_140);
  not1 I033_248(w_033_248, w_010_316);
  not1 I033_249(w_033_249, w_003_156);
  not1 I033_260(w_033_260, w_007_214);
  or2  I033_276(w_033_276, w_003_311, w_030_679);
  nand2 I033_283(w_033_283, w_009_058, w_011_424);
  nand2 I033_284(w_033_284, w_024_1327, w_024_616);
  nand2 I033_294(w_033_294, w_007_358, w_028_678);
  not1 I033_307(w_033_307, w_020_924);
  not1 I033_314(w_033_314, w_000_825);
  nand2 I033_320(w_033_320, w_005_809, w_015_226);
  not1 I033_322(w_033_322, w_018_280);
  and2 I033_323(w_033_323, w_026_1008, w_021_027);
  nand2 I033_326(w_033_326, w_001_371, w_007_021);
  nand2 I033_332(w_033_332, w_024_168, w_000_1809);
  and2 I033_341(w_033_341, w_013_286, w_016_024);
  nand2 I033_347(w_033_347, w_029_387, w_012_270);
  not1 I033_355(w_033_355, w_025_232);
  nand2 I033_361(w_033_361, w_027_052, w_014_101);
  or2  I033_370(w_033_370, w_012_336, w_030_504);
  nand2 I033_373(w_033_373, w_022_078, w_022_386);
  nand2 I033_390(w_033_390, w_018_070, w_004_1011);
  nand2 I033_391(w_033_391, w_029_391, w_032_126);
  nand2 I033_393(w_033_393, w_017_917, w_008_017);
  not1 I033_397(w_033_397, w_014_022);
  and2 I033_413(w_033_413, w_001_1655, w_017_457);
  and2 I033_423(w_033_423, w_002_488, w_013_289);
  nand2 I033_453(w_033_453, w_006_189, w_000_1058);
  or2  I033_457(w_033_457, w_011_816, w_015_071);
  not1 I033_476(w_033_476, w_017_616);
  nand2 I033_478(w_033_478, w_020_991, w_010_013);
  and2 I033_482(w_033_482, w_016_017, w_014_181);
  or2  I033_485(w_033_485, w_017_1407, w_023_1594);
  not1 I033_498(w_033_498, w_025_712);
  and2 I033_501(w_033_501, w_016_007, w_028_256);
  or2  I033_523(w_033_523, w_022_182, w_024_1094);
  or2  I033_528(w_033_528, w_006_191, w_029_308);
  and2 I033_539(w_033_539, w_025_035, w_004_251);
  not1 I033_550(w_033_550, w_019_024);
  or2  I033_563(w_033_563, w_031_027, w_016_019);
  or2  I033_574(w_033_574, w_018_070, w_014_504);
  or2  I033_595(w_033_595, w_000_663, w_015_060);
  nand2 I033_600(w_033_600, w_031_536, w_017_1116);
  not1 I033_602(w_033_602, w_012_550);
  and2 I033_605(w_033_605, w_011_674, w_011_128);
  not1 I033_629(w_033_629, w_015_074);
  or2  I033_631(w_033_631, w_032_210, w_012_666);
  or2  I033_634(w_033_634, w_023_1019, w_010_020);
  not1 I033_638(w_033_638, w_020_1060);
  not1 I033_643(w_033_643, w_008_639);
  nand2 I033_649(w_033_649, w_001_915, w_008_293);
  not1 I033_655(w_033_655, w_001_517);
  nand2 I033_660(w_033_660, w_004_724, w_013_240);
  not1 I033_672(w_033_672, w_026_1006);
  and2 I033_682(w_033_682, w_007_203, w_021_251);
  and2 I033_697(w_033_697, w_016_018, w_011_022);
  or2  I033_708(w_033_708, w_002_121, w_029_206);
  nand2 I033_713(w_033_713, w_012_405, w_022_178);
  not1 I033_722(w_033_722, w_025_1192);
  nand2 I033_730(w_033_730, w_001_1538, w_010_347);
  nand2 I033_752(w_033_752, w_021_228, w_020_667);
  or2  I033_755(w_033_755, w_012_255, w_006_066);
  or2  I033_801(w_033_801, w_009_050, w_022_230);
  and2 I033_803(w_033_803, w_005_523, w_032_092);
  and2 I033_805(w_033_805, w_019_757, w_014_768);
  or2  I033_845(w_033_845, w_010_017, w_015_210);
  or2  I033_847(w_033_847, w_031_062, w_009_025);
  or2  I033_869(w_033_869, w_032_098, w_021_033);
  and2 I033_876(w_033_876, w_002_559, w_001_981);
  not1 I033_895(w_033_895, w_021_063);
  and2 I033_923(w_033_923, w_019_571, w_000_1852);
  nand2 I033_927(w_033_927, w_013_327, w_027_403);
  and2 I033_944(w_033_944, w_004_235, w_011_725);
  nand2 I033_949(w_033_949, w_027_530, w_001_1536);
  nand2 I033_970(w_033_970, w_016_020, w_031_617);
  not1 I033_979(w_033_979, w_012_388);
  not1 I033_987(w_033_987, w_017_1006);
  not1 I033_999(w_033_999, w_019_130);
  and2 I033_1001(w_033_1001, w_000_243, w_012_159);
  or2  I033_1015(w_033_1015, w_022_354, w_015_282);
  and2 I033_1018(w_033_1018, w_030_228, w_025_314);
  and2 I033_1032(w_033_1032, w_024_488, w_005_1448);
  not1 I033_1033(w_033_1033, w_013_086);
  or2  I033_1044(w_033_1044, w_014_102, w_025_342);
  and2 I033_1049(w_033_1049, w_029_471, w_008_143);
  not1 I033_1060(w_033_1060, w_013_044);
  not1 I033_1068(w_033_1068, w_002_176);
  and2 I033_1076(w_033_1076, w_000_1082, w_010_225);
  not1 I033_1077(w_033_1077, w_016_019);
  and2 I033_1098(w_033_1098, w_015_189, w_023_1460);
  not1 I033_1099(w_033_1099, w_008_714);
  not1 I033_1104(w_033_1104, w_014_443);
  and2 I033_1112(w_033_1112, w_031_284, w_023_135);
  or2  I033_1116(w_033_1116, w_004_1107, w_009_008);
  or2  I033_1136(w_033_1136, w_024_1568, w_011_001);
  and2 I033_1142(w_033_1142, w_028_823, w_000_467);
  not1 I033_1156(w_033_1156, w_022_101);
  and2 I033_1187(w_033_1187, w_032_020, w_028_852);
  and2 I033_1193(w_033_1193, w_009_031, w_026_159);
  and2 I033_1205(w_033_1205, w_023_447, w_031_037);
  or2  I033_1210(w_033_1210, w_009_006, w_030_816);
  not1 I033_1214(w_033_1214, w_001_1333);
  or2  I033_1235(w_033_1235, w_004_737, w_020_064);
  or2  I033_1239(w_033_1239, w_016_019, w_015_140);
  and2 I033_1243(w_033_1243, w_001_266, w_031_252);
  or2  I033_1249(w_033_1249, w_010_124, w_011_583);
  and2 I033_1268(w_033_1268, w_012_111, w_030_175);
  nand2 I033_1277(w_033_1277, w_016_020, w_002_587);
  nand2 I033_1280(w_033_1280, w_027_178, w_008_748);
  nand2 I033_1284(w_033_1284, w_029_051, w_012_587);
  nand2 I033_1291(w_033_1291, w_027_215, w_032_095);
  not1 I033_1295(w_033_1295, w_003_312);
  and2 I033_1305(w_033_1305, w_007_1497, w_031_1130);
  not1 I033_1307(w_033_1307, w_006_310);
  nand2 I033_1318(w_033_1318, w_026_1111, w_031_076);
  nand2 I033_1324(w_033_1324, w_032_077, w_017_1381);
  not1 I033_1357(w_033_1357, w_015_033);
  and2 I033_1375(w_033_1375, w_000_1114, w_024_222);
  nand2 I033_1376(w_033_1376, w_015_176, w_003_004);
  nand2 I033_1405(w_033_1405, w_014_341, w_021_088);
  or2  I033_1406(w_033_1406, w_008_550, w_028_028);
  or2  I033_1409(w_033_1409, w_012_650, w_024_683);
  nand2 I033_1411(w_033_1411, w_018_118, w_024_163);
  or2  I033_1417(w_033_1417, w_007_786, w_029_1053);
  not1 I033_1421(w_033_1421, w_030_658);
  nand2 I033_1429(w_033_1429, w_016_006, w_024_126);
  not1 I033_1436(w_033_1436, w_007_1554);
  and2 I033_1438(w_033_1438, w_014_787, w_019_547);
  not1 I033_1444(w_033_1444, w_030_245);
  or2  I033_1448(w_033_1448, w_030_578, w_010_102);
  and2 I033_1461(w_033_1461, w_022_342, w_029_1272);
  and2 I033_1489(w_033_1489, w_024_062, w_024_194);
  nand2 I033_1498(w_033_1498, w_031_529, w_015_006);
  and2 I033_1507(w_033_1507, w_001_822, w_002_495);
  not1 I033_1512(w_033_1512, w_002_537);
  nand2 I033_1523(w_033_1523, w_020_1258, w_032_127);
  and2 I033_1524(w_033_1524, w_030_667, w_028_565);
  nand2 I033_1551(w_033_1551, w_028_809, w_024_055);
  nand2 I033_1577(w_033_1577, w_031_990, w_030_477);
  and2 I033_1605(w_033_1605, w_016_035, w_030_070);
  not1 I033_1619(w_033_1619, w_002_086);
  and2 I033_1624(w_033_1624, w_008_836, w_013_085);
  and2 I033_1634(w_033_1634, w_015_189, w_001_156);
  or2  I033_1635(w_033_1635, w_023_301, w_025_877);
  and2 I033_1638(w_033_1638, w_025_1125, w_013_027);
  not1 I033_1643(w_033_1643, w_029_579);
  nand2 I033_1647(w_033_1647, w_011_872, w_031_949);
  nand2 I033_1650(w_033_1650, w_024_677, w_007_1594);
  or2  I034_006(w_034_006, w_023_1266, w_027_529);
  nand2 I034_007(w_034_007, w_002_336, w_029_632);
  and2 I034_009(w_034_009, w_029_416, w_021_092);
  nand2 I034_011(w_034_011, w_010_359, w_030_459);
  and2 I034_016(w_034_016, w_025_683, w_031_825);
  and2 I034_022(w_034_022, w_019_666, w_008_705);
  nand2 I034_031(w_034_031, w_008_743, w_004_322);
  or2  I034_034(w_034_034, w_025_1037, w_009_060);
  nand2 I034_044(w_034_044, w_001_947, w_024_059);
  and2 I034_057(w_034_057, w_003_243, w_022_070);
  or2  I034_061(w_034_061, w_015_229, w_012_101);
  or2  I034_066(w_034_066, w_001_149, w_008_418);
  nand2 I034_067(w_034_067, w_017_549, w_018_213);
  not1 I034_072(w_034_072, w_021_065);
  not1 I034_074(w_034_074, w_020_1121);
  and2 I034_079(w_034_079, w_020_643, w_003_207);
  nand2 I034_083(w_034_083, w_015_153, w_019_926);
  or2  I034_089(w_034_089, w_007_1412, w_017_1531);
  nand2 I034_090(w_034_090, w_032_018, w_012_323);
  or2  I034_099(w_034_099, w_033_1421, w_005_793);
  not1 I034_104(w_034_104, w_010_272);
  and2 I034_109(w_034_109, w_027_158, w_017_1852);
  and2 I034_114(w_034_114, w_013_194, w_025_1124);
  not1 I034_115(w_034_115, w_005_1370);
  and2 I034_116(w_034_116, w_030_716, w_030_183);
  and2 I034_121(w_034_121, w_006_262, w_008_087);
  and2 I034_122(w_034_122, w_026_1043, w_010_014);
  or2  I034_125(w_034_125, w_001_998, w_001_765);
  nand2 I034_130(w_034_130, w_000_1636, w_016_016);
  or2  I034_133(w_034_133, w_016_035, w_022_383);
  not1 I034_134(w_034_134, w_030_852);
  nand2 I034_140(w_034_140, w_005_256, w_033_1551);
  and2 I034_144(w_034_144, w_009_110, w_031_718);
  or2  I034_145(w_034_145, w_033_501, w_000_366);
  and2 I034_161(w_034_161, w_007_279, w_007_289);
  not1 I034_166(w_034_166, w_024_887);
  or2  I034_178(w_034_178, w_022_179, w_013_235);
  nand2 I034_182(w_034_182, w_012_284, w_021_060);
  or2  I034_185(w_034_185, w_019_580, w_019_900);
  or2  I034_189(w_034_189, w_021_234, w_013_048);
  nand2 I034_196(w_034_196, w_003_079, w_005_734);
  not1 I034_199(w_034_199, w_016_020);
  nand2 I034_201(w_034_201, w_008_721, w_004_738);
  nand2 I034_203(w_034_203, w_026_300, w_023_1503);
  and2 I034_204(w_034_204, w_014_110, w_013_289);
  and2 I034_205(w_034_205, w_014_104, w_029_166);
  nand2 I034_213(w_034_213, w_006_197, w_030_012);
  or2  I034_214(w_034_214, w_022_143, w_024_120);
  and2 I034_216(w_034_216, w_025_1249, w_000_1514);
  or2  I034_225(w_034_225, w_026_268, w_023_076);
  or2  I034_226(w_034_226, w_003_193, w_010_070);
  and2 I034_227(w_034_227, w_033_234, w_007_068);
  or2  I034_241(w_034_241, w_012_238, w_000_1917);
  nand2 I034_245(w_034_245, w_030_206, w_005_148);
  nand2 I034_248(w_034_248, w_017_1895, w_017_1129);
  nand2 I034_252(w_034_252, w_026_1158, w_013_170);
  and2 I034_254(w_034_254, w_004_1187, w_027_419);
  not1 I034_268(w_034_268, w_009_059);
  or2  I034_269(w_034_269, w_013_177, w_032_215);
  or2  I034_273(w_034_273, w_024_1226, w_027_383);
  and2 I034_274(w_034_274, w_010_285, w_017_1354);
  or2  I034_276(w_034_276, w_009_020, w_006_098);
  and2 I034_281(w_034_281, w_022_186, w_001_1670);
  nand2 I034_289(w_034_289, w_028_623, w_028_169);
  not1 I034_292(w_034_292, w_024_723);
  or2  I034_297(w_034_297, w_028_007, w_018_141);
  and2 I034_300(w_034_300, w_015_287, w_009_004);
  or2  I034_305(w_034_305, w_025_358, w_012_083);
  and2 I034_308(w_034_308, w_000_316, w_004_1664);
  or2  I034_309(w_034_309, w_010_205, w_019_344);
  not1 I034_314(w_034_314, w_005_257);
  not1 I034_315(w_034_315, w_033_137);
  nand2 I034_316(w_034_316, w_006_093, w_025_307);
  or2  I034_322(w_034_322, w_029_414, w_018_049);
  or2  I034_323(w_034_323, w_009_054, w_030_110);
  nand2 I034_328(w_034_328, w_031_040, w_010_305);
  and2 I034_329(w_034_329, w_028_404, w_004_059);
  nand2 I034_330(w_034_330, w_008_515, w_016_014);
  nand2 I034_336(w_034_336, w_007_018, w_031_315);
  or2  I034_339(w_034_339, w_026_909, w_009_104);
  nand2 I034_345(w_034_345, w_033_523, w_016_015);
  or2  I034_347(w_034_347, w_006_170, w_028_257);
  not1 I034_350(w_034_350, w_017_914);
  or2  I034_351(w_034_351, w_031_743, w_008_240);
  not1 I034_354(w_034_354, w_017_1809);
  nand2 I034_358(w_034_358, w_000_1813, w_028_418);
  nand2 I034_363(w_034_363, w_020_250, w_006_074);
  and2 I034_368(w_034_368, w_030_559, w_023_1421);
  nand2 I034_369(w_034_369, w_001_1093, w_006_191);
  nand2 I034_371(w_034_371, w_012_535, w_003_107);
  not1 I034_372(w_034_372, w_017_155);
  nand2 I034_376(w_034_376, w_019_627, w_028_120);
  not1 I034_377(w_034_377, w_016_038);
  or2  I034_378(w_034_378, w_032_185, w_001_769);
  not1 I034_379(w_034_379, w_020_465);
  nand2 I034_382(w_034_382, w_008_266, w_029_210);
  and2 I034_391(w_034_391, w_015_212, w_001_1508);
  and2 I034_398(w_034_398, w_009_040, w_033_755);
  and2 I034_400(w_034_400, w_018_141, w_001_1132);
  and2 I034_403(w_034_403, w_008_433, w_020_1097);
  not1 I034_404(w_034_404, w_014_169);
  not1 I034_405(w_034_405, w_023_1569);
  or2  I034_406(w_034_406, w_018_242, w_001_1037);
  nand2 I034_407(w_034_407, w_020_256, w_029_274);
  or2  I034_410(w_034_410, w_000_192, w_011_405);
  and2 I034_412(w_034_412, w_022_057, w_002_218);
  or2  I034_415(w_034_415, w_033_390, w_010_264);
  or2  I034_416(w_034_416, w_032_223, w_017_334);
  or2  I034_418(w_034_418, w_002_020, w_000_1118);
  and2 I034_419(w_034_419, w_010_073, w_002_367);
  and2 I034_420(w_034_420, w_010_367, w_008_771);
  and2 I034_422(w_034_422, w_010_054, w_007_348);
  and2 I034_424(w_034_424, w_018_254, w_028_237);
  not1 I034_430(w_034_430, w_021_270);
  not1 I034_433(w_034_433, w_028_655);
  or2  I034_434(w_034_434, w_005_1139, w_012_581);
  and2 I034_439(w_034_439, w_032_043, w_004_1805);
  or2  I034_441(w_034_441, w_028_690, w_033_1284);
  and2 I034_442(w_034_442, w_000_1138, w_033_1060);
  and2 I034_452(w_034_452, w_029_766, w_011_098);
  or2  I034_459(w_034_459, w_029_1106, w_008_019);
  nand2 I034_460(w_034_460, w_033_1076, w_023_181);
  nand2 I034_462(w_034_462, w_016_024, w_004_1115);
  and2 I034_463(w_034_463, w_011_058, w_033_1156);
  nand2 I034_471(w_034_471, w_015_196, w_018_057);
  not1 I034_475(w_034_475, w_027_183);
  not1 I034_476(w_034_476, w_031_137);
  not1 I034_486(w_034_486, w_027_345);
  nand2 I034_488(w_034_488, w_011_838, w_022_133);
  nand2 I034_494(w_034_494, w_009_107, w_002_209);
  nand2 I034_498(w_034_498, w_029_202, w_032_126);
  and2 I034_500(w_034_500, w_002_277, w_029_650);
  or2  I034_504(w_034_504, w_013_025, w_032_235);
  not1 I034_506(w_034_506, w_025_1483);
  or2  I034_511(w_034_511, w_000_1654, w_024_009);
  and2 I034_513(w_034_513, w_028_077, w_015_277);
  or2  I034_521(w_034_521, w_002_342, w_014_534);
  or2  I034_526(w_034_526, w_029_004, w_008_624);
  nand2 I034_527(w_034_527, w_027_093, w_026_991);
  and2 I034_528(w_034_528, w_006_157, w_023_996);
  or2  I034_545(w_034_545, w_022_094, w_018_212);
  or2  I034_551(w_034_551, w_019_962, w_012_036);
  and2 I034_555(w_034_555, w_007_892, w_032_065);
  nand2 I034_557(w_034_557, w_028_698, w_019_229);
  nand2 I034_558(w_034_558, w_002_070, w_009_002);
  and2 I034_559(w_034_559, w_008_117, w_029_291);
  nand2 I034_563(w_034_563, w_007_1484, w_028_026);
  nand2 I034_564(w_034_564, w_022_103, w_025_617);
  nand2 I034_566(w_034_566, w_032_175, w_013_291);
  and2 I034_568(w_034_568, w_030_305, w_008_404);
  and2 I034_569(w_034_569, w_029_1244, w_008_490);
  nand2 I034_570(w_034_570, w_005_290, w_009_000);
  nand2 I034_575(w_034_575, w_021_016, w_001_553);
  or2  I034_577(w_034_577, w_016_030, w_027_054);
  or2  I034_578(w_034_578, w_009_004, w_011_837);
  or2  I034_582(w_034_582, w_011_878, w_033_1461);
  not1 I034_583(w_034_583, w_019_618);
  nand2 I034_584(w_034_584, w_007_447, w_006_308);
  or2  I034_585(w_034_585, w_010_265, w_022_101);
  not1 I034_590(w_034_590, w_008_345);
  nand2 I034_592(w_034_592, w_033_1068, w_011_081);
  not1 I034_595(w_034_595, w_002_538);
  or2  I034_599(w_034_599, w_012_413, w_016_038);
  and2 I034_607(w_034_607, w_019_748, w_012_585);
  or2  I034_608(w_034_608, w_022_371, w_007_002);
  and2 I034_610(w_034_610, w_017_1640, w_000_1899);
  or2  I034_612(w_034_612, w_017_1517, w_008_077);
  nand2 I034_613(w_034_613, w_012_472, w_026_1296);
  and2 I034_620(w_034_620, w_005_1429, w_023_1412);
  not1 I034_621(w_034_621, w_033_655);
  not1 I034_630(w_034_630, w_005_072);
  or2  I034_649(w_034_649, w_018_192, w_031_848);
  nand2 I034_653(w_034_653, w_000_1226, w_029_718);
  or2  I034_657(w_034_657, w_024_125, w_026_020);
  nand2 I034_664(w_034_664, w_004_046, w_031_184);
  or2  I034_665(w_034_665, w_009_082, w_021_142);
  or2  I034_669(w_034_669, w_024_1438, w_007_563);
  nand2 I034_674(w_034_674, w_033_373, w_032_127);
  not1 I034_677(w_034_677, w_008_603);
  nand2 I034_680(w_034_680, w_005_1549, w_018_203);
  or2  I034_686(w_034_686, w_024_304, w_021_216);
  and2 I034_690(w_034_690, w_012_023, w_004_177);
  nand2 I035_003(w_035_003, w_015_176, w_022_368);
  nand2 I035_004(w_035_004, w_003_086, w_026_905);
  and2 I035_026(w_035_026, w_011_160, w_033_1098);
  nand2 I035_028(w_035_028, w_008_187, w_021_216);
  and2 I035_029(w_035_029, w_030_112, w_033_1523);
  and2 I035_036(w_035_036, w_028_783, w_009_044);
  nand2 I035_037(w_035_037, w_019_753, w_004_832);
  or2  I035_050(w_035_050, w_026_813, w_032_081);
  nand2 I035_051(w_035_051, w_033_361, w_032_036);
  or2  I035_052(w_035_052, w_025_1211, w_016_031);
  and2 I035_061(w_035_061, w_027_018, w_022_068);
  or2  I035_064(w_035_064, w_005_709, w_027_172);
  and2 I035_066(w_035_066, w_015_007, w_027_011);
  or2  I035_076(w_035_076, w_018_132, w_007_963);
  or2  I035_077(w_035_077, w_015_040, w_004_1292);
  and2 I035_083(w_035_083, w_029_243, w_031_038);
  nand2 I035_084(w_035_084, w_014_061, w_001_700);
  not1 I035_087(w_035_087, w_005_420);
  and2 I035_088(w_035_088, w_026_324, w_027_437);
  nand2 I035_091(w_035_091, w_006_156, w_034_227);
  not1 I035_095(w_035_095, w_034_613);
  nand2 I035_096(w_035_096, w_019_585, w_017_507);
  or2  I035_101(w_035_101, w_033_600, w_028_335);
  not1 I035_102(w_035_102, w_004_1300);
  or2  I035_103(w_035_103, w_000_1886, w_005_1007);
  not1 I035_104(w_035_104, w_029_1077);
  and2 I035_109(w_035_109, w_028_480, w_023_235);
  or2  I035_111(w_035_111, w_008_632, w_031_152);
  and2 I035_116(w_035_116, w_029_005, w_029_215);
  or2  I035_117(w_035_117, w_015_282, w_002_161);
  not1 I035_130(w_035_130, w_020_1017);
  and2 I035_134(w_035_134, w_017_159, w_029_1176);
  or2  I035_136(w_035_136, w_000_1838, w_008_108);
  nand2 I035_138(w_035_138, w_034_513, w_022_081);
  and2 I035_139(w_035_139, w_012_105, w_021_072);
  not1 I035_144(w_035_144, w_025_579);
  or2  I035_149(w_035_149, w_004_637, w_002_354);
  and2 I035_152(w_035_152, w_001_461, w_025_1280);
  and2 I035_160(w_035_160, w_004_1573, w_028_365);
  and2 I035_167(w_035_167, w_029_136, w_028_111);
  nand2 I035_168(w_035_168, w_034_379, w_031_643);
  or2  I035_175(w_035_175, w_033_1033, w_024_647);
  nand2 I035_188(w_035_188, w_001_244, w_004_837);
  or2  I035_194(w_035_194, w_031_778, w_024_1617);
  and2 I035_203(w_035_203, w_013_235, w_023_123);
  not1 I035_208(w_035_208, w_004_321);
  or2  I035_209(w_035_209, w_012_411, w_001_074);
  not1 I035_212(w_035_212, w_020_659);
  and2 I035_213(w_035_213, w_018_212, w_016_004);
  not1 I035_217(w_035_217, w_007_258);
  or2  I035_225(w_035_225, w_004_1731, w_000_361);
  or2  I035_228(w_035_228, w_005_208, w_020_231);
  nand2 I035_235(w_035_235, w_003_057, w_008_115);
  not1 I035_238(w_035_238, w_017_014);
  and2 I035_240(w_035_240, w_000_1910, w_026_443);
  nand2 I035_255(w_035_255, w_016_036, w_020_183);
  not1 I035_263(w_035_263, w_001_404);
  or2  I035_274(w_035_274, w_018_008, w_000_350);
  not1 I035_276(w_035_276, w_022_397);
  and2 I035_301(w_035_301, w_015_214, w_005_527);
  or2  I035_323(w_035_323, w_034_486, w_014_203);
  nand2 I035_328(w_035_328, w_014_184, w_010_280);
  nand2 I035_343(w_035_343, w_013_287, w_003_163);
  nand2 I035_349(w_035_349, w_029_022, w_028_674);
  nand2 I035_350(w_035_350, w_007_1313, w_015_149);
  or2  I035_351(w_035_351, w_020_582, w_026_079);
  and2 I035_352(w_035_352, w_011_016, w_027_038);
  nand2 I035_358(w_035_358, w_022_005, w_007_1294);
  or2  I035_397(w_035_397, w_030_696, w_021_097);
  and2 I035_433(w_035_433, w_009_013, w_001_330);
  nand2 I035_440(w_035_440, w_004_796, w_011_122);
  and2 I035_446(w_035_446, w_012_421, w_033_453);
  nand2 I035_460(w_035_460, w_016_003, w_015_236);
  or2  I035_467(w_035_467, w_008_207, w_029_1126);
  or2  I035_516(w_035_516, w_032_015, w_030_705);
  nand2 I035_520(w_035_520, w_034_526, w_020_650);
  and2 I035_546(w_035_546, w_000_1186, w_019_124);
  not1 I035_574(w_035_574, w_020_784);
  or2  I035_600(w_035_600, w_010_125, w_034_415);
  and2 I035_608(w_035_608, w_023_1004, w_008_434);
  nand2 I035_626(w_035_626, w_020_593, w_020_315);
  or2  I035_637(w_035_637, w_012_578, w_002_354);
  and2 I035_640(w_035_640, w_002_097, w_015_041);
  and2 I035_642(w_035_642, w_007_1175, w_016_002);
  or2  I035_643(w_035_643, w_005_129, w_000_100);
  nand2 I035_644(w_035_644, w_015_160, w_012_042);
  not1 I035_647(w_035_647, w_009_045);
  not1 I035_657(w_035_657, w_019_305);
  and2 I035_671(w_035_671, w_019_790, w_010_168);
  nand2 I035_678(w_035_678, w_025_1564, w_011_696);
  or2  I035_712(w_035_712, w_009_014, w_007_148);
  nand2 I035_722(w_035_722, w_031_848, w_023_1194);
  not1 I035_760(w_035_760, w_030_559);
  or2  I035_772(w_035_772, w_023_775, w_006_244);
  and2 I035_777(w_035_777, w_018_028, w_013_183);
  nand2 I035_804(w_035_804, w_013_121, w_032_025);
  not1 I035_805(w_035_805, w_014_314);
  nand2 I035_815(w_035_815, w_028_907, w_001_902);
  and2 I035_818(w_035_818, w_002_190, w_018_142);
  nand2 I035_832(w_035_832, w_014_436, w_021_136);
  or2  I035_840(w_035_840, w_017_684, w_017_1583);
  not1 I035_844(w_035_844, w_006_241);
  nand2 I035_848(w_035_848, w_030_412, w_014_213);
  and2 I035_861(w_035_861, w_003_060, w_029_1171);
  not1 I035_866(w_035_866, w_015_243);
  or2  I035_894(w_035_894, w_018_081, w_031_864);
  nand2 I035_908(w_035_908, w_017_528, w_004_1215);
  or2  I035_921(w_035_921, w_001_1603, w_007_1470);
  nand2 I035_936(w_035_936, w_007_135, w_033_631);
  and2 I035_938(w_035_938, w_017_158, w_004_1637);
  nand2 I035_941(w_035_941, w_020_440, w_008_256);
  or2  I035_976(w_035_976, w_022_173, w_029_470);
  not1 I035_987(w_035_987, w_020_093);
  and2 I035_991(w_035_991, w_010_102, w_018_103);
  or2  I035_996(w_035_996, w_009_059, w_013_184);
  and2 I035_997(w_035_997, w_011_144, w_004_1539);
  not1 I035_998(w_035_998, w_018_117);
  nand2 I035_999(w_035_999, w_013_119, w_021_036);
  or2  I035_1010(w_035_1010, w_015_127, w_002_315);
  and2 I035_1016(w_035_1016, w_025_253, w_020_480);
  not1 I035_1017(w_035_1017, w_027_563);
  or2  I035_1023(w_035_1023, w_012_663, w_010_359);
  or2  I035_1037(w_035_1037, w_012_469, w_000_1942);
  nand2 I035_1040(w_035_1040, w_012_369, w_023_088);
  or2  I035_1041(w_035_1041, w_017_240, w_009_039);
  not1 I035_1053(w_035_1053, w_027_422);
  not1 I035_1054(w_035_1054, w_031_150);
  not1 I035_1079(w_035_1079, w_021_075);
  or2  I035_1098(w_035_1098, w_026_1483, w_009_011);
  nand2 I035_1102(w_035_1102, w_028_705, w_007_002);
  and2 I035_1107(w_035_1107, w_000_1346, w_030_098);
  nand2 I035_1112(w_035_1112, w_002_360, w_019_1036);
  or2  I035_1119(w_035_1119, w_026_1070, w_027_408);
  nand2 I035_1125(w_035_1125, w_019_488, w_017_1556);
  or2  I035_1135(w_035_1135, w_006_117, w_023_236);
  nand2 I035_1146(w_035_1146, w_034_213, w_011_079);
  not1 I035_1147(w_035_1147, w_015_073);
  not1 I035_1176(w_035_1176, w_025_888);
  or2  I035_1198(w_035_1198, w_017_1269, w_034_557);
  nand2 I035_1203(w_035_1203, w_004_1017, w_032_000);
  or2  I035_1226(w_035_1226, w_018_172, w_002_155);
  not1 I035_1227(w_035_1227, w_013_292);
  and2 I035_1234(w_035_1234, w_020_085, w_030_220);
  or2  I035_1255(w_035_1255, w_002_222, w_004_530);
  nand2 I035_1267(w_035_1267, w_008_275, w_029_782);
  and2 I035_1273(w_035_1273, w_003_101, w_005_293);
  nand2 I035_1281(w_035_1281, w_033_923, w_031_422);
  and2 I035_1303(w_035_1303, w_017_558, w_034_677);
  and2 I035_1335(w_035_1335, w_021_242, w_024_869);
  or2  I035_1357(w_035_1357, w_028_070, w_013_077);
  nand2 I035_1371(w_035_1371, w_017_1000, w_028_668);
  not1 I035_1391(w_035_1391, w_030_071);
  nand2 I035_1397(w_035_1397, w_021_107, w_002_085);
  not1 I035_1425(w_035_1425, w_023_1569);
  or2  I035_1428(w_035_1428, w_000_1894, w_002_308);
  or2  I035_1431(w_035_1431, w_015_032, w_013_160);
  or2  I035_1437(w_035_1437, w_008_396, w_030_364);
  or2  I035_1450(w_035_1450, w_012_272, w_004_1128);
  not1 I035_1464(w_035_1464, w_010_074);
  nand2 I035_1471(w_035_1471, w_006_310, w_013_159);
  nand2 I035_1475(w_035_1475, w_005_1265, w_006_199);
  or2  I035_1484(w_035_1484, w_031_917, w_028_760);
  not1 I035_1485(w_035_1485, w_007_567);
  not1 I035_1487(w_035_1487, w_012_642);
  not1 I035_1502(w_035_1502, w_019_055);
  not1 I035_1506(w_035_1506, w_022_353);
  not1 I035_1510(w_035_1510, w_023_538);
  not1 I035_1513(w_035_1513, w_021_263);
  nand2 I035_1518(w_035_1518, w_024_480, w_003_249);
  or2  I035_1527(w_035_1527, w_026_450, w_013_300);
  or2  I035_1530(w_035_1530, w_019_229, w_013_044);
  nand2 I035_1546(w_035_1546, w_014_772, w_018_075);
  and2 I035_1585(w_035_1585, w_028_219, w_007_1492);
  not1 I035_1596(w_035_1596, w_011_109);
  not1 I035_1601(w_035_1601, w_005_766);
  and2 I035_1619(w_035_1619, w_022_298, w_011_578);
  or2  I035_1621(w_035_1621, w_015_160, w_001_044);
  nand2 I035_1646(w_035_1646, w_028_004, w_014_796);
  nand2 I035_1664(w_035_1664, w_006_322, w_003_148);
  nand2 I035_1671(w_035_1671, w_028_680, w_014_310);
  not1 I035_1673(w_035_1673, w_002_523);
  nand2 I035_1685(w_035_1685, w_029_631, w_029_792);
  nand2 I035_1707(w_035_1707, w_003_129, w_019_812);
  nand2 I035_1713(w_035_1713, w_003_274, w_034_686);
  or2  I035_1720(w_035_1720, w_028_666, w_024_164);
  not1 I036_018(w_036_018, w_006_120);
  not1 I036_025(w_036_025, w_023_759);
  not1 I036_029(w_036_029, w_028_317);
  or2  I036_032(w_036_032, w_025_479, w_012_531);
  not1 I036_033(w_036_033, w_016_019);
  not1 I036_037(w_036_037, w_011_094);
  not1 I036_045(w_036_045, w_009_078);
  not1 I036_047(w_036_047, w_034_203);
  nand2 I036_049(w_036_049, w_029_475, w_004_1537);
  not1 I036_056(w_036_056, w_026_1178);
  not1 I036_071(w_036_071, w_005_381);
  nand2 I036_079(w_036_079, w_027_091, w_020_750);
  and2 I036_085(w_036_085, w_004_1745, w_015_089);
  or2  I036_101(w_036_101, w_026_1155, w_034_418);
  not1 I036_107(w_036_107, w_026_227);
  not1 I036_114(w_036_114, w_001_1300);
  or2  I036_123(w_036_123, w_025_630, w_009_051);
  and2 I036_124(w_036_124, w_024_977, w_018_178);
  and2 I036_133(w_036_133, w_012_222, w_025_290);
  and2 I036_137(w_036_137, w_031_726, w_026_337);
  or2  I036_143(w_036_143, w_013_219, w_032_175);
  not1 I036_147(w_036_147, w_034_274);
  not1 I036_148(w_036_148, w_012_298);
  and2 I036_149(w_036_149, w_014_475, w_012_290);
  and2 I036_151(w_036_151, w_033_1619, w_030_630);
  and2 I036_161(w_036_161, w_023_986, w_028_592);
  not1 I036_166(w_036_166, w_003_027);
  or2  I036_169(w_036_169, w_013_132, w_028_311);
  or2  I036_170(w_036_170, w_015_222, w_007_1080);
  and2 I036_173(w_036_173, w_028_568, w_000_1422);
  nand2 I036_179(w_036_179, w_020_569, w_015_136);
  not1 I036_180(w_036_180, w_013_278);
  and2 I036_194(w_036_194, w_011_004, w_021_138);
  nand2 I036_196(w_036_196, w_003_289, w_014_342);
  or2  I036_199(w_036_199, w_013_090, w_024_1569);
  not1 I036_200(w_036_200, w_024_1545);
  nand2 I036_206(w_036_206, w_012_400, w_032_132);
  and2 I036_207(w_036_207, w_029_836, w_008_461);
  or2  I036_218(w_036_218, w_026_154, w_020_203);
  not1 I036_222(w_036_222, w_009_093);
  nand2 I036_226(w_036_226, w_028_641, w_003_281);
  not1 I036_238(w_036_238, w_011_883);
  nand2 I036_252(w_036_252, w_003_067, w_026_1202);
  and2 I036_255(w_036_255, w_022_015, w_006_126);
  not1 I036_256(w_036_256, w_012_438);
  nand2 I036_258(w_036_258, w_013_169, w_002_433);
  not1 I036_272(w_036_272, w_024_055);
  not1 I036_273(w_036_273, w_013_252);
  not1 I036_281(w_036_281, w_007_779);
  nand2 I036_282(w_036_282, w_021_253, w_006_241);
  nand2 I036_283(w_036_283, w_025_1094, w_028_716);
  and2 I036_297(w_036_297, w_006_342, w_012_205);
  or2  I036_310(w_036_310, w_026_1169, w_035_848);
  not1 I036_319(w_036_319, w_006_221);
  not1 I036_322(w_036_322, w_031_1021);
  or2  I036_323(w_036_323, w_021_010, w_010_375);
  nand2 I036_337(w_036_337, w_006_102, w_011_286);
  and2 I036_353(w_036_353, w_023_156, w_010_363);
  not1 I036_355(w_036_355, w_019_204);
  or2  I036_361(w_036_361, w_001_869, w_007_1515);
  not1 I036_369(w_036_369, w_023_136);
  and2 I036_374(w_036_374, w_007_1360, w_028_719);
  or2  I036_375(w_036_375, w_016_025, w_033_643);
  or2  I036_379(w_036_379, w_007_348, w_034_268);
  or2  I036_390(w_036_390, w_028_727, w_033_040);
  or2  I036_398(w_036_398, w_026_533, w_033_322);
  or2  I036_405(w_036_405, w_016_025, w_019_237);
  or2  I036_408(w_036_408, w_014_586, w_001_395);
  not1 I036_435(w_036_435, w_020_589);
  nand2 I036_441(w_036_441, w_019_864, w_034_578);
  and2 I036_450(w_036_450, w_011_037, w_002_413);
  not1 I036_451(w_036_451, w_000_1682);
  and2 I036_452(w_036_452, w_010_277, w_004_1905);
  nand2 I036_454(w_036_454, w_004_368, w_011_194);
  nand2 I036_456(w_036_456, w_003_046, w_008_318);
  or2  I036_481(w_036_481, w_028_070, w_009_034);
  or2  I036_482(w_036_482, w_009_006, w_032_081);
  and2 I036_486(w_036_486, w_000_880, w_015_080);
  or2  I036_488(w_036_488, w_009_051, w_022_331);
  nand2 I036_492(w_036_492, w_018_256, w_010_231);
  and2 I036_493(w_036_493, w_010_244, w_024_610);
  not1 I036_495(w_036_495, w_012_561);
  and2 I036_496(w_036_496, w_011_771, w_035_050);
  and2 I036_505(w_036_505, w_000_039, w_023_474);
  nand2 I036_513(w_036_513, w_023_414, w_013_025);
  nand2 I036_525(w_036_525, w_011_093, w_019_284);
  or2  I036_538(w_036_538, w_033_314, w_034_308);
  nand2 I036_543(w_036_543, w_027_184, w_020_191);
  or2  I036_577(w_036_577, w_016_012, w_012_020);
  and2 I036_580(w_036_580, w_001_873, w_020_381);
  nand2 I036_585(w_036_585, w_009_076, w_018_049);
  and2 I036_589(w_036_589, w_023_624, w_011_811);
  and2 I036_594(w_036_594, w_024_082, w_009_097);
  nand2 I036_596(w_036_596, w_012_322, w_005_771);
  or2  I036_650(w_036_650, w_005_1616, w_035_076);
  or2  I036_652(w_036_652, w_001_1607, w_008_208);
  nand2 I036_657(w_036_657, w_018_113, w_017_1738);
  not1 I036_692(w_036_692, w_026_699);
  nand2 I036_696(w_036_696, w_025_707, w_012_129);
  and2 I036_697(w_036_697, w_002_264, w_003_027);
  not1 I036_702(w_036_702, w_013_021);
  and2 I036_712(w_036_712, w_018_012, w_006_146);
  or2  I036_713(w_036_713, w_015_171, w_016_000);
  or2  I036_723(w_036_723, w_015_077, w_007_715);
  not1 I036_728(w_036_728, w_005_072);
  or2  I036_764(w_036_764, w_032_046, w_007_051);
  or2  I036_778(w_036_778, w_003_308, w_016_013);
  nand2 I036_781(w_036_781, w_024_1225, w_003_103);
  or2  I036_786(w_036_786, w_033_081, w_014_393);
  and2 I036_790(w_036_790, w_024_830, w_004_057);
  nand2 I036_803(w_036_803, w_014_169, w_002_412);
  not1 I036_813(w_036_813, w_010_126);
  or2  I036_815(w_036_815, w_025_081, w_013_132);
  nand2 I036_826(w_036_826, w_018_092, w_006_110);
  nand2 I036_837(w_036_837, w_013_100, w_028_463);
  and2 I036_842(w_036_842, w_003_052, w_015_034);
  or2  I036_850(w_036_850, w_018_132, w_018_143);
  or2  I036_866(w_036_866, w_020_1202, w_030_781);
  or2  I036_875(w_036_875, w_034_528, w_014_235);
  nand2 I036_880(w_036_880, w_017_436, w_014_486);
  and2 I036_895(w_036_895, w_026_097, w_002_138);
  and2 I036_914(w_036_914, w_018_139, w_001_139);
  nand2 I036_924(w_036_924, w_011_193, w_034_665);
  nand2 I036_937(w_036_937, w_010_105, w_019_338);
  nand2 I036_939(w_036_939, w_033_064, w_004_1288);
  or2  I036_953(w_036_953, w_019_273, w_035_350);
  nand2 I036_965(w_036_965, w_031_546, w_004_1530);
  nand2 I036_972(w_036_972, w_027_364, w_014_780);
  or2  I036_978(w_036_978, w_033_869, w_009_004);
  not1 I036_982(w_036_982, w_023_635);
  nand2 I036_992(w_036_992, w_011_242, w_027_328);
  not1 I036_1005(w_036_1005, w_029_129);
  not1 I036_1014(w_036_1014, w_012_159);
  not1 I036_1023(w_036_1023, w_029_755);
  and2 I036_1034(w_036_1034, w_003_218, w_014_416);
  and2 I036_1043(w_036_1043, w_021_250, w_019_843);
  or2  I036_1049(w_036_1049, w_004_587, w_014_481);
  and2 I036_1071(w_036_1071, w_002_385, w_023_1275);
  nand2 I036_1076(w_036_1076, w_019_1089, w_029_589);
  and2 I036_1104(w_036_1104, w_011_345, w_023_282);
  nand2 I036_1107(w_036_1107, w_016_019, w_001_1128);
  nand2 I036_1114(w_036_1114, w_033_1318, w_032_089);
  or2  I036_1115(w_036_1115, w_031_712, w_029_453);
  or2  I036_1129(w_036_1129, w_015_133, w_035_134);
  not1 I036_1139(w_036_1139, w_006_310);
  not1 I036_1140(w_036_1140, w_012_400);
  not1 I036_1149(w_036_1149, w_035_1135);
  or2  I036_1150(w_036_1150, w_009_023, w_027_523);
  and2 I036_1153(w_036_1153, w_002_433, w_020_068);
  nand2 I036_1174(w_036_1174, w_024_606, w_024_044);
  or2  I036_1210(w_036_1210, w_015_015, w_032_032);
  or2  I036_1217(w_036_1217, w_029_693, w_016_004);
  not1 I036_1218(w_036_1218, w_006_129);
  and2 I036_1220(w_036_1220, w_011_539, w_017_821);
  not1 I036_1222(w_036_1222, w_034_545);
  and2 I036_1226(w_036_1226, w_014_197, w_011_074);
  not1 I036_1227(w_036_1227, w_016_005);
  and2 I036_1234(w_036_1234, w_007_1176, w_016_009);
  nand2 I036_1237(w_036_1237, w_033_195, w_002_568);
  and2 I036_1239(w_036_1239, w_000_581, w_035_084);
  and2 I036_1273(w_036_1273, w_003_019, w_033_979);
  and2 I036_1289(w_036_1289, w_027_440, w_016_037);
  or2  I036_1294(w_036_1294, w_008_762, w_007_941);
  not1 I036_1306(w_036_1306, w_015_238);
  and2 I036_1309(w_036_1309, w_025_100, w_018_268);
  or2  I036_1320(w_036_1320, w_021_149, w_019_817);
  or2  I036_1325(w_036_1325, w_031_087, w_003_101);
  nand2 I036_1336(w_036_1336, w_002_492, w_007_1227);
  nand2 I036_1339(w_036_1339, w_005_1153, w_008_417);
  and2 I036_1341(w_036_1341, w_020_228, w_029_494);
  or2  I036_1346(w_036_1346, w_001_1144, w_013_154);
  and2 I036_1356(w_036_1356, w_020_333, w_033_191);
  and2 I036_1366(w_036_1366, w_017_360, w_025_230);
  not1 I036_1373(w_036_1373, w_004_1445);
  or2  I036_1379(w_036_1379, w_026_1016, w_010_261);
  nand2 I036_1397(w_036_1397, w_009_076, w_021_047);
  nand2 I036_1399(w_036_1399, w_027_585, w_022_367);
  or2  I036_1406(w_036_1406, w_013_097, w_028_243);
  not1 I036_1426(w_036_1426, w_008_796);
  not1 I036_1438(w_036_1438, w_008_197);
  or2  I036_1440(w_036_1440, w_010_127, w_019_097);
  and2 I036_1454(w_036_1454, w_008_005, w_022_129);
  or2  I036_1457(w_036_1457, w_016_028, w_016_014);
  and2 I036_1464(w_036_1464, w_029_347, w_009_082);
  not1 I036_1473(w_036_1473, w_001_1323);
  nand2 I036_1475(w_036_1475, w_022_109, w_000_270);
  nand2 I036_1481(w_036_1481, w_003_225, w_022_053);
  or2  I036_1493(w_036_1493, w_001_413, w_020_727);
  not1 I037_001(w_037_001, w_030_633);
  nand2 I037_007(w_037_007, w_000_1962, w_026_1277);
  and2 I037_028(w_037_028, w_006_317, w_024_1050);
  not1 I037_046(w_037_046, w_014_728);
  or2  I037_055(w_037_055, w_010_250, w_025_1549);
  not1 I037_072(w_037_072, w_008_090);
  nand2 I037_076(w_037_076, w_003_077, w_027_032);
  and2 I037_081(w_037_081, w_018_061, w_019_776);
  and2 I037_085(w_037_085, w_015_011, w_007_564);
  not1 I037_090(w_037_090, w_009_100);
  and2 I037_098(w_037_098, w_031_983, w_020_298);
  or2  I037_111(w_037_111, w_025_938, w_006_148);
  not1 I037_114(w_037_114, w_021_061);
  not1 I037_119(w_037_119, w_015_243);
  not1 I037_137(w_037_137, w_018_152);
  nand2 I037_143(w_037_143, w_003_034, w_027_447);
  not1 I037_145(w_037_145, w_001_014);
  and2 I037_155(w_037_155, w_002_220, w_020_549);
  nand2 I037_156(w_037_156, w_032_195, w_023_1612);
  nand2 I037_157(w_037_157, w_033_283, w_034_564);
  and2 I037_160(w_037_160, w_004_512, w_017_1139);
  nand2 I037_161(w_037_161, w_036_1341, w_017_1351);
  and2 I037_175(w_037_175, w_019_395, w_027_371);
  not1 I037_188(w_037_188, w_027_057);
  not1 I037_190(w_037_190, w_017_1422);
  and2 I037_193(w_037_193, w_030_082, w_030_641);
  and2 I037_197(w_037_197, w_021_193, w_009_078);
  and2 I037_201(w_037_201, w_024_1624, w_036_226);
  or2  I037_210(w_037_210, w_019_960, w_004_402);
  not1 I037_219(w_037_219, w_021_169);
  nand2 I037_222(w_037_222, w_006_083, w_023_004);
  nand2 I037_226(w_037_226, w_035_255, w_008_049);
  nand2 I037_262(w_037_262, w_026_1456, w_003_002);
  or2  I037_303(w_037_303, w_015_227, w_009_050);
  or2  I037_324(w_037_324, w_019_849, w_003_121);
  not1 I037_328(w_037_328, w_018_045);
  not1 I037_352(w_037_352, w_010_061);
  nand2 I037_355(w_037_355, w_007_839, w_033_847);
  or2  I037_363(w_037_363, w_005_597, w_008_836);
  or2  I037_372(w_037_372, w_007_1132, w_009_038);
  or2  I037_387(w_037_387, w_029_1124, w_034_044);
  and2 I037_407(w_037_407, w_013_335, w_017_1586);
  and2 I037_438(w_037_438, w_025_573, w_027_524);
  and2 I037_446(w_037_446, w_011_503, w_005_875);
  not1 I037_496(w_037_496, w_001_631);
  not1 I037_502(w_037_502, w_011_100);
  not1 I037_508(w_037_508, w_019_551);
  not1 I037_510(w_037_510, w_026_257);
  or2  I037_517(w_037_517, w_004_1900, w_008_104);
  or2  I037_519(w_037_519, w_004_1643, w_035_626);
  nand2 I037_535(w_037_535, w_031_337, w_027_109);
  or2  I037_541(w_037_541, w_029_1092, w_025_1597);
  or2  I037_547(w_037_547, w_025_679, w_021_020);
  not1 I037_553(w_037_553, w_019_860);
  not1 I037_563(w_037_563, w_003_201);
  nand2 I037_567(w_037_567, w_014_118, w_016_019);
  nand2 I037_594(w_037_594, w_005_253, w_028_024);
  or2  I037_604(w_037_604, w_007_1484, w_023_010);
  not1 I037_607(w_037_607, w_007_155);
  or2  I037_627(w_037_627, w_017_1379, w_001_208);
  nand2 I037_629(w_037_629, w_019_706, w_000_008);
  or2  I037_633(w_037_633, w_003_088, w_001_045);
  or2  I037_649(w_037_649, w_006_040, w_003_250);
  nand2 I037_669(w_037_669, w_022_248, w_031_517);
  and2 I037_670(w_037_670, w_004_661, w_027_475);
  not1 I037_674(w_037_674, w_002_181);
  not1 I037_675(w_037_675, w_007_682);
  and2 I037_679(w_037_679, w_029_402, w_013_186);
  not1 I037_684(w_037_684, w_013_167);
  or2  I037_690(w_037_690, w_005_600, w_011_117);
  or2  I037_702(w_037_702, w_024_1203, w_018_171);
  and2 I037_705(w_037_705, w_027_276, w_032_042);
  nand2 I037_706(w_037_706, w_004_900, w_036_1222);
  not1 I037_713(w_037_713, w_027_081);
  or2  I037_741(w_037_741, w_008_349, w_016_010);
  nand2 I037_745(w_037_745, w_021_018, w_002_206);
  nand2 I037_765(w_037_765, w_002_293, w_002_486);
  and2 I037_774(w_037_774, w_030_572, w_008_537);
  and2 I037_777(w_037_777, w_012_435, w_003_113);
  nand2 I037_778(w_037_778, w_011_107, w_029_130);
  not1 I037_793(w_037_793, w_031_145);
  nand2 I037_804(w_037_804, w_033_004, w_007_1328);
  nand2 I037_807(w_037_807, w_023_187, w_036_1218);
  not1 I037_812(w_037_812, w_019_409);
  nand2 I037_849(w_037_849, w_007_834, w_017_299);
  not1 I037_876(w_037_876, w_005_096);
  not1 I037_879(w_037_879, w_019_478);
  and2 I037_884(w_037_884, w_012_100, w_001_544);
  not1 I037_900(w_037_900, w_018_230);
  not1 I037_901(w_037_901, w_030_638);
  or2  I037_906(w_037_906, w_021_095, w_019_745);
  or2  I037_923(w_037_923, w_036_1454, w_017_896);
  not1 I037_939(w_037_939, w_001_529);
  or2  I037_942(w_037_942, w_003_245, w_023_776);
  nand2 I037_949(w_037_949, w_014_380, w_006_325);
  not1 I037_953(w_037_953, w_030_169);
  not1 I037_982(w_037_982, w_006_251);
  and2 I037_998(w_037_998, w_000_803, w_000_823);
  nand2 I037_999(w_037_999, w_033_485, w_005_098);
  or2  I037_1000(w_037_1000, w_031_123, w_029_440);
  not1 I037_1035(w_037_1035, w_011_307);
  not1 I037_1050(w_037_1050, w_025_1084);
  or2  I037_1054(w_037_1054, w_022_075, w_013_271);
  nand2 I037_1076(w_037_1076, w_015_166, w_009_053);
  not1 I037_1081(w_037_1081, w_018_146);
  not1 I037_1083(w_037_1083, w_014_161);
  not1 I037_1084(w_037_1084, w_029_550);
  not1 I037_1088(w_037_1088, w_034_182);
  not1 I037_1103(w_037_1103, w_036_1115);
  nand2 I037_1106(w_037_1106, w_015_164, w_023_1567);
  not1 I037_1108(w_037_1108, w_036_1149);
  or2  I037_1128(w_037_1128, w_004_080, w_030_017);
  nand2 I037_1132(w_037_1132, w_013_181, w_032_009);
  nand2 I037_1140(w_037_1140, w_011_508, w_025_1575);
  not1 I037_1149(w_037_1149, w_029_033);
  and2 I037_1177(w_037_1177, w_004_1720, w_031_359);
  not1 I037_1186(w_037_1186, w_007_210);
  not1 I037_1194(w_037_1194, w_031_370);
  and2 I037_1210(w_037_1210, w_005_1243, w_020_371);
  and2 I037_1211(w_037_1211, w_010_250, w_031_713);
  not1 I037_1234(w_037_1234, w_010_172);
  nand2 I037_1238(w_037_1238, w_013_062, w_029_136);
  nand2 I037_1254(w_037_1254, w_017_457, w_034_504);
  and2 I037_1259(w_037_1259, w_022_329, w_032_153);
  and2 I037_1278(w_037_1278, w_022_225, w_016_030);
  nand2 I037_1290(w_037_1290, w_031_815, w_004_1320);
  not1 I037_1292(w_037_1292, w_032_155);
  not1 I037_1307(w_037_1307, w_028_095);
  or2  I037_1309(w_037_1309, w_014_383, w_021_166);
  not1 I037_1320(w_037_1320, w_003_153);
  nand2 I037_1329(w_037_1329, w_002_498, w_014_478);
  not1 I037_1339(w_037_1339, w_029_477);
  not1 I037_1340(w_037_1340, w_000_1086);
  and2 I037_1343(w_037_1343, w_028_889, w_017_631);
  nand2 I037_1344(w_037_1344, w_021_107, w_004_186);
  nand2 I037_1349(w_037_1349, w_007_152, w_000_1526);
  and2 I037_1357(w_037_1357, w_035_168, w_019_383);
  nand2 I037_1389(w_037_1389, w_012_555, w_018_216);
  or2  I037_1406(w_037_1406, w_023_176, w_023_459);
  and2 I037_1421(w_037_1421, w_024_874, w_001_1025);
  or2  I037_1422(w_037_1422, w_018_181, w_024_153);
  or2  I037_1432(w_037_1432, w_031_521, w_013_260);
  and2 I037_1441(w_037_1441, w_028_155, w_033_1436);
  and2 I037_1451(w_037_1451, w_010_357, w_024_313);
  or2  I037_1461(w_037_1461, w_022_059, w_017_1397);
  nand2 I037_1462(w_037_1462, w_002_399, w_014_270);
  or2  I037_1488(w_037_1488, w_010_398, w_011_204);
  nand2 I037_1489(w_037_1489, w_009_039, w_026_1376);
  and2 I037_1494(w_037_1494, w_022_023, w_024_1055);
  not1 I037_1500(w_037_1500, w_011_213);
  not1 I037_1520(w_037_1520, w_013_154);
  and2 I037_1528(w_037_1528, w_018_030, w_013_073);
  nand2 I037_1531(w_037_1531, w_025_1452, w_007_1405);
  and2 I037_1532(w_037_1532, w_014_387, w_009_012);
  not1 I037_1541(w_037_1541, w_014_124);
  not1 I037_1554(w_037_1554, w_027_155);
  and2 I037_1602(w_037_1602, w_026_1253, w_001_660);
  not1 I037_1625(w_037_1625, w_009_019);
  or2  I037_1637(w_037_1637, w_017_427, w_004_063);
  nand2 I037_1646(w_037_1646, w_033_326, w_019_206);
  and2 I037_1656(w_037_1656, w_010_059, w_014_089);
  and2 I037_1659(w_037_1659, w_009_042, w_009_078);
  nand2 I037_1674(w_037_1674, w_030_549, w_030_706);
  not1 I037_1676(w_037_1676, w_035_066);
  not1 I037_1678(w_037_1678, w_009_027);
  and2 I037_1679(w_037_1679, w_000_620, w_035_358);
  nand2 I037_1689(w_037_1689, w_028_589, w_021_147);
  or2  I037_1694(w_037_1694, w_011_094, w_020_714);
  not1 I037_1711(w_037_1711, w_011_369);
  not1 I037_1730(w_037_1730, w_005_1157);
  nand2 I038_002(w_038_002, w_018_205, w_008_795);
  not1 I038_006(w_038_006, w_031_917);
  or2  I038_007(w_038_007, w_023_029, w_004_1616);
  or2  I038_012(w_038_012, w_032_202, w_010_190);
  and2 I038_015(w_038_015, w_013_217, w_001_657);
  and2 I038_019(w_038_019, w_017_556, w_027_226);
  not1 I038_021(w_038_021, w_009_025);
  not1 I038_022(w_038_022, w_022_251);
  or2  I038_027(w_038_027, w_002_338, w_014_677);
  or2  I038_028(w_038_028, w_022_123, w_000_1125);
  or2  I038_031(w_038_031, w_028_114, w_032_239);
  and2 I038_034(w_038_034, w_015_181, w_005_1180);
  not1 I038_039(w_038_039, w_006_048);
  and2 I038_043(w_038_043, w_035_235, w_030_716);
  or2  I038_045(w_038_045, w_033_069, w_013_313);
  and2 I038_048(w_038_048, w_035_866, w_034_418);
  nand2 I038_049(w_038_049, w_016_010, w_017_1622);
  or2  I038_052(w_038_052, w_020_290, w_002_500);
  nand2 I038_055(w_038_055, w_036_652, w_013_296);
  or2  I038_058(w_038_058, w_034_513, w_008_547);
  not1 I038_061(w_038_061, w_024_178);
  or2  I038_063(w_038_063, w_036_585, w_033_1444);
  nand2 I038_065(w_038_065, w_029_110, w_024_072);
  or2  I038_068(w_038_068, w_012_451, w_005_841);
  nand2 I038_073(w_038_073, w_003_043, w_021_082);
  or2  I038_076(w_038_076, w_025_1222, w_023_169);
  not1 I038_077(w_038_077, w_032_032);
  and2 I038_081(w_038_081, w_003_025, w_001_488);
  nand2 I038_084(w_038_084, w_025_1309, w_020_178);
  and2 I038_100(w_038_100, w_030_309, w_017_944);
  not1 I038_108(w_038_108, w_011_262);
  not1 I038_109(w_038_109, w_026_317);
  not1 I038_111(w_038_111, w_018_148);
  and2 I038_112(w_038_112, w_036_252, w_033_482);
  or2  I038_113(w_038_113, w_030_525, w_033_260);
  not1 I038_118(w_038_118, w_002_569);
  nand2 I038_122(w_038_122, w_037_076, w_035_1671);
  and2 I038_130(w_038_130, w_015_218, w_021_191);
  or2  I038_134(w_038_134, w_010_391, w_000_1246);
  or2  I038_136(w_038_136, w_028_530, w_009_063);
  and2 I038_141(w_038_141, w_020_1121, w_020_295);
  and2 I038_144(w_038_144, w_008_570, w_021_093);
  not1 I038_148(w_038_148, w_004_345);
  or2  I038_150(w_038_150, w_016_026, w_012_288);
  nand2 I038_152(w_038_152, w_002_505, w_013_335);
  not1 I038_153(w_038_153, w_008_470);
  or2  I038_155(w_038_155, w_023_1196, w_035_1226);
  and2 I038_158(w_038_158, w_034_090, w_000_1011);
  and2 I038_160(w_038_160, w_005_706, w_036_1473);
  not1 I038_161(w_038_161, w_027_411);
  nand2 I038_170(w_038_170, w_002_204, w_022_085);
  or2  I038_173(w_038_173, w_031_500, w_034_034);
  not1 I038_175(w_038_175, w_034_513);
  and2 I038_178(w_038_178, w_015_144, w_011_652);
  not1 I038_181(w_038_181, w_025_1048);
  not1 I038_183(w_038_183, w_020_1131);
  and2 I038_186(w_038_186, w_031_210, w_003_079);
  not1 I038_192(w_038_192, w_012_287);
  and2 I038_196(w_038_196, w_025_1174, w_005_1478);
  not1 I038_198(w_038_198, w_005_1420);
  and2 I038_200(w_038_200, w_012_233, w_024_288);
  or2  I038_201(w_038_201, w_018_180, w_004_590);
  or2  I038_207(w_038_207, w_008_764, w_007_077);
  and2 I038_208(w_038_208, w_015_061, w_002_225);
  nand2 I038_211(w_038_211, w_036_924, w_023_1046);
  not1 I038_221(w_038_221, w_009_033);
  and2 I038_224(w_038_224, w_007_1531, w_010_276);
  not1 I038_227(w_038_227, w_037_098);
  nand2 I038_233(w_038_233, w_003_042, w_024_003);
  or2  I038_235(w_038_235, w_035_1596, w_005_052);
  or2  I038_236(w_038_236, w_019_487, w_014_323);
  or2  I038_239(w_038_239, w_025_101, w_018_241);
  and2 I038_255(w_038_255, w_033_244, w_000_459);
  or2  I038_256(w_038_256, w_031_510, w_035_160);
  and2 I038_258(w_038_258, w_022_281, w_008_457);
  or2  I038_260(w_038_260, w_003_050, w_033_1018);
  and2 I038_263(w_038_263, w_010_270, w_002_146);
  and2 I038_265(w_038_265, w_013_021, w_006_220);
  not1 I038_269(w_038_269, w_002_087);
  nand2 I038_276(w_038_276, w_009_008, w_024_1473);
  nand2 I038_281(w_038_281, w_036_390, w_028_855);
  not1 I038_287(w_038_287, w_026_218);
  or2  I038_290(w_038_290, w_019_386, w_011_870);
  and2 I038_299(w_038_299, w_033_107, w_032_193);
  and2 I038_300(w_038_300, w_031_513, w_035_832);
  and2 I038_302(w_038_302, w_014_005, w_035_351);
  nand2 I038_304(w_038_304, w_027_258, w_008_424);
  or2  I038_308(w_038_308, w_000_857, w_015_129);
  not1 I038_317(w_038_317, w_023_299);
  not1 I038_319(w_038_319, w_016_017);
  not1 I038_320(w_038_320, w_033_1280);
  or2  I038_325(w_038_325, w_009_108, w_019_729);
  and2 I038_327(w_038_327, w_008_172, w_005_149);
  nand2 I038_331(w_038_331, w_037_949, w_008_185);
  not1 I038_332(w_038_332, w_034_599);
  nand2 I038_333(w_038_333, w_031_597, w_030_079);
  or2  I038_335(w_038_335, w_016_012, w_037_1290);
  nand2 I038_337(w_038_337, w_029_273, w_002_459);
  nand2 I038_338(w_038_338, w_027_376, w_027_209);
  nand2 I038_339(w_038_339, w_007_1524, w_034_407);
  not1 I038_345(w_038_345, w_011_046);
  nand2 I038_348(w_038_348, w_021_233, w_022_393);
  and2 I038_353(w_038_353, w_023_1007, w_002_327);
  not1 I038_362(w_038_362, w_008_009);
  not1 I038_364(w_038_364, w_022_213);
  nand2 I038_366(w_038_366, w_000_1080, w_030_181);
  not1 I038_367(w_038_367, w_006_244);
  and2 I038_368(w_038_368, w_000_1525, w_012_375);
  not1 I038_372(w_038_372, w_029_810);
  nand2 I038_378(w_038_378, w_030_248, w_028_653);
  nand2 I038_382(w_038_382, w_004_620, w_008_813);
  nand2 I038_384(w_038_384, w_032_211, w_015_077);
  or2  I038_385(w_038_385, w_008_342, w_037_1088);
  not1 I038_387(w_038_387, w_029_450);
  not1 I038_390(w_038_390, w_015_173);
  and2 I038_391(w_038_391, w_018_246, w_006_098);
  and2 I038_392(w_038_392, w_037_324, w_016_022);
  or2  I038_395(w_038_395, w_035_1621, w_016_022);
  or2  I038_397(w_038_397, w_037_627, w_017_324);
  not1 I038_400(w_038_400, w_023_277);
  and2 I038_401(w_038_401, w_034_406, w_035_1040);
  nand2 I038_402(w_038_402, w_016_034, w_036_1071);
  and2 I038_404(w_038_404, w_024_035, w_017_885);
  and2 I038_405(w_038_405, w_013_053, w_016_022);
  and2 I038_410(w_038_410, w_025_1350, w_013_125);
  not1 I038_412(w_038_412, w_015_039);
  or2  I038_413(w_038_413, w_004_785, w_003_212);
  and2 I038_429(w_038_429, w_023_1573, w_026_671);
  or2  I038_438(w_038_438, w_007_1304, w_027_129);
  or2  I038_439(w_038_439, w_000_1311, w_012_567);
  and2 I038_448(w_038_448, w_018_040, w_011_698);
  and2 I038_451(w_038_451, w_024_146, w_028_217);
  or2  I038_454(w_038_454, w_023_280, w_007_444);
  or2  I038_457(w_038_457, w_024_842, w_031_611);
  and2 I038_458(w_038_458, w_032_236, w_029_901);
  nand2 I038_459(w_038_459, w_022_267, w_025_1671);
  or2  I038_464(w_038_464, w_012_590, w_021_087);
  nand2 I038_473(w_038_473, w_030_804, w_005_1101);
  not1 I038_475(w_038_475, w_008_165);
  or2  I038_479(w_038_479, w_017_1098, w_026_1097);
  not1 I038_480(w_038_480, w_034_419);
  nand2 I038_484(w_038_484, w_018_003, w_010_108);
  and2 I038_485(w_038_485, w_000_054, w_022_298);
  and2 I038_486(w_038_486, w_010_273, w_002_086);
  not1 I039_007(w_039_007, w_037_1340);
  nand2 I039_018(w_039_018, w_033_332, w_004_399);
  not1 I039_024(w_039_024, w_004_1211);
  nand2 I039_025(w_039_025, w_008_233, w_008_286);
  or2  I039_027(w_039_027, w_021_088, w_029_354);
  not1 I039_033(w_039_033, w_037_1694);
  not1 I039_065(w_039_065, w_029_178);
  and2 I039_075(w_039_075, w_011_103, w_038_112);
  and2 I039_087(w_039_087, w_021_147, w_000_1861);
  nand2 I039_092(w_039_092, w_013_198, w_036_1114);
  nand2 I039_100(w_039_100, w_013_155, w_028_528);
  nand2 I039_113(w_039_113, w_024_1478, w_035_301);
  nand2 I039_133(w_039_133, w_024_1032, w_024_277);
  nand2 I039_135(w_039_135, w_005_1321, w_028_160);
  or2  I039_142(w_039_142, w_013_073, w_035_1428);
  nand2 I039_167(w_039_167, w_009_102, w_013_144);
  or2  I039_178(w_039_178, w_017_303, w_017_838);
  not1 I039_198(w_039_198, w_033_1249);
  nand2 I039_199(w_039_199, w_030_218, w_012_133);
  not1 I039_204(w_039_204, w_035_274);
  nand2 I039_250(w_039_250, w_029_1281, w_016_025);
  not1 I039_252(w_039_252, w_012_393);
  and2 I039_259(w_039_259, w_022_113, w_028_004);
  and2 I039_260(w_039_260, w_020_668, w_031_250);
  and2 I039_266(w_039_266, w_028_683, w_001_1167);
  and2 I039_272(w_039_272, w_004_1267, w_024_888);
  nand2 I039_289(w_039_289, w_034_248, w_003_191);
  nand2 I039_306(w_039_306, w_019_953, w_016_021);
  and2 I039_310(w_039_310, w_016_035, w_026_288);
  and2 I039_313(w_039_313, w_013_061, w_009_016);
  and2 I039_347(w_039_347, w_019_409, w_012_139);
  nand2 I039_351(w_039_351, w_023_818, w_018_219);
  nand2 I039_415(w_039_415, w_027_040, w_007_393);
  not1 I039_429(w_039_429, w_020_652);
  and2 I039_466(w_039_466, w_017_1423, w_028_275);
  or2  I039_470(w_039_470, w_011_070, w_019_250);
  or2  I039_477(w_039_477, w_031_766, w_005_143);
  not1 I039_482(w_039_482, w_002_466);
  nand2 I039_490(w_039_490, w_031_635, w_034_297);
  not1 I039_501(w_039_501, w_038_061);
  not1 I039_507(w_039_507, w_002_218);
  not1 I039_516(w_039_516, w_007_1469);
  and2 I039_526(w_039_526, w_026_1507, w_024_269);
  nand2 I039_530(w_039_530, w_019_791, w_020_606);
  and2 I039_533(w_039_533, w_010_056, w_013_133);
  and2 I039_558(w_039_558, w_020_745, w_011_221);
  or2  I039_568(w_039_568, w_007_576, w_005_596);
  or2  I039_595(w_039_595, w_024_000, w_000_995);
  nand2 I039_597(w_039_597, w_023_667, w_016_002);
  not1 I039_599(w_039_599, w_029_477);
  nand2 I039_610(w_039_610, w_003_300, w_017_317);
  not1 I039_612(w_039_612, w_016_025);
  and2 I039_614(w_039_614, w_012_204, w_001_029);
  not1 I039_618(w_039_618, w_005_262);
  nand2 I039_629(w_039_629, w_036_702, w_001_153);
  nand2 I039_631(w_039_631, w_022_219, w_002_346);
  or2  I039_648(w_039_648, w_027_074, w_000_1198);
  or2  I039_650(w_039_650, w_038_077, w_015_176);
  nand2 I039_665(w_039_665, w_027_413, w_036_965);
  and2 I039_676(w_039_676, w_013_217, w_017_023);
  not1 I039_687(w_039_687, w_019_717);
  and2 I039_707(w_039_707, w_023_049, w_038_402);
  or2  I039_714(w_039_714, w_007_269, w_002_504);
  and2 I039_721(w_039_721, w_022_008, w_017_984);
  not1 I039_726(w_039_726, w_009_102);
  or2  I039_752(w_039_752, w_022_210, w_006_004);
  or2  I039_759(w_039_759, w_016_021, w_016_033);
  and2 I039_775(w_039_775, w_023_111, w_012_442);
  not1 I039_782(w_039_782, w_025_1538);
  or2  I039_788(w_039_788, w_022_409, w_025_1633);
  or2  I039_793(w_039_793, w_020_662, w_033_1136);
  or2  I039_805(w_039_805, w_029_258, w_018_259);
  nand2 I039_834(w_039_834, w_030_173, w_026_024);
  nand2 I039_835(w_039_835, w_003_302, w_011_297);
  not1 I039_842(w_039_842, w_031_394);
  or2  I039_847(w_039_847, w_017_1051, w_021_009);
  not1 I039_879(w_039_879, w_038_239);
  not1 I039_881(w_039_881, w_037_1500);
  or2  I039_895(w_039_895, w_010_125, w_030_314);
  not1 I039_910(w_039_910, w_028_727);
  and2 I039_915(w_039_915, w_032_009, w_019_699);
  nand2 I039_932(w_039_932, w_008_108, w_013_251);
  or2  I039_933(w_039_933, w_017_085, w_019_353);
  or2  I039_936(w_039_936, w_026_1467, w_010_328);
  and2 I039_938(w_039_938, w_009_027, w_015_218);
  not1 I039_969(w_039_969, w_026_110);
  or2  I039_977(w_039_977, w_006_082, w_020_488);
  not1 I039_1009(w_039_1009, w_015_186);
  or2  I039_1059(w_039_1059, w_012_362, w_002_461);
  and2 I039_1065(w_039_1065, w_011_246, w_037_1541);
  and2 I039_1078(w_039_1078, w_007_130, w_028_853);
  or2  I039_1097(w_039_1097, w_010_067, w_027_190);
  not1 I039_1126(w_039_1126, w_004_724);
  not1 I039_1145(w_039_1145, w_014_025);
  nand2 I039_1151(w_039_1151, w_023_546, w_019_420);
  not1 I039_1162(w_039_1162, w_009_020);
  nand2 I039_1213(w_039_1213, w_018_170, w_022_175);
  nand2 I039_1227(w_039_1227, w_014_316, w_006_192);
  not1 I039_1232(w_039_1232, w_004_1801);
  and2 I039_1235(w_039_1235, w_032_196, w_038_457);
  or2  I039_1273(w_039_1273, w_006_200, w_005_116);
  and2 I039_1280(w_039_1280, w_016_028, w_029_098);
  nand2 I039_1295(w_039_1295, w_001_1640, w_025_1508);
  or2  I039_1297(w_039_1297, w_033_539, w_004_1782);
  not1 I039_1308(w_039_1308, w_014_344);
  not1 I039_1311(w_039_1311, w_004_286);
  and2 I039_1335(w_039_1335, w_000_1345, w_036_1289);
  or2  I039_1361(w_039_1361, w_011_290, w_007_550);
  nand2 I039_1362(w_039_1362, w_001_603, w_025_1170);
  nand2 I039_1372(w_039_1372, w_000_607, w_004_1094);
  nand2 I039_1392(w_039_1392, w_026_1268, w_011_727);
  or2  I039_1407(w_039_1407, w_022_417, w_022_405);
  not1 I039_1446(w_039_1446, w_035_343);
  and2 I039_1457(w_039_1457, w_037_774, w_004_775);
  or2  I039_1470(w_039_1470, w_020_1068, w_021_023);
  not1 I039_1496(w_039_1496, w_031_270);
  not1 I039_1509(w_039_1509, w_026_1257);
  not1 I039_1530(w_039_1530, w_030_496);
  not1 I039_1548(w_039_1548, w_031_159);
  and2 I039_1551(w_039_1551, w_022_013, w_017_895);
  not1 I039_1577(w_039_1577, w_002_106);
  not1 I039_1582(w_039_1582, w_030_229);
  not1 I039_1588(w_039_1588, w_030_620);
  and2 I039_1597(w_039_1597, w_029_132, w_038_173);
  not1 I039_1600(w_039_1600, w_035_1720);
  or2  I039_1605(w_039_1605, w_002_281, w_036_033);
  not1 I039_1611(w_039_1611, w_006_185);
  not1 I039_1634(w_039_1634, w_028_029);
  and2 I039_1643(w_039_1643, w_022_188, w_005_131);
  not1 I039_1654(w_039_1654, w_000_489);
  and2 I039_1699(w_039_1699, w_037_765, w_036_1043);
  and2 I039_1726(w_039_1726, w_038_325, w_035_1303);
  not1 I039_1731(w_039_1731, w_008_184);
  not1 I039_1753(w_039_1753, w_013_169);
  and2 I039_1768(w_039_1768, w_029_274, w_001_229);
  not1 I039_1770(w_039_1770, w_007_1090);
  or2  I039_1788(w_039_1788, w_013_299, w_021_119);
  nand2 I039_1835(w_039_1835, w_007_247, w_013_283);
  or2  I039_1836(w_039_1836, w_026_219, w_027_067);
  or2  I039_1856(w_039_1856, w_038_302, w_026_440);
  nand2 I039_1869(w_039_1869, w_010_170, w_031_117);
  and2 I039_1890(w_039_1890, w_023_726, w_032_042);
  and2 I039_1891(w_039_1891, w_026_1094, w_014_438);
  nand2 I039_1906(w_039_1906, w_030_557, w_028_721);
  or2  I039_1907(w_039_1907, w_034_378, w_020_274);
  or2  I039_1919(w_039_1919, w_014_581, w_036_937);
  or2  I039_1932(w_039_1932, w_031_351, w_020_074);
  or2  I040_011(w_040_011, w_039_477, w_012_109);
  not1 I040_015(w_040_015, w_016_022);
  and2 I040_016(w_040_016, w_034_569, w_004_100);
  and2 I040_019(w_040_019, w_002_068, w_035_777);
  nand2 I040_020(w_040_020, w_023_1153, w_013_206);
  and2 I040_024(w_040_024, w_024_303, w_015_273);
  nand2 I040_030(w_040_030, w_021_060, w_026_588);
  not1 I040_037(w_040_037, w_038_109);
  and2 I040_044(w_040_044, w_026_144, w_027_237);
  not1 I040_048(w_040_048, w_007_207);
  not1 I040_052(w_040_052, w_001_1676);
  nand2 I040_055(w_040_055, w_008_491, w_008_278);
  not1 I040_056(w_040_056, w_023_216);
  not1 I040_059(w_040_059, w_006_194);
  nand2 I040_060(w_040_060, w_013_167, w_008_491);
  nand2 I040_061(w_040_061, w_031_389, w_012_075);
  and2 I040_068(w_040_068, w_002_228, w_019_189);
  and2 I040_075(w_040_075, w_012_599, w_021_080);
  not1 I040_080(w_040_080, w_013_137);
  or2  I040_086(w_040_086, w_029_180, w_030_837);
  not1 I040_093(w_040_093, w_027_347);
  or2  I040_096(w_040_096, w_008_277, w_004_1020);
  nand2 I040_102(w_040_102, w_023_091, w_016_028);
  not1 I040_121(w_040_121, w_035_1098);
  nand2 I040_127(w_040_127, w_031_102, w_030_315);
  nand2 I040_134(w_040_134, w_003_171, w_026_195);
  or2  I040_148(w_040_148, w_008_644, w_015_232);
  and2 I040_165(w_040_165, w_017_1165, w_036_1356);
  or2  I040_172(w_040_172, w_005_1347, w_018_146);
  and2 I040_183(w_040_183, w_029_090, w_016_034);
  nand2 I040_189(w_040_189, w_014_271, w_019_449);
  nand2 I040_203(w_040_203, w_023_882, w_003_248);
  not1 I040_208(w_040_208, w_028_067);
  and2 I040_210(w_040_210, w_030_174, w_003_104);
  or2  I040_212(w_040_212, w_006_271, w_039_1577);
  not1 I040_220(w_040_220, w_021_148);
  and2 I040_225(w_040_225, w_005_1574, w_036_1294);
  or2  I040_226(w_040_226, w_010_377, w_027_574);
  not1 I040_227(w_040_227, w_009_014);
  nand2 I040_239(w_040_239, w_015_076, w_026_1463);
  not1 I040_255(w_040_255, w_024_453);
  not1 I040_260(w_040_260, w_034_657);
  and2 I040_272(w_040_272, w_018_027, w_006_043);
  not1 I040_273(w_040_273, w_025_1042);
  and2 I040_278(w_040_278, w_017_1284, w_024_1408);
  and2 I040_294(w_040_294, w_021_104, w_024_542);
  nand2 I040_297(w_040_297, w_009_098, w_015_103);
  nand2 I040_306(w_040_306, w_002_457, w_010_235);
  not1 I040_307(w_040_307, w_029_227);
  nand2 I040_312(w_040_312, w_021_150, w_010_089);
  and2 I040_314(w_040_314, w_030_396, w_005_240);
  and2 I040_315(w_040_315, w_023_880, w_005_473);
  and2 I040_320(w_040_320, w_026_074, w_038_007);
  nand2 I040_323(w_040_323, w_035_1487, w_001_757);
  nand2 I040_324(w_040_324, w_031_350, w_004_1563);
  or2  I040_325(w_040_325, w_000_734, w_033_602);
  nand2 I040_333(w_040_333, w_033_1405, w_001_853);
  nand2 I040_353(w_040_353, w_036_803, w_019_303);
  and2 I040_356(w_040_356, w_023_347, w_016_035);
  or2  I040_364(w_040_364, w_038_019, w_019_879);
  or2  I040_365(w_040_365, w_027_211, w_011_640);
  and2 I040_380(w_040_380, w_001_288, w_019_445);
  or2  I040_387(w_040_387, w_012_034, w_004_510);
  or2  I040_390(w_040_390, w_032_003, w_001_210);
  and2 I040_407(w_040_407, w_012_129, w_013_265);
  nand2 I040_411(w_040_411, w_007_451, w_011_014);
  or2  I040_423(w_040_423, w_003_304, w_015_078);
  and2 I040_427(w_040_427, w_001_140, w_018_251);
  and2 I040_436(w_040_436, w_008_147, w_009_075);
  and2 I040_447(w_040_447, w_017_687, w_029_149);
  or2  I040_461(w_040_461, w_022_225, w_017_960);
  or2  I040_462(w_040_462, w_035_1198, w_028_092);
  or2  I040_463(w_040_463, w_038_007, w_005_123);
  and2 I040_468(w_040_468, w_016_016, w_033_803);
  nand2 I040_472(w_040_472, w_000_347, w_037_188);
  nand2 I040_473(w_040_473, w_031_676, w_010_154);
  and2 I040_482(w_040_482, w_021_227, w_000_796);
  nand2 I040_489(w_040_489, w_013_018, w_017_1666);
  or2  I040_495(w_040_495, w_034_607, w_020_355);
  and2 I040_512(w_040_512, w_024_1001, w_004_000);
  and2 I040_521(w_040_521, w_008_511, w_034_225);
  not1 I040_526(w_040_526, w_002_247);
  and2 I040_527(w_040_527, w_001_1441, w_020_516);
  or2  I040_539(w_040_539, w_039_726, w_009_083);
  or2  I040_568(w_040_568, w_006_026, w_034_412);
  nand2 I040_577(w_040_577, w_024_301, w_023_1363);
  and2 I040_583(w_040_583, w_006_198, w_015_106);
  nand2 I040_585(w_040_585, w_025_1041, w_029_148);
  nand2 I040_590(w_040_590, w_016_005, w_031_634);
  not1 I040_593(w_040_593, w_019_368);
  nand2 I040_632(w_040_632, w_008_858, w_013_185);
  not1 I040_663(w_040_663, w_028_082);
  not1 I040_667(w_040_667, w_017_1763);
  and2 I040_673(w_040_673, w_016_008, w_023_367);
  and2 I040_679(w_040_679, w_004_970, w_012_320);
  and2 I040_683(w_040_683, w_001_532, w_033_260);
  and2 I040_695(w_040_695, w_031_645, w_025_1169);
  or2  I040_700(w_040_700, w_002_185, w_024_1193);
  and2 I040_724(w_040_724, w_035_671, w_005_1592);
  or2  I040_729(w_040_729, w_021_124, w_002_405);
  not1 I040_737(w_040_737, w_023_123);
  or2  I040_754(w_040_754, w_024_539, w_004_1765);
  not1 I040_757(w_040_757, w_010_078);
  and2 I040_759(w_040_759, w_017_722, w_021_172);
  and2 I040_764(w_040_764, w_025_235, w_000_1622);
  and2 I040_766(w_040_766, w_011_147, w_018_249);
  not1 I040_770(w_040_770, w_031_1027);
  not1 I040_771(w_040_771, w_031_1001);
  or2  I040_791(w_040_791, w_018_194, w_009_055);
  nand2 I040_813(w_040_813, w_036_151, w_022_066);
  and2 I040_823(w_040_823, w_012_453, w_039_759);
  not1 I040_832(w_040_832, w_021_144);
  and2 I040_848(w_040_848, w_003_122, w_007_1101);
  and2 I040_852(w_040_852, w_022_001, w_013_036);
  and2 I040_854(w_040_854, w_035_029, w_023_345);
  nand2 I040_856(w_040_856, w_005_1015, w_024_092);
  not1 I040_869(w_040_869, w_026_1084);
  not1 I040_904(w_040_904, w_010_029);
  nand2 I040_911(w_040_911, w_028_258, w_006_038);
  not1 I040_914(w_040_914, w_026_654);
  not1 I040_938(w_040_938, w_025_1126);
  not1 I040_959(w_040_959, w_023_1090);
  and2 I040_978(w_040_978, w_005_167, w_005_1329);
  and2 I040_979(w_040_979, w_035_328, w_027_323);
  or2  I040_981(w_040_981, w_024_009, w_029_1006);
  and2 I040_984(w_040_984, w_004_828, w_036_281);
  nand2 I040_987(w_040_987, w_017_203, w_032_051);
  and2 I040_1003(w_040_1003, w_013_003, w_003_239);
  not1 I040_1005(w_040_1005, w_026_045);
  not1 I040_1013(w_040_1013, w_015_177);
  nand2 I040_1028(w_040_1028, w_027_220, w_018_228);
  and2 I040_1038(w_040_1038, w_023_1156, w_013_105);
  and2 I040_1046(w_040_1046, w_011_862, w_001_1207);
  or2  I040_1076(w_040_1076, w_001_1507, w_009_028);
  and2 I040_1082(w_040_1082, w_038_186, w_035_076);
  nand2 I040_1084(w_040_1084, w_037_303, w_026_998);
  and2 I040_1102(w_040_1102, w_031_645, w_014_333);
  not1 I040_1119(w_040_1119, w_018_246);
  and2 I040_1125(w_040_1125, w_006_034, w_002_262);
  and2 I040_1134(w_040_1134, w_002_526, w_000_798);
  not1 I040_1138(w_040_1138, w_010_076);
  and2 I040_1156(w_040_1156, w_029_1245, w_030_533);
  not1 I040_1178(w_040_1178, w_012_100);
  nand2 I040_1195(w_040_1195, w_032_231, w_036_728);
  and2 I040_1213(w_040_1213, w_020_277, w_022_023);
  not1 I040_1232(w_040_1232, w_035_144);
  not1 I040_1237(w_040_1237, w_031_937);
  not1 I040_1263(w_040_1263, w_007_159);
  and2 I040_1276(w_040_1276, w_032_138, w_025_300);
  nand2 I040_1286(w_040_1286, w_006_026, w_027_280);
  nand2 I040_1291(w_040_1291, w_033_1643, w_036_505);
  and2 I040_1294(w_040_1294, w_004_1807, w_035_104);
  not1 I040_1304(w_040_1304, w_032_194);
  nand2 I040_1314(w_040_1314, w_020_722, w_034_511);
  and2 I040_1320(w_040_1320, w_025_552, w_023_1318);
  nand2 I040_1327(w_040_1327, w_039_1530, w_029_142);
  or2  I040_1350(w_040_1350, w_029_985, w_034_309);
  not1 I040_1352(w_040_1352, w_000_1647);
  or2  I040_1383(w_040_1383, w_029_319, w_000_809);
  or2  I041_002(w_041_002, w_031_770, w_026_609);
  not1 I041_004(w_041_004, w_030_435);
  or2  I041_007(w_041_007, w_010_221, w_015_278);
  nand2 I041_008(w_041_008, w_039_415, w_020_369);
  nand2 I041_010(w_041_010, w_013_072, w_038_338);
  not1 I041_012(w_041_012, w_022_032);
  and2 I041_017(w_041_017, w_030_613, w_032_009);
  not1 I041_018(w_041_018, w_023_748);
  or2  I041_021(w_041_021, w_030_042, w_018_227);
  or2  I041_022(w_041_022, w_035_1530, w_028_083);
  and2 I041_025(w_041_025, w_028_084, w_018_234);
  and2 I041_026(w_041_026, w_028_757, w_007_062);
  not1 I041_035(w_041_035, w_014_334);
  or2  I041_037(w_041_037, w_021_139, w_004_535);
  not1 I041_042(w_041_042, w_002_256);
  nand2 I041_043(w_041_043, w_022_354, w_035_1054);
  not1 I041_044(w_041_044, w_040_468);
  and2 I041_045(w_041_045, w_013_338, w_032_072);
  nand2 I041_049(w_041_049, w_028_580, w_027_006);
  not1 I041_052(w_041_052, w_000_395);
  not1 I041_053(w_041_053, w_006_322);
  nand2 I041_055(w_041_055, w_024_017, w_021_130);
  or2  I041_059(w_041_059, w_003_061, w_033_276);
  or2  I041_062(w_041_062, w_018_030, w_040_1294);
  and2 I041_063(w_041_063, w_030_789, w_005_1398);
  nand2 I041_064(w_041_064, w_015_171, w_020_620);
  and2 I041_065(w_041_065, w_029_311, w_018_085);
  not1 I041_066(w_041_066, w_010_230);
  nand2 I041_069(w_041_069, w_025_1265, w_039_1446);
  or2  I041_071(w_041_071, w_029_1087, w_011_140);
  and2 I041_073(w_041_073, w_040_255, w_017_003);
  nand2 I041_074(w_041_074, w_030_105, w_022_391);
  not1 I041_077(w_041_077, w_036_657);
  or2  I041_081(w_041_081, w_034_116, w_031_485);
  not1 I041_082(w_041_082, w_011_512);
  not1 I041_084(w_041_084, w_038_148);
  nand2 I041_085(w_041_085, w_029_245, w_009_086);
  and2 I041_087(w_041_087, w_027_531, w_013_302);
  or2  I041_090(w_041_090, w_003_190, w_036_1325);
  and2 I041_091(w_041_091, w_035_225, w_019_480);
  and2 I041_092(w_041_092, w_028_470, w_005_1171);
  or2  I041_096(w_041_096, w_023_013, w_040_423);
  or2  I041_098(w_041_098, w_020_397, w_022_172);
  not1 I041_107(w_041_107, w_036_1227);
  and2 I041_108(w_041_108, w_030_840, w_014_366);
  nand2 I041_110(w_041_110, w_016_026, w_026_352);
  nand2 I041_111(w_041_111, w_024_415, w_033_1305);
  nand2 I041_113(w_041_113, w_014_704, w_006_212);
  nand2 I041_114(w_041_114, w_014_691, w_002_276);
  or2  I041_115(w_041_115, w_004_644, w_029_475);
  or2  I041_118(w_041_118, w_021_141, w_033_127);
  not1 I041_121(w_041_121, w_010_149);
  not1 I041_122(w_041_122, w_040_1232);
  or2  I041_124(w_041_124, w_003_034, w_003_287);
  or2  I041_126(w_041_126, w_008_186, w_001_421);
  nand2 I041_127(w_041_127, w_017_1679, w_038_043);
  nand2 I041_128(w_041_128, w_031_853, w_038_366);
  nand2 I041_131(w_041_131, w_022_056, w_035_138);
  nand2 I041_132(w_041_132, w_038_224, w_028_088);
  or2  I041_134(w_041_134, w_005_901, w_000_110);
  not1 I041_140(w_041_140, w_031_300);
  nand2 I041_146(w_041_146, w_016_034, w_019_659);
  or2  I041_149(w_041_149, w_022_036, w_034_144);
  or2  I041_150(w_041_150, w_036_029, w_000_645);
  and2 I041_152(w_041_152, w_013_234, w_037_669);
  and2 I041_154(w_041_154, w_022_286, w_003_008);
  and2 I041_155(w_041_155, w_003_230, w_025_1374);
  nand2 I041_156(w_041_156, w_019_153, w_025_173);
  nand2 I041_157(w_041_157, w_025_527, w_025_959);
  not1 I041_158(w_041_158, w_030_780);
  and2 I041_161(w_041_161, w_002_312, w_001_877);
  or2  I041_169(w_041_169, w_005_097, w_014_673);
  nand2 I041_171(w_041_171, w_001_151, w_025_1472);
  nand2 I041_178(w_041_178, w_017_1379, w_036_180);
  nand2 I041_180(w_041_180, w_003_148, w_009_072);
  and2 I041_181(w_041_181, w_040_667, w_011_173);
  or2  I041_183(w_041_183, w_040_210, w_027_207);
  nand2 I041_186(w_041_186, w_028_725, w_040_278);
  or2  I041_187(w_041_187, w_005_1076, w_036_133);
  or2  I041_188(w_041_188, w_030_344, w_040_527);
  or2  I041_191(w_041_191, w_019_302, w_018_186);
  or2  I041_193(w_041_193, w_038_039, w_038_335);
  and2 I041_194(w_041_194, w_006_173, w_023_191);
  nand2 I041_197(w_041_197, w_000_1082, w_035_1016);
  or2  I041_198(w_041_198, w_023_114, w_009_012);
  and2 I041_199(w_041_199, w_008_666, w_035_1506);
  not1 I041_200(w_041_200, w_012_228);
  and2 I041_201(w_041_201, w_036_255, w_002_215);
  not1 I041_202(w_041_202, w_027_120);
  and2 I041_204(w_041_204, w_037_1343, w_030_385);
  and2 I041_205(w_041_205, w_009_096, w_032_197);
  and2 I041_206(w_041_206, w_011_576, w_023_347);
  and2 I041_207(w_041_207, w_028_258, w_027_059);
  nand2 I041_208(w_041_208, w_024_166, w_006_225);
  or2  I041_211(w_041_211, w_013_221, w_037_702);
  or2  I041_212(w_041_212, w_030_614, w_023_1357);
  and2 I041_217(w_041_217, w_002_125, w_018_220);
  and2 I041_219(w_041_219, w_017_1223, w_025_824);
  and2 I041_229(w_041_229, w_014_487, w_008_018);
  and2 I041_230(w_041_230, w_008_243, w_027_174);
  and2 I041_231(w_041_231, w_000_767, w_001_1489);
  not1 I041_232(w_041_232, w_005_134);
  not1 I041_235(w_041_235, w_027_553);
  or2  I041_237(w_041_237, w_032_027, w_025_565);
  nand2 I041_245(w_041_245, w_027_560, w_014_118);
  nand2 I041_246(w_041_246, w_015_188, w_017_1655);
  nand2 I041_247(w_041_247, w_013_101, w_028_298);
  not1 I041_248(w_041_248, w_010_101);
  not1 I041_249(w_041_249, w_005_1139);
  nand2 I041_250(w_041_250, w_012_213, w_008_429);
  nand2 I041_253(w_041_253, w_025_434, w_032_067);
  nand2 I041_254(w_041_254, w_005_1554, w_024_1638);
  nand2 I041_257(w_041_257, w_013_067, w_014_324);
  not1 I041_258(w_041_258, w_013_247);
  nand2 I041_264(w_041_264, w_016_001, w_022_098);
  and2 I041_265(w_041_265, w_002_178, w_035_091);
  and2 I041_267(w_041_267, w_017_1373, w_038_404);
  and2 I041_268(w_041_268, w_027_079, w_003_167);
  or2  I041_271(w_041_271, w_037_1000, w_001_980);
  not1 I041_273(w_041_273, w_040_1350);
  nand2 I041_275(w_041_275, w_036_323, w_010_351);
  and2 I041_278(w_041_278, w_023_238, w_017_649);
  not1 I041_279(w_041_279, w_021_015);
  and2 I041_282(w_041_282, w_033_012, w_005_736);
  not1 I041_285(w_041_285, w_029_567);
  not1 I041_288(w_041_288, w_031_934);
  not1 I041_289(w_041_289, w_026_610);
  nand2 I041_294(w_041_294, w_009_062, w_016_000);
  not1 I042_000(w_042_000, w_025_064);
  nand2 I042_001(w_042_001, w_031_040, w_003_316);
  not1 I042_002(w_042_002, w_008_597);
  and2 I042_003(w_042_003, w_012_199, w_015_137);
  or2  I042_007(w_042_007, w_027_472, w_034_442);
  and2 I042_008(w_042_008, w_035_1079, w_006_098);
  or2  I042_009(w_042_009, w_012_628, w_008_773);
  not1 I042_014(w_042_014, w_011_037);
  and2 I042_016(w_042_016, w_004_009, w_010_230);
  or2  I042_017(w_042_017, w_036_1464, w_009_111);
  and2 I042_018(w_042_018, w_031_296, w_005_068);
  or2  I042_019(w_042_019, w_031_712, w_015_184);
  and2 I042_021(w_042_021, w_011_846, w_008_785);
  not1 I042_022(w_042_022, w_006_028);
  nand2 I042_023(w_042_023, w_017_1670, w_040_059);
  not1 I042_025(w_042_025, w_039_1788);
  and2 I042_026(w_042_026, w_022_353, w_017_346);
  or2  I042_027(w_042_027, w_022_320, w_039_676);
  not1 I042_028(w_042_028, w_010_238);
  nand2 I042_029(w_042_029, w_008_018, w_014_752);
  not1 I042_030(w_042_030, w_030_191);
  nand2 I042_031(w_042_031, w_019_583, w_022_088);
  nand2 I042_034(w_042_034, w_027_371, w_003_148);
  or2  I042_035(w_042_035, w_013_301, w_004_032);
  and2 I042_036(w_042_036, w_017_1882, w_004_1829);
  not1 I042_037(w_042_037, w_017_100);
  not1 I042_040(w_042_040, w_021_238);
  nand2 I042_041(w_042_041, w_040_208, w_031_356);
  nand2 I042_044(w_042_044, w_005_1283, w_036_513);
  not1 I042_046(w_042_046, w_011_217);
  not1 I042_047(w_042_047, w_029_1135);
  or2  I042_048(w_042_048, w_018_222, w_008_253);
  and2 I042_051(w_042_051, w_003_304, w_029_146);
  and2 I042_052(w_042_052, w_002_183, w_004_085);
  or2  I042_053(w_042_053, w_016_031, w_026_127);
  or2  I042_054(w_042_054, w_035_1037, w_005_039);
  nand2 I042_055(w_042_055, w_015_211, w_036_369);
  nand2 I042_058(w_042_058, w_013_154, w_030_454);
  nand2 I042_060(w_042_060, w_032_106, w_009_013);
  and2 I042_062(w_042_062, w_019_965, w_004_537);
  or2  I042_063(w_042_063, w_031_228, w_010_397);
  and2 I042_064(w_042_064, w_029_251, w_030_147);
  or2  I042_065(w_042_065, w_035_1176, w_037_438);
  and2 I042_068(w_042_068, w_003_255, w_040_226);
  not1 I042_072(w_042_072, w_034_471);
  not1 I042_073(w_042_073, w_019_864);
  nand2 I042_074(w_042_074, w_011_574, w_034_347);
  nand2 I042_076(w_042_076, w_012_471, w_041_090);
  or2  I042_077(w_042_077, w_029_567, w_020_476);
  and2 I042_079(w_042_079, w_030_830, w_016_014);
  not1 I042_081(w_042_081, w_024_1137);
  and2 I042_084(w_042_084, w_019_025, w_000_614);
  not1 I042_085(w_042_085, w_025_711);
  not1 I042_086(w_042_086, w_012_557);
  or2  I042_088(w_042_088, w_035_1518, w_029_496);
  not1 I042_089(w_042_089, w_003_005);
  and2 I042_093(w_042_093, w_035_051, w_004_328);
  nand2 I042_094(w_042_094, w_006_026, w_038_300);
  and2 I042_095(w_042_095, w_029_802, w_029_308);
  or2  I042_096(w_042_096, w_033_249, w_021_231);
  not1 I042_097(w_042_097, w_038_084);
  not1 I042_100(w_042_100, w_034_475);
  nand2 I042_102(w_042_102, w_026_1243, w_027_102);
  or2  I042_103(w_042_103, w_005_1499, w_024_250);
  not1 I042_104(w_042_104, w_003_102);
  and2 I042_105(w_042_105, w_009_042, w_009_076);
  and2 I042_107(w_042_107, w_009_049, w_027_114);
  or2  I042_109(w_042_109, w_003_229, w_024_934);
  or2  I042_110(w_042_110, w_006_154, w_013_013);
  and2 I042_111(w_042_111, w_024_1576, w_008_058);
  and2 I042_112(w_042_112, w_025_649, w_014_430);
  nand2 I042_113(w_042_113, w_013_112, w_007_546);
  and2 I042_115(w_042_115, w_041_248, w_004_1656);
  nand2 I042_117(w_042_117, w_033_112, w_034_664);
  and2 I042_118(w_042_118, w_016_007, w_004_1698);
  or2  I042_119(w_042_119, w_030_699, w_024_316);
  or2  I042_121(w_042_121, w_039_167, w_039_259);
  nand2 I042_122(w_042_122, w_041_127, w_013_116);
  not1 I042_124(w_042_124, w_027_587);
  nand2 I042_125(w_042_125, w_041_066, w_041_183);
  not1 I042_127(w_042_127, w_016_024);
  or2  I042_128(w_042_128, w_010_090, w_040_683);
  nand2 I042_129(w_042_129, w_007_373, w_040_1213);
  and2 I042_130(w_042_130, w_036_322, w_012_392);
  or2  I042_132(w_042_132, w_025_823, w_025_1675);
  and2 I042_134(w_042_134, w_028_041, w_004_1047);
  not1 I042_135(w_042_135, w_003_000);
  and2 I042_137(w_042_137, w_016_033, w_035_208);
  not1 I042_139(w_042_139, w_031_743);
  and2 I042_140(w_042_140, w_041_275, w_039_614);
  or2  I042_141(w_042_141, w_024_473, w_039_1059);
  nand2 I042_142(w_042_142, w_001_659, w_015_119);
  and2 I043_000(w_043_000, w_032_148, w_021_260);
  nand2 I043_001(w_043_001, w_041_247, w_032_187);
  and2 I043_004(w_043_004, w_010_156, w_031_429);
  and2 I043_005(w_043_005, w_021_256, w_036_218);
  or2  I043_006(w_043_006, w_003_061, w_018_064);
  not1 I043_010(w_043_010, w_029_747);
  or2  I043_011(w_043_011, w_010_239, w_041_132);
  or2  I043_012(w_043_012, w_026_446, w_005_1415);
  and2 I043_013(w_043_013, w_015_103, w_039_648);
  or2  I043_014(w_043_014, w_032_169, w_028_583);
  and2 I043_015(w_043_015, w_004_1157, w_000_1811);
  and2 I043_016(w_043_016, w_027_578, w_006_173);
  and2 I043_019(w_043_019, w_041_294, w_004_1534);
  not1 I043_020(w_043_020, w_013_211);
  or2  I043_021(w_043_021, w_034_166, w_018_134);
  and2 I043_022(w_043_022, w_018_015, w_041_063);
  not1 I043_023(w_043_023, w_039_879);
  nand2 I043_024(w_043_024, w_011_298, w_036_170);
  not1 I043_025(w_043_025, w_041_264);
  or2  I043_026(w_043_026, w_008_370, w_032_176);
  and2 I043_027(w_043_027, w_019_485, w_008_332);
  not1 I043_028(w_043_028, w_042_068);
  and2 I043_029(w_043_029, w_030_182, w_023_357);
  and2 I043_030(w_043_030, w_018_104, w_016_003);
  and2 I043_031(w_043_031, w_019_1057, w_018_176);
  and2 I043_032(w_043_032, w_016_018, w_020_483);
  nand2 I043_034(w_043_034, w_033_320, w_028_863);
  and2 I043_035(w_043_035, w_033_1235, w_023_1608);
  not1 I043_036(w_043_036, w_034_252);
  nand2 I043_037(w_043_037, w_042_127, w_030_224);
  nand2 I043_039(w_043_039, w_006_274, w_013_046);
  and2 I043_040(w_043_040, w_030_362, w_036_374);
  and2 I043_041(w_043_041, w_022_059, w_005_1674);
  or2  I043_042(w_043_042, w_028_373, w_039_933);
  not1 I043_043(w_043_043, w_001_585);
  not1 I043_046(w_043_046, w_020_806);
  nand2 I043_048(w_043_048, w_040_695, w_024_282);
  or2  I043_049(w_043_049, w_002_134, w_025_137);
  nand2 I043_050(w_043_050, w_019_722, w_040_764);
  and2 I043_051(w_043_051, w_007_045, w_029_541);
  or2  I043_052(w_043_052, w_036_101, w_016_006);
  nand2 I043_053(w_043_053, w_041_154, w_009_025);
  or2  I043_054(w_043_054, w_028_553, w_040_904);
  nand2 I043_055(w_043_055, w_018_108, w_012_274);
  or2  I043_056(w_043_056, w_000_905, w_027_243);
  not1 I043_057(w_043_057, w_032_201);
  nand2 I043_058(w_043_058, w_010_321, w_009_093);
  nand2 I043_059(w_043_059, w_017_723, w_029_070);
  and2 I043_060(w_043_060, w_039_1361, w_024_944);
  or2  I043_062(w_043_062, w_031_308, w_023_1371);
  or2  I043_063(w_043_063, w_015_276, w_009_106);
  not1 I043_064(w_043_064, w_033_1444);
  not1 I043_065(w_043_065, w_000_186);
  nand2 I043_066(w_043_066, w_038_390, w_021_259);
  and2 I043_067(w_043_067, w_028_546, w_017_753);
  and2 I043_068(w_043_068, w_034_328, w_007_097);
  nand2 I043_070(w_043_070, w_001_281, w_041_246);
  or2  I043_071(w_043_071, w_023_1180, w_032_234);
  not1 I043_073(w_043_073, w_022_142);
  and2 I043_075(w_043_075, w_004_1812, w_016_012);
  not1 I043_077(w_043_077, w_038_201);
  not1 I043_078(w_043_078, w_028_054);
  and2 I043_079(w_043_079, w_006_222, w_024_066);
  and2 I043_081(w_043_081, w_005_917, w_011_594);
  nand2 I043_082(w_043_082, w_034_630, w_022_169);
  nand2 I043_083(w_043_083, w_006_296, w_037_1050);
  not1 I043_084(w_043_084, w_024_095);
  or2  I043_085(w_043_085, w_010_147, w_022_030);
  or2  I043_088(w_043_088, w_033_053, w_011_872);
  nand2 I043_089(w_043_089, w_025_1242, w_006_023);
  and2 I043_091(w_043_091, w_024_1504, w_019_290);
  nand2 I043_092(w_043_092, w_018_255, w_034_130);
  nand2 I043_093(w_043_093, w_033_355, w_037_604);
  nand2 I043_094(w_043_094, w_022_161, w_003_163);
  and2 I043_095(w_043_095, w_001_1123, w_015_151);
  not1 I043_096(w_043_096, w_018_255);
  nand2 I043_097(w_043_097, w_014_013, w_032_233);
  or2  I043_098(w_043_098, w_008_760, w_038_122);
  or2  I043_099(w_043_099, w_021_002, w_023_190);
  and2 I043_100(w_043_100, w_009_077, w_041_146);
  and2 I043_101(w_043_101, w_036_781, w_018_132);
  and2 I043_102(w_043_102, w_026_172, w_038_304);
  and2 I043_103(w_043_103, w_029_999, w_020_897);
  not1 I043_105(w_043_105, w_014_524);
  nand2 I044_018(w_044_018, w_043_041, w_025_031);
  nand2 I044_022(w_044_022, w_006_020, w_028_175);
  not1 I044_030(w_044_030, w_005_1370);
  and2 I044_033(w_044_033, w_024_1250, w_023_290);
  or2  I044_035(w_044_035, w_009_067, w_020_358);
  nand2 I044_047(w_044_047, w_002_113, w_010_246);
  and2 I044_056(w_044_056, w_017_1665, w_022_041);
  nand2 I044_074(w_044_074, w_026_882, w_037_210);
  nand2 I044_087(w_044_087, w_000_178, w_030_774);
  or2  I044_107(w_044_107, w_014_516, w_028_731);
  or2  I044_112(w_044_112, w_009_082, w_002_082);
  and2 I044_115(w_044_115, w_001_067, w_031_985);
  nand2 I044_129(w_044_129, w_001_449, w_020_631);
  and2 I044_132(w_044_132, w_026_1489, w_021_232);
  and2 I044_134(w_044_134, w_041_232, w_037_145);
  and2 I044_137(w_044_137, w_038_007, w_020_154);
  or2  I044_142(w_044_142, w_006_077, w_017_408);
  nand2 I044_147(w_044_147, w_018_135, w_032_241);
  nand2 I044_156(w_044_156, w_034_578, w_010_103);
  and2 I044_166(w_044_166, w_002_138, w_015_217);
  not1 I044_175(w_044_175, w_038_384);
  or2  I044_176(w_044_176, w_032_001, w_011_412);
  nand2 I044_184(w_044_184, w_029_468, w_004_171);
  not1 I044_189(w_044_189, w_027_356);
  and2 I044_196(w_044_196, w_021_216, w_017_871);
  or2  I044_199(w_044_199, w_030_196, w_009_032);
  or2  I044_201(w_044_201, w_029_244, w_019_770);
  not1 I044_226(w_044_226, w_007_638);
  and2 I044_264(w_044_264, w_025_097, w_037_1329);
  or2  I044_308(w_044_308, w_009_059, w_012_066);
  nand2 I044_309(w_044_309, w_002_018, w_003_059);
  nand2 I044_314(w_044_314, w_021_205, w_024_1187);
  nand2 I044_324(w_044_324, w_022_108, w_022_171);
  or2  I044_342(w_044_342, w_013_242, w_029_281);
  nand2 I044_355(w_044_355, w_002_342, w_033_276);
  nand2 I044_357(w_044_357, w_016_024, w_036_1239);
  not1 I044_374(w_044_374, w_036_1320);
  not1 I044_390(w_044_390, w_023_289);
  not1 I044_393(w_044_393, w_014_457);
  and2 I044_414(w_044_414, w_018_271, w_036_697);
  not1 I044_443(w_044_443, w_032_053);
  or2  I044_462(w_044_462, w_037_633, w_013_266);
  or2  I044_465(w_044_465, w_035_1107, w_028_809);
  nand2 I044_466(w_044_466, w_019_613, w_008_651);
  or2  I044_475(w_044_475, w_022_235, w_000_631);
  or2  I044_538(w_044_538, w_028_469, w_024_262);
  and2 I044_541(w_044_541, w_030_826, w_026_820);
  nand2 I044_542(w_044_542, w_026_1177, w_030_774);
  nand2 I044_569(w_044_569, w_016_013, w_027_076);
  and2 I044_607(w_044_607, w_032_042, w_016_000);
  and2 I044_613(w_044_613, w_031_409, w_037_804);
  not1 I044_618(w_044_618, w_002_106);
  or2  I044_665(w_044_665, w_005_409, w_005_162);
  nand2 I044_675(w_044_675, w_000_1511, w_038_077);
  or2  I044_682(w_044_682, w_005_1168, w_017_1636);
  or2  I044_697(w_044_697, w_017_117, w_022_140);
  not1 I044_718(w_044_718, w_043_030);
  nand2 I044_724(w_044_724, w_008_128, w_026_233);
  and2 I044_764(w_044_764, w_017_1201, w_043_000);
  nand2 I044_777(w_044_777, w_016_031, w_013_072);
  nand2 I044_778(w_044_778, w_022_156, w_004_1787);
  not1 I044_784(w_044_784, w_038_332);
  or2  I044_788(w_044_788, w_000_1356, w_029_163);
  and2 I044_790(w_044_790, w_019_239, w_022_286);
  and2 I044_791(w_044_791, w_015_195, w_032_138);
  and2 I044_794(w_044_794, w_025_547, w_037_1343);
  and2 I044_795(w_044_795, w_013_022, w_019_842);
  not1 I044_831(w_044_831, w_031_425);
  nand2 I044_870(w_044_870, w_043_048, w_035_1273);
  and2 I044_897(w_044_897, w_013_159, w_016_034);
  and2 I044_907(w_044_907, w_004_770, w_029_106);
  or2  I044_908(w_044_908, w_035_1119, w_040_771);
  nand2 I044_913(w_044_913, w_040_1327, w_041_197);
  or2  I044_914(w_044_914, w_018_211, w_008_174);
  or2  I044_931(w_044_931, w_034_090, w_015_283);
  not1 I044_951(w_044_951, w_029_533);
  nand2 I044_954(w_044_954, w_013_068, w_012_298);
  nand2 I044_963(w_044_963, w_025_1004, w_010_372);
  or2  I044_972(w_044_972, w_001_052, w_022_194);
  and2 I044_990(w_044_990, w_001_1661, w_038_429);
  or2  I044_1077(w_044_1077, w_039_1235, w_011_184);
  not1 I044_1093(w_044_1093, w_021_265);
  or2  I044_1095(w_044_1095, w_003_138, w_018_249);
  and2 I044_1108(w_044_1108, w_020_164, w_012_536);
  or2  I044_1116(w_044_1116, w_039_631, w_033_708);
  not1 I044_1117(w_044_1117, w_014_491);
  not1 I044_1134(w_044_1134, w_020_934);
  or2  I044_1139(w_044_1139, w_015_161, w_041_268);
  or2  I044_1141(w_044_1141, w_036_1226, w_014_574);
  and2 I044_1146(w_044_1146, w_042_097, w_013_053);
  nand2 I044_1152(w_044_1152, w_030_723, w_040_436);
  or2  I044_1176(w_044_1176, w_013_192, w_010_163);
  nand2 I044_1197(w_044_1197, w_038_161, w_022_208);
  nand2 I044_1209(w_044_1209, w_035_722, w_033_115);
  not1 I044_1217(w_044_1217, w_016_024);
  nand2 I044_1224(w_044_1224, w_000_286, w_018_012);
  nand2 I044_1230(w_044_1230, w_020_949, w_038_429);
  nand2 I044_1251(w_044_1251, w_043_067, w_036_525);
  nand2 I044_1261(w_044_1261, w_027_550, w_028_880);
  nand2 I044_1268(w_044_1268, w_031_480, w_011_879);
  and2 I044_1274(w_044_1274, w_016_033, w_032_239);
  not1 I044_1327(w_044_1327, w_028_095);
  or2  I044_1330(w_044_1330, w_038_048, w_043_056);
  not1 I044_1342(w_044_1342, w_024_032);
  nand2 I044_1344(w_044_1344, w_026_331, w_042_007);
  nand2 I044_1377(w_044_1377, w_027_523, w_029_135);
  not1 I044_1379(w_044_1379, w_013_084);
  and2 I044_1383(w_044_1383, w_042_021, w_023_232);
  and2 I044_1386(w_044_1386, w_013_175, w_038_337);
  or2  I044_1405(w_044_1405, w_017_381, w_042_060);
  or2  I044_1417(w_044_1417, w_012_406, w_000_479);
  nand2 I044_1426(w_044_1426, w_041_071, w_002_453);
  or2  I044_1427(w_044_1427, w_028_170, w_012_666);
  and2 I044_1446(w_044_1446, w_018_072, w_041_134);
  and2 I044_1447(w_044_1447, w_037_363, w_007_676);
  or2  I044_1459(w_044_1459, w_026_330, w_043_048);
  and2 I044_1465(w_044_1465, w_013_123, w_009_102);
  or2  I044_1481(w_044_1481, w_030_229, w_038_136);
  and2 I044_1505(w_044_1505, w_023_334, w_018_227);
  nand2 I044_1523(w_044_1523, w_015_032, w_005_014);
  or2  I044_1550(w_044_1550, w_010_415, w_012_257);
  or2  I044_1566(w_044_1566, w_038_227, w_017_846);
  or2  I044_1580(w_044_1580, w_007_1566, w_017_540);
  and2 I044_1614(w_044_1614, w_041_049, w_006_140);
  not1 I044_1616(w_044_1616, w_019_326);
  or2  I044_1629(w_044_1629, w_013_272, w_030_769);
  or2  I044_1630(w_044_1630, w_031_564, w_009_062);
  not1 I044_1635(w_044_1635, w_030_757);
  not1 I044_1639(w_044_1639, w_007_1379);
  not1 I044_1684(w_044_1684, w_026_119);
  or2  I044_1690(w_044_1690, w_005_319, w_033_1624);
  nand2 I044_1695(w_044_1695, w_031_609, w_026_481);
  and2 I044_1723(w_044_1723, w_000_1178, w_007_823);
  nand2 I044_1750(w_044_1750, w_007_388, w_017_673);
  not1 I044_1751(w_044_1751, w_032_021);
  and2 I044_1752(w_044_1752, w_008_036, w_041_268);
  not1 I044_1769(w_044_1769, w_024_200);
  or2  I044_1781(w_044_1781, w_035_712, w_027_322);
  nand2 I044_1783(w_044_1783, w_035_1713, w_009_101);
  or2  I044_1792(w_044_1792, w_033_1268, w_014_032);
  not1 I045_005(w_045_005, w_024_290);
  or2  I045_009(w_045_009, w_026_1072, w_020_219);
  nand2 I045_023(w_045_023, w_030_050, w_015_268);
  nand2 I045_041(w_045_041, w_009_009, w_016_002);
  or2  I045_065(w_045_065, w_001_1207, w_000_1971);
  and2 I045_066(w_045_066, w_013_108, w_039_969);
  nand2 I045_070(w_045_070, w_033_114, w_012_607);
  not1 I045_072(w_045_072, w_028_780);
  and2 I045_077(w_045_077, w_009_052, w_033_123);
  or2  I045_082(w_045_082, w_005_1099, w_027_201);
  or2  I045_093(w_045_093, w_003_133, w_010_189);
  and2 I045_110(w_045_110, w_022_407, w_040_427);
  not1 I045_163(w_045_163, w_032_004);
  and2 I045_170(w_045_170, w_010_173, w_037_1106);
  or2  I045_171(w_045_171, w_002_441, w_003_091);
  not1 I045_199(w_045_199, w_005_759);
  or2  I045_209(w_045_209, w_011_076, w_030_783);
  or2  I045_213(w_045_213, w_040_911, w_015_244);
  or2  I045_224(w_045_224, w_013_024, w_020_457);
  or2  I045_226(w_045_226, w_034_511, w_027_001);
  and2 I045_251(w_045_251, w_000_474, w_000_422);
  not1 I045_255(w_045_255, w_017_385);
  or2  I045_266(w_045_266, w_039_490, w_031_184);
  nand2 I045_288(w_045_288, w_019_772, w_043_101);
  nand2 I045_290(w_045_290, w_016_035, w_023_836);
  nand2 I045_303(w_045_303, w_014_757, w_015_209);
  not1 I045_310(w_045_310, w_019_700);
  and2 I045_331(w_045_331, w_002_055, w_010_164);
  not1 I045_335(w_045_335, w_008_815);
  and2 I045_338(w_045_338, w_031_1025, w_005_622);
  or2  I045_344(w_045_344, w_025_352, w_015_038);
  nand2 I045_346(w_045_346, w_018_141, w_000_1311);
  or2  I045_365(w_045_365, w_017_1656, w_009_035);
  and2 I045_398(w_045_398, w_022_041, w_028_397);
  or2  I045_405(w_045_405, w_003_103, w_021_162);
  and2 I045_424(w_045_424, w_033_1001, w_002_158);
  nand2 I045_437(w_045_437, w_002_523, w_032_142);
  not1 I045_452(w_045_452, w_024_1544);
  not1 I045_475(w_045_475, w_014_271);
  nand2 I045_483(w_045_483, w_027_219, w_012_068);
  nand2 I045_490(w_045_490, w_025_435, w_000_865);
  and2 I045_495(w_045_495, w_001_619, w_012_628);
  nand2 I045_524(w_045_524, w_042_040, w_009_030);
  or2  I045_547(w_045_547, w_040_987, w_012_536);
  nand2 I045_548(w_045_548, w_040_134, w_026_276);
  nand2 I045_574(w_045_574, w_037_193, w_032_038);
  or2  I045_578(w_045_578, w_001_486, w_020_1001);
  nand2 I045_580(w_045_580, w_004_599, w_007_054);
  and2 I045_583(w_045_583, w_042_124, w_020_325);
  or2  I045_588(w_045_588, w_017_1666, w_008_184);
  nand2 I045_599(w_045_599, w_017_1870, w_034_551);
  nand2 I045_607(w_045_607, w_003_175, w_042_037);
  and2 I045_617(w_045_617, w_018_045, w_044_913);
  not1 I045_635(w_045_635, w_022_217);
  not1 I045_662(w_045_662, w_032_036);
  nand2 I045_666(w_045_666, w_013_174, w_000_559);
  and2 I045_710(w_045_710, w_008_577, w_003_289);
  or2  I045_711(w_045_711, w_010_037, w_026_449);
  or2  I045_721(w_045_721, w_030_048, w_035_323);
  nand2 I045_731(w_045_731, w_030_434, w_006_007);
  and2 I045_747(w_045_747, w_023_045, w_003_279);
  nand2 I045_752(w_045_752, w_018_255, w_033_391);
  nand2 I045_766(w_045_766, w_032_176, w_017_305);
  and2 I045_786(w_045_786, w_043_039, w_039_895);
  not1 I045_796(w_045_796, w_005_694);
  nand2 I045_802(w_045_802, w_013_073, w_006_133);
  and2 I045_805(w_045_805, w_027_580, w_019_000);
  and2 I045_830(w_045_830, w_036_148, w_011_854);
  or2  I045_874(w_045_874, w_004_162, w_033_1512);
  nand2 I045_937(w_045_937, w_009_069, w_015_147);
  and2 I045_957(w_045_957, w_012_100, w_008_172);
  nand2 I045_962(w_045_962, w_040_068, w_015_232);
  not1 I045_1002(w_045_1002, w_000_943);
  or2  I045_1015(w_045_1015, w_017_1238, w_012_425);
  and2 I045_1052(w_045_1052, w_038_175, w_007_044);
  and2 I045_1064(w_045_1064, w_026_1136, w_014_032);
  and2 I045_1066(w_045_1066, w_036_493, w_015_154);
  or2  I045_1071(w_045_1071, w_006_234, w_041_187);
  nand2 I045_1086(w_045_1086, w_031_963, w_006_032);
  not1 I045_1102(w_045_1102, w_043_100);
  and2 I045_1104(w_045_1104, w_013_214, w_041_085);
  or2  I045_1139(w_045_1139, w_044_1750, w_008_463);
  and2 I045_1153(w_045_1153, w_000_725, w_032_077);
  nand2 I045_1161(w_045_1161, w_006_006, w_020_585);
  not1 I045_1181(w_045_1181, w_008_553);
  nand2 I045_1189(w_045_1189, w_020_628, w_036_1217);
  nand2 I045_1203(w_045_1203, w_039_204, w_021_151);
  and2 I045_1229(w_045_1229, w_007_423, w_002_576);
  and2 I045_1231(w_045_1231, w_016_016, w_044_226);
  or2  I045_1242(w_045_1242, w_027_287, w_024_165);
  not1 I045_1264(w_045_1264, w_002_350);
  not1 I045_1313(w_045_1313, w_029_178);
  not1 I045_1328(w_045_1328, w_044_963);
  and2 I045_1333(w_045_1333, w_029_072, w_003_241);
  not1 I045_1349(w_045_1349, w_040_527);
  not1 I045_1414(w_045_1414, w_031_1006);
  nand2 I045_1467(w_045_1467, w_044_074, w_021_020);
  and2 I045_1486(w_045_1486, w_028_010, w_032_190);
  or2  I045_1488(w_045_1488, w_025_1053, w_040_770);
  and2 I045_1489(w_045_1489, w_014_780, w_041_197);
  nand2 I045_1507(w_045_1507, w_034_368, w_010_160);
  and2 I045_1538(w_045_1538, w_041_187, w_008_187);
  or2  I045_1551(w_045_1551, w_022_131, w_002_059);
  not1 I045_1561(w_045_1561, w_000_1792);
  not1 I045_1590(w_045_1590, w_044_1695);
  not1 I045_1596(w_045_1596, w_035_1685);
  not1 I045_1599(w_045_1599, w_015_229);
  not1 I045_1622(w_045_1622, w_041_194);
  nand2 I045_1646(w_045_1646, w_043_037, w_036_650);
  and2 I045_1650(w_045_1650, w_017_179, w_005_1090);
  and2 I045_1653(w_045_1653, w_009_027, w_029_296);
  and2 I045_1659(w_045_1659, w_028_610, w_008_210);
  nand2 I045_1677(w_045_1677, w_020_174, w_019_071);
  or2  I045_1693(w_045_1693, w_019_001, w_026_1221);
  and2 I045_1704(w_045_1704, w_038_413, w_020_387);
  or2  I045_1715(w_045_1715, w_040_472, w_020_539);
  and2 I045_1718(w_045_1718, w_021_151, w_040_024);
  and2 I045_1738(w_045_1738, w_043_004, w_040_080);
  nand2 I045_1756(w_045_1756, w_025_396, w_008_207);
  and2 I045_1806(w_045_1806, w_012_505, w_041_113);
  not1 I045_1824(w_045_1824, w_015_088);
  and2 I045_1830(w_045_1830, w_016_001, w_040_482);
  not1 I045_1833(w_045_1833, w_001_141);
  not1 I045_1878(w_045_1878, w_009_010);
  not1 I046_005(w_046_005, w_032_099);
  or2  I046_008(w_046_008, w_027_326, w_002_054);
  nand2 I046_011(w_046_011, w_019_201, w_025_1399);
  and2 I046_012(w_046_012, w_021_011, w_005_479);
  or2  I046_014(w_046_014, w_033_595, w_006_026);
  and2 I046_017(w_046_017, w_030_000, w_008_488);
  and2 I046_018(w_046_018, w_027_459, w_011_414);
  not1 I046_020(w_046_020, w_018_257);
  nand2 I046_028(w_046_028, w_036_283, w_019_920);
  not1 I046_029(w_046_029, w_034_178);
  not1 I046_030(w_046_030, w_007_036);
  and2 I046_034(w_046_034, w_006_050, w_042_031);
  and2 I046_040(w_046_040, w_007_168, w_041_091);
  and2 I046_042(w_046_042, w_003_056, w_019_213);
  or2  I046_045(w_046_045, w_036_353, w_023_147);
  or2  I046_048(w_046_048, w_044_056, w_040_914);
  nand2 I046_049(w_046_049, w_007_1127, w_022_144);
  nand2 I046_052(w_046_052, w_009_063, w_040_1102);
  not1 I046_054(w_046_054, w_029_504);
  nand2 I046_056(w_046_056, w_015_141, w_033_1417);
  not1 I046_060(w_046_060, w_010_291);
  and2 I046_062(w_046_062, w_042_014, w_019_665);
  not1 I046_066(w_046_066, w_017_1109);
  nand2 I046_070(w_046_070, w_011_208, w_033_629);
  not1 I046_072(w_046_072, w_033_022);
  or2  I046_074(w_046_074, w_029_1328, w_026_195);
  and2 I046_075(w_046_075, w_003_188, w_002_171);
  not1 I046_076(w_046_076, w_005_1393);
  nand2 I046_077(w_046_077, w_014_532, w_035_861);
  not1 I046_078(w_046_078, w_002_240);
  nand2 I046_079(w_046_079, w_037_1238, w_039_1297);
  not1 I046_082(w_046_082, w_039_1906);
  and2 I046_083(w_046_083, w_004_425, w_022_053);
  not1 I046_087(w_046_087, w_010_056);
  or2  I046_090(w_046_090, w_011_204, w_005_101);
  and2 I046_098(w_046_098, w_020_1255, w_010_246);
  nand2 I046_099(w_046_099, w_004_1254, w_042_016);
  not1 I046_105(w_046_105, w_023_553);
  nand2 I046_109(w_046_109, w_012_451, w_004_959);
  or2  I046_114(w_046_114, w_040_1005, w_007_463);
  not1 I046_118(w_046_118, w_002_023);
  nand2 I046_119(w_046_119, w_036_1107, w_014_312);
  nand2 I046_120(w_046_120, w_020_583, w_031_1021);
  and2 I046_121(w_046_121, w_019_027, w_001_1460);
  nand2 I046_122(w_046_122, w_044_675, w_010_278);
  or2  I046_123(w_046_123, w_035_987, w_029_1002);
  or2  I046_124(w_046_124, w_010_095, w_001_107);
  not1 I046_127(w_046_127, w_024_460);
  not1 I046_128(w_046_128, w_043_097);
  and2 I046_130(w_046_130, w_030_354, w_007_171);
  or2  I046_131(w_046_131, w_041_122, w_019_958);
  not1 I046_133(w_046_133, w_008_821);
  not1 I046_134(w_046_134, w_023_333);
  and2 I046_136(w_046_136, w_008_413, w_042_047);
  and2 I046_138(w_046_138, w_043_066, w_005_180);
  nand2 I046_139(w_046_139, w_026_090, w_008_266);
  and2 I046_140(w_046_140, w_025_704, w_026_234);
  or2  I046_145(w_046_145, w_023_625, w_041_131);
  nand2 I046_147(w_046_147, w_003_028, w_020_1143);
  and2 I046_148(w_046_148, w_011_406, w_041_212);
  not1 I046_149(w_046_149, w_001_185);
  or2  I046_156(w_046_156, w_027_006, w_023_708);
  nand2 I046_159(w_046_159, w_032_028, w_034_114);
  and2 I046_168(w_046_168, w_000_163, w_045_251);
  and2 I046_170(w_046_170, w_031_1110, w_016_020);
  not1 I046_171(w_046_171, w_000_1190);
  nand2 I046_173(w_046_173, w_035_600, w_032_023);
  not1 I046_174(w_046_174, w_021_193);
  and2 I046_178(w_046_178, w_039_466, w_017_1534);
  not1 I046_180(w_046_180, w_035_168);
  nand2 I046_181(w_046_181, w_016_029, w_032_030);
  not1 I046_191(w_046_191, w_026_341);
  and2 I046_192(w_046_192, w_044_764, w_017_1453);
  nand2 I046_193(w_046_193, w_033_393, w_018_235);
  nand2 I046_195(w_046_195, w_036_1399, w_019_317);
  and2 I046_198(w_046_198, w_031_786, w_016_012);
  nand2 I046_202(w_046_202, w_037_222, w_022_188);
  nand2 I046_203(w_046_203, w_025_016, w_022_010);
  nand2 I046_207(w_046_207, w_000_494, w_002_086);
  nand2 I046_208(w_046_208, w_000_821, w_032_075);
  nand2 I046_213(w_046_213, w_028_159, w_019_619);
  nand2 I046_215(w_046_215, w_021_111, w_014_255);
  or2  I046_216(w_046_216, w_005_1265, w_032_002);
  and2 I046_218(w_046_218, w_040_447, w_020_135);
  and2 I046_219(w_046_219, w_044_1465, w_032_054);
  and2 I046_220(w_046_220, w_008_748, w_011_109);
  not1 I046_223(w_046_223, w_039_782);
  nand2 I046_225(w_046_225, w_027_207, w_003_259);
  and2 I046_226(w_046_226, w_029_1155, w_045_662);
  or2  I046_228(w_046_228, w_029_565, w_036_238);
  and2 I046_230(w_046_230, w_035_1585, w_028_126);
  or2  I046_231(w_046_231, w_035_1664, w_002_006);
  nand2 I046_232(w_046_232, w_045_617, w_025_300);
  and2 I046_233(w_046_233, w_018_113, w_015_151);
  or2  I046_236(w_046_236, w_037_706, w_008_143);
  nand2 I046_237(w_046_237, w_015_220, w_009_019);
  not1 I046_238(w_046_238, w_028_705);
  not1 I046_247(w_046_247, w_037_1676);
  not1 I046_248(w_046_248, w_003_138);
  or2  I046_250(w_046_250, w_022_416, w_019_407);
  and2 I046_251(w_046_251, w_025_177, w_029_095);
  and2 I046_252(w_046_252, w_029_935, w_040_134);
  nand2 I046_254(w_046_254, w_010_216, w_023_161);
  or2  I046_255(w_046_255, w_019_530, w_014_798);
  or2  I046_258(w_046_258, w_018_088, w_022_069);
  and2 I046_259(w_046_259, w_014_333, w_003_238);
  or2  I046_266(w_046_266, w_005_339, w_040_1286);
  not1 I046_267(w_046_267, w_042_044);
  nand2 I046_270(w_046_270, w_034_269, w_013_258);
  or2  I046_274(w_046_274, w_000_1844, w_027_444);
  and2 I046_276(w_046_276, w_043_063, w_019_614);
  not1 I046_277(w_046_277, w_001_267);
  or2  I046_278(w_046_278, w_017_1686, w_007_627);
  or2  I046_279(w_046_279, w_015_243, w_042_073);
  and2 I046_280(w_046_280, w_026_1135, w_025_137);
  or2  I046_282(w_046_282, w_019_127, w_005_862);
  not1 I047_000(w_047_000, w_034_398);
  or2  I047_007(w_047_007, w_011_611, w_036_450);
  not1 I047_013(w_047_013, w_011_230);
  not1 I047_015(w_047_015, w_030_317);
  or2  I047_019(w_047_019, w_025_913, w_012_652);
  and2 I047_022(w_047_022, w_044_201, w_034_585);
  or2  I047_028(w_047_028, w_005_1638, w_020_1129);
  nand2 I047_031(w_047_031, w_006_177, w_036_482);
  nand2 I047_046(w_047_046, w_035_1601, w_004_1399);
  nand2 I047_054(w_047_054, w_003_262, w_039_1126);
  and2 I047_056(w_047_056, w_044_1093, w_004_042);
  nand2 I047_057(w_047_057, w_003_214, w_009_028);
  and2 I047_059(w_047_059, w_008_289, w_007_828);
  and2 I047_060(w_047_060, w_025_1678, w_032_090);
  or2  I047_062(w_047_062, w_036_492, w_033_218);
  and2 I047_065(w_047_065, w_039_1907, w_030_146);
  and2 I047_073(w_047_073, w_034_109, w_006_176);
  nand2 I047_074(w_047_074, w_007_1467, w_017_1504);
  and2 I047_100(w_047_100, w_012_614, w_018_087);
  not1 I047_103(w_047_103, w_003_028);
  nand2 I047_107(w_047_107, w_026_1418, w_035_760);
  nand2 I047_115(w_047_115, w_000_1132, w_005_1360);
  and2 I047_119(w_047_119, w_044_542, w_030_208);
  nand2 I047_129(w_047_129, w_016_032, w_039_558);
  and2 I047_139(w_047_139, w_031_456, w_016_004);
  or2  I047_140(w_047_140, w_008_747, w_008_620);
  and2 I047_141(w_047_141, w_046_042, w_037_1186);
  nand2 I047_149(w_047_149, w_042_017, w_039_252);
  or2  I047_174(w_047_174, w_010_042, w_032_147);
  and2 I047_175(w_047_175, w_031_468, w_018_204);
  nand2 I047_190(w_047_190, w_017_368, w_022_184);
  or2  I047_194(w_047_194, w_046_156, w_021_241);
  nand2 I047_195(w_047_195, w_014_123, w_028_426);
  not1 I047_196(w_047_196, w_001_165);
  and2 I047_224(w_047_224, w_011_449, w_032_130);
  or2  I047_226(w_047_226, w_023_205, w_002_334);
  nand2 I047_230(w_047_230, w_005_128, w_025_815);
  nand2 I047_231(w_047_231, w_036_282, w_001_1310);
  and2 I047_233(w_047_233, w_023_294, w_038_479);
  not1 I047_235(w_047_235, w_037_1081);
  or2  I047_241(w_047_241, w_036_1034, w_009_017);
  not1 I047_251(w_047_251, w_015_059);
  and2 I047_253(w_047_253, w_020_015, w_018_078);
  nand2 I047_259(w_047_259, w_035_1281, w_019_190);
  or2  I047_262(w_047_262, w_036_488, w_046_052);
  not1 I047_280(w_047_280, w_015_046);
  not1 I047_283(w_047_283, w_044_951);
  or2  I047_288(w_047_288, w_020_875, w_029_490);
  and2 I047_291(w_047_291, w_037_1254, w_021_256);
  nand2 I047_301(w_047_301, w_016_035, w_017_513);
  nand2 I047_303(w_047_303, w_037_906, w_026_879);
  nand2 I047_319(w_047_319, w_025_1611, w_006_276);
  and2 I047_320(w_047_320, w_027_130, w_005_1185);
  and2 I047_329(w_047_329, w_045_365, w_021_182);
  nand2 I047_331(w_047_331, w_032_080, w_013_119);
  or2  I047_332(w_047_332, w_009_015, w_001_1308);
  nand2 I047_335(w_047_335, w_003_233, w_005_1028);
  or2  I047_338(w_047_338, w_037_1344, w_028_777);
  not1 I047_340(w_047_340, w_029_256);
  nand2 I047_341(w_047_341, w_040_312, w_008_051);
  nand2 I047_345(w_047_345, w_018_234, w_034_351);
  and2 I047_362(w_047_362, w_013_203, w_001_1563);
  nand2 I047_363(w_047_363, w_040_273, w_021_111);
  or2  I047_372(w_047_372, w_002_025, w_029_507);
  and2 I047_375(w_047_375, w_028_513, w_023_1179);
  not1 I047_384(w_047_384, w_018_107);
  nand2 I047_386(w_047_386, w_010_023, w_001_028);
  and2 I047_387(w_047_387, w_025_1674, w_021_027);
  and2 I047_391(w_047_391, w_023_902, w_026_1244);
  and2 I047_400(w_047_400, w_020_860, w_008_769);
  or2  I047_404(w_047_404, w_008_268, w_005_137);
  and2 I047_415(w_047_415, w_034_289, w_020_360);
  or2  I047_418(w_047_418, w_002_290, w_016_037);
  and2 I047_419(w_047_419, w_036_200, w_044_1108);
  nand2 I047_425(w_047_425, w_029_899, w_025_355);
  not1 I047_428(w_047_428, w_035_460);
  or2  I047_434(w_047_434, w_004_486, w_012_260);
  or2  I047_441(w_047_441, w_028_552, w_005_608);
  and2 I047_442(w_047_442, w_025_718, w_039_470);
  or2  I047_462(w_047_462, w_043_081, w_023_266);
  or2  I047_465(w_047_465, w_039_568, w_025_1626);
  nand2 I047_475(w_047_475, w_023_349, w_019_692);
  not1 I047_480(w_047_480, w_037_1646);
  or2  I047_489(w_047_489, w_000_1975, w_024_054);
  or2  I047_491(w_047_491, w_041_257, w_013_085);
  and2 I047_496(w_047_496, w_011_865, w_029_042);
  and2 I047_500(w_047_500, w_024_200, w_040_1237);
  not1 I047_501(w_047_501, w_006_197);
  or2  I047_503(w_047_503, w_034_430, w_015_161);
  nand2 I047_518(w_047_518, w_038_317, w_023_820);
  and2 I047_524(w_047_524, w_041_026, w_043_100);
  and2 I047_532(w_047_532, w_016_001, w_018_008);
  and2 I047_537(w_047_537, w_003_041, w_011_118);
  not1 I047_543(w_047_543, w_011_533);
  not1 I047_545(w_047_545, w_019_105);
  or2  I047_548(w_047_548, w_040_015, w_024_189);
  not1 I047_550(w_047_550, w_046_128);
  or2  I047_552(w_047_552, w_027_130, w_004_112);
  not1 I047_558(w_047_558, w_000_491);
  or2  I047_562(w_047_562, w_013_248, w_045_1561);
  not1 I047_568(w_047_568, w_045_226);
  not1 I047_569(w_047_569, w_009_060);
  nand2 I047_570(w_047_570, w_032_087, w_004_1524);
  and2 I047_573(w_047_573, w_014_337, w_003_244);
  not1 I047_577(w_047_577, w_025_1540);
  nand2 I047_579(w_047_579, w_011_112, w_003_066);
  not1 I047_585(w_047_585, w_009_084);
  and2 I047_594(w_047_594, w_030_592, w_018_068);
  nand2 I047_595(w_047_595, w_017_736, w_005_778);
  not1 I047_599(w_047_599, w_020_606);
  nand2 I047_606(w_047_606, w_037_081, w_046_208);
  nand2 I047_632(w_047_632, w_003_220, w_025_036);
  not1 I047_639(w_047_639, w_029_414);
  nand2 I047_640(w_047_640, w_007_084, w_032_091);
  not1 I047_641(w_047_641, w_019_430);
  not1 I047_653(w_047_653, w_008_073);
  nand2 I047_675(w_047_675, w_000_1274, w_031_981);
  nand2 I047_692(w_047_692, w_006_030, w_038_405);
  and2 I047_698(w_047_698, w_033_099, w_017_1900);
  or2  I048_000(w_048_000, w_005_281, w_031_495);
  or2  I048_007(w_048_007, w_036_408, w_039_1634);
  not1 I048_010(w_048_010, w_027_063);
  and2 I048_018(w_048_018, w_010_169, w_033_1429);
  not1 I048_021(w_048_021, w_006_272);
  and2 I048_033(w_048_033, w_046_202, w_033_722);
  nand2 I048_053(w_048_053, w_019_772, w_033_1438);
  and2 I048_054(w_048_054, w_002_531, w_020_687);
  nand2 I048_057(w_048_057, w_040_959, w_016_021);
  or2  I048_072(w_048_072, w_036_1493, w_021_010);
  nand2 I048_073(w_048_073, w_037_1234, w_018_187);
  not1 I048_077(w_048_077, w_008_096);
  and2 I048_090(w_048_090, w_029_553, w_020_220);
  or2  I048_092(w_048_092, w_000_827, w_036_1273);
  not1 I048_098(w_048_098, w_023_1283);
  or2  I048_117(w_048_117, w_000_1557, w_025_1321);
  or2  I048_132(w_048_132, w_003_062, w_001_232);
  nand2 I048_134(w_048_134, w_044_1481, w_047_139);
  not1 I048_135(w_048_135, w_018_013);
  not1 I048_142(w_048_142, w_001_1491);
  or2  I048_148(w_048_148, w_037_1211, w_035_358);
  not1 I048_159(w_048_159, w_030_181);
  and2 I048_162(w_048_162, w_005_905, w_042_022);
  or2  I048_171(w_048_171, w_019_091, w_013_267);
  and2 I048_194(w_048_194, w_016_031, w_013_040);
  and2 I048_202(w_048_202, w_015_127, w_008_163);
  and2 I048_204(w_048_204, w_047_491, w_017_1103);
  or2  I048_209(w_048_209, w_044_1077, w_005_1464);
  or2  I048_213(w_048_213, w_043_001, w_014_121);
  or2  I048_229(w_048_229, w_021_199, w_030_161);
  nand2 I048_230(w_048_230, w_047_363, w_034_345);
  not1 I048_236(w_048_236, w_009_088);
  or2  I048_243(w_048_243, w_047_335, w_010_194);
  nand2 I048_250(w_048_250, w_045_1489, w_002_418);
  not1 I048_253(w_048_253, w_030_003);
  nand2 I048_276(w_048_276, w_003_253, w_040_306);
  nand2 I048_312(w_048_312, w_030_007, w_032_126);
  nand2 I048_317(w_048_317, w_028_871, w_037_1140);
  or2  I048_326(w_048_326, w_021_221, w_042_001);
  or2  I048_328(w_048_328, w_023_012, w_007_1443);
  or2  I048_345(w_048_345, w_045_547, w_034_583);
  nand2 I048_348(w_048_348, w_011_401, w_030_261);
  not1 I048_354(w_048_354, w_018_168);
  and2 I048_358(w_048_358, w_043_023, w_032_197);
  and2 I048_373(w_048_373, w_040_568, w_006_322);
  and2 I048_383(w_048_383, w_037_953, w_023_1265);
  not1 I048_405(w_048_405, w_028_292);
  and2 I048_406(w_048_406, w_038_459, w_014_229);
  or2  I048_409(w_048_409, w_027_427, w_029_644);
  nand2 I048_415(w_048_415, w_024_197, w_024_243);
  and2 I048_416(w_048_416, w_021_053, w_003_248);
  nand2 I048_421(w_048_421, w_039_1273, w_025_015);
  or2  I048_431(w_048_431, w_006_011, w_047_332);
  and2 I048_432(w_048_432, w_022_122, w_002_022);
  or2  I048_436(w_048_436, w_007_017, w_022_135);
  nand2 I048_439(w_048_439, w_021_033, w_021_249);
  or2  I048_440(w_048_440, w_009_071, w_036_047);
  nand2 I048_446(w_048_446, w_017_471, w_037_1674);
  nand2 I048_447(w_048_447, w_041_231, w_007_1292);
  and2 I048_472(w_048_472, w_026_001, w_021_044);
  or2  I048_473(w_048_473, w_024_345, w_047_375);
  or2  I048_479(w_048_479, w_045_1181, w_007_1110);
  not1 I048_487(w_048_487, w_026_1316);
  or2  I048_520(w_048_520, w_022_146, w_044_166);
  not1 I048_527(w_048_527, w_044_1723);
  or2  I048_536(w_048_536, w_022_323, w_000_449);
  not1 I048_546(w_048_546, w_038_395);
  nand2 I048_548(w_048_548, w_045_731, w_017_033);
  or2  I048_551(w_048_551, w_037_072, w_037_137);
  nand2 I048_553(w_048_553, w_030_069, w_045_1596);
  or2  I048_554(w_048_554, w_005_126, w_000_038);
  and2 I048_560(w_048_560, w_000_970, w_029_085);
  and2 I048_561(w_048_561, w_045_475, w_047_331);
  or2  I048_564(w_048_564, w_003_067, w_031_1019);
  not1 I048_567(w_048_567, w_040_127);
  and2 I048_583(w_048_583, w_035_1450, w_027_461);
  or2  I048_584(w_048_584, w_017_1416, w_036_692);
  nand2 I048_588(w_048_588, w_032_059, w_013_127);
  or2  I048_593(w_048_593, w_025_668, w_029_1127);
  and2 I048_597(w_048_597, w_000_1341, w_009_017);
  not1 I048_598(w_048_598, w_016_020);
  not1 I048_622(w_048_622, w_002_060);
  nand2 I048_623(w_048_623, w_022_136, w_021_169);
  and2 I048_627(w_048_627, w_026_069, w_046_139);
  nand2 I048_629(w_048_629, w_032_084, w_030_411);
  not1 I048_637(w_048_637, w_015_234);
  nand2 I048_649(w_048_649, w_034_205, w_026_661);
  and2 I048_651(w_048_651, w_025_747, w_035_657);
  not1 I048_652(w_048_652, w_012_056);
  not1 I048_668(w_048_668, w_007_838);
  nand2 I048_671(w_048_671, w_008_362, w_021_081);
  and2 I048_672(w_048_672, w_035_647, w_043_004);
  or2  I048_676(w_048_676, w_031_874, w_024_1221);
  or2  I048_677(w_048_677, w_011_721, w_029_017);
  not1 I048_694(w_048_694, w_011_830);
  and2 I048_705(w_048_705, w_010_293, w_029_554);
  or2  I048_713(w_048_713, w_006_099, w_035_1397);
  and2 I048_724(w_048_724, w_015_125, w_024_1570);
  or2  I048_742(w_048_742, w_011_610, w_011_190);
  and2 I048_746(w_048_746, w_014_467, w_012_241);
  nand2 I048_751(w_048_751, w_032_015, w_000_577);
  nand2 I048_752(w_048_752, w_047_573, w_047_386);
  or2  I048_758(w_048_758, w_004_677, w_017_867);
  and2 I048_762(w_048_762, w_036_045, w_008_288);
  and2 I048_770(w_048_770, w_034_308, w_032_156);
  not1 I048_777(w_048_777, w_007_744);
  not1 I048_781(w_048_781, w_007_1481);
  not1 I048_783(w_048_783, w_001_120);
  or2  I048_787(w_048_787, w_038_076, w_046_191);
  or2  I048_792(w_048_792, w_019_608, w_007_309);
  and2 I048_797(w_048_797, w_033_113, w_016_021);
  not1 I048_799(w_048_799, w_012_524);
  and2 I048_802(w_048_802, w_004_1835, w_032_092);
  and2 I048_824(w_048_824, w_033_713, w_006_048);
  not1 I048_827(w_048_827, w_037_1451);
  or2  I048_849(w_048_849, w_046_173, w_001_662);
  nand2 I048_850(w_048_850, w_002_545, w_007_107);
  nand2 I048_881(w_048_881, w_025_1426, w_020_395);
  and2 I048_884(w_048_884, w_028_152, w_021_083);
  nand2 I048_897(w_048_897, w_001_196, w_003_139);
  and2 I048_901(w_048_901, w_040_061, w_016_010);
  not1 I048_904(w_048_904, w_046_122);
  nand2 I048_908(w_048_908, w_001_1425, w_044_1566);
  not1 I048_909(w_048_909, w_016_030);
  and2 I048_918(w_048_918, w_030_715, w_002_275);
  not1 I048_963(w_048_963, w_009_088);
  not1 I048_966(w_048_966, w_043_075);
  or2  I048_974(w_048_974, w_000_1951, w_021_221);
  nand2 I049_008(w_049_008, w_018_214, w_015_211);
  or2  I049_013(w_049_013, w_015_159, w_000_654);
  or2  I049_020(w_049_020, w_048_564, w_014_150);
  or2  I049_031(w_049_031, w_005_1324, w_030_262);
  and2 I049_043(w_049_043, w_007_1543, w_023_359);
  or2  I049_047(w_049_047, w_046_178, w_038_153);
  not1 I049_055(w_049_055, w_026_650);
  and2 I049_076(w_049_076, w_026_1223, w_048_010);
  not1 I049_077(w_049_077, w_039_881);
  or2  I049_080(w_049_080, w_036_992, w_013_328);
  nand2 I049_087(w_049_087, w_018_280, w_004_345);
  nand2 I049_095(w_049_095, w_017_1393, w_040_512);
  and2 I049_099(w_049_099, w_014_643, w_029_119);
  not1 I049_110(w_049_110, w_029_739);
  or2  I049_112(w_049_112, w_048_439, w_004_725);
  not1 I049_132(w_049_132, w_047_585);
  not1 I049_157(w_049_157, w_040_1076);
  nand2 I049_169(w_049_169, w_046_180, w_029_731);
  or2  I049_190(w_049_190, w_008_280, w_048_622);
  nand2 I049_206(w_049_206, w_044_033, w_001_017);
  nand2 I049_213(w_049_213, w_000_471, w_007_109);
  nand2 I049_220(w_049_220, w_041_115, w_040_1013);
  nand2 I049_241(w_049_241, w_014_814, w_048_348);
  or2  I049_252(w_049_252, w_008_262, w_034_441);
  not1 I049_253(w_049_253, w_007_1617);
  or2  I049_255(w_049_255, w_028_664, w_045_1203);
  or2  I049_260(w_049_260, w_020_545, w_021_035);
  or2  I049_272(w_049_272, w_036_375, w_038_364);
  or2  I049_275(w_049_275, w_014_643, w_048_421);
  not1 I049_277(w_049_277, w_025_1469);
  not1 I049_282(w_049_282, w_031_050);
  nand2 I049_289(w_049_289, w_034_122, w_039_100);
  not1 I049_300(w_049_300, w_009_101);
  or2  I049_306(w_049_306, w_004_093, w_017_524);
  nand2 I049_309(w_049_309, w_005_1223, w_046_109);
  or2  I049_311(w_049_311, w_006_135, w_038_236);
  not1 I049_315(w_049_315, w_028_038);
  nand2 I049_327(w_049_327, w_021_118, w_043_028);
  nand2 I049_335(w_049_335, w_041_279, w_046_078);
  nand2 I049_336(w_049_336, w_016_000, w_006_298);
  not1 I049_345(w_049_345, w_002_138);
  and2 I049_347(w_049_347, w_000_491, w_015_113);
  not1 I049_370(w_049_370, w_014_130);
  and2 I049_377(w_049_377, w_012_122, w_044_682);
  not1 I049_378(w_049_378, w_032_233);
  nand2 I049_393(w_049_393, w_027_146, w_020_1115);
  or2  I049_403(w_049_403, w_016_011, w_044_443);
  nand2 I049_404(w_049_404, w_025_080, w_022_015);
  not1 I049_429(w_049_429, w_011_021);
  not1 I049_433(w_049_433, w_033_876);
  or2  I049_447(w_049_447, w_045_786, w_012_632);
  nand2 I049_454(w_049_454, w_004_1815, w_048_431);
  or2  I049_457(w_049_457, w_046_147, w_033_232);
  nand2 I049_488(w_049_488, w_039_516, w_010_132);
  or2  I049_489(w_049_489, w_046_237, w_041_126);
  or2  I049_494(w_049_494, w_008_692, w_024_247);
  or2  I049_515(w_049_515, w_016_006, w_036_1104);
  or2  I049_519(w_049_519, w_012_507, w_047_428);
  or2  I049_521(w_049_521, w_023_026, w_015_163);
  and2 I049_529(w_049_529, w_042_002, w_041_081);
  and2 I049_530(w_049_530, w_008_252, w_031_012);
  not1 I049_537(w_049_537, w_025_1668);
  not1 I049_541(w_049_541, w_031_287);
  or2  I049_542(w_049_542, w_016_024, w_028_586);
  or2  I049_543(w_049_543, w_014_251, w_003_011);
  nand2 I049_548(w_049_548, w_032_112, w_035_1707);
  nand2 I049_554(w_049_554, w_010_071, w_043_025);
  and2 I049_571(w_049_571, w_024_349, w_026_156);
  and2 I049_584(w_049_584, w_025_639, w_009_047);
  and2 I049_594(w_049_594, w_018_260, w_017_744);
  nand2 I049_595(w_049_595, w_047_362, w_025_521);
  and2 I049_601(w_049_601, w_045_580, w_015_291);
  or2  I049_606(w_049_606, w_040_294, w_020_134);
  nand2 I049_616(w_049_616, w_042_102, w_010_268);
  nand2 I049_620(w_049_620, w_015_212, w_018_155);
  or2  I049_634(w_049_634, w_030_392, w_040_823);
  or2  I049_651(w_049_651, w_005_479, w_006_014);
  not1 I049_700(w_049_700, w_036_258);
  or2  I049_710(w_049_710, w_006_228, w_019_202);
  and2 I049_738(w_049_738, w_033_168, w_034_204);
  or2  I049_786(w_049_786, w_020_423, w_038_368);
  not1 I049_803(w_049_803, w_009_007);
  and2 I049_813(w_049_813, w_045_874, w_012_242);
  nand2 I049_869(w_049_869, w_011_117, w_017_1220);
  or2  I049_871(w_049_871, w_021_271, w_033_109);
  or2  I049_882(w_049_882, w_008_734, w_013_104);
  or2  I049_909(w_049_909, w_018_251, w_006_201);
  and2 I049_929(w_049_929, w_029_263, w_042_064);
  nand2 I049_962(w_049_962, w_041_149, w_042_062);
  nand2 I049_971(w_049_971, w_006_285, w_039_1280);
  and2 I049_999(w_049_999, w_017_863, w_044_1417);
  not1 I049_1001(w_049_1001, w_016_034);
  or2  I049_1006(w_049_1006, w_007_381, w_003_311);
  nand2 I049_1033(w_049_1033, w_016_022, w_025_1425);
  nand2 I049_1041(w_049_1041, w_018_038, w_013_116);
  nand2 I049_1057(w_049_1057, w_017_896, w_047_319);
  nand2 I049_1058(w_049_1058, w_042_009, w_010_109);
  not1 I049_1067(w_049_1067, w_041_245);
  or2  I049_1075(w_049_1075, w_024_1297, w_008_110);
  and2 I049_1111(w_049_1111, w_014_729, w_004_101);
  and2 I049_1129(w_049_1129, w_040_323, w_002_227);
  or2  I049_1136(w_049_1136, w_045_1806, w_032_235);
  and2 I049_1140(w_049_1140, w_017_1464, w_030_334);
  nand2 I049_1143(w_049_1143, w_008_289, w_012_310);
  or2  I049_1157(w_049_1157, w_000_1663, w_012_653);
  and2 I049_1165(w_049_1165, w_037_942, w_025_573);
  not1 I049_1167(w_049_1167, w_025_782);
  and2 I049_1169(w_049_1169, w_016_006, w_028_079);
  not1 I049_1207(w_049_1207, w_008_549);
  nand2 I049_1221(w_049_1221, w_043_079, w_041_282);
  not1 I049_1227(w_049_1227, w_024_435);
  or2  I049_1243(w_049_1243, w_003_205, w_038_118);
  or2  I049_1303(w_049_1303, w_032_092, w_046_225);
  not1 I049_1320(w_049_1320, w_028_195);
  nand2 I049_1359(w_049_1359, w_009_018, w_026_152);
  and2 I050_010(w_050_010, w_037_1084, w_014_121);
  or2  I050_015(w_050_015, w_034_276, w_006_064);
  and2 I050_016(w_050_016, w_000_1883, w_016_036);
  not1 I050_020(w_050_020, w_027_465);
  nand2 I050_032(w_050_032, w_033_895, w_017_525);
  not1 I050_033(w_050_033, w_038_395);
  not1 I050_038(w_050_038, w_016_014);
  not1 I050_041(w_050_041, w_006_226);
  or2  I050_044(w_050_044, w_003_289, w_017_325);
  and2 I050_045(w_050_045, w_032_134, w_023_257);
  and2 I050_052(w_050_052, w_007_081, w_017_914);
  and2 I050_066(w_050_066, w_001_043, w_011_062);
  and2 I050_069(w_050_069, w_037_999, w_007_109);
  or2  I050_071(w_050_071, w_009_059, w_033_1650);
  not1 I050_079(w_050_079, w_007_205);
  and2 I050_090(w_050_090, w_013_255, w_026_106);
  nand2 I050_097(w_050_097, w_001_447, w_037_155);
  not1 I050_101(w_050_101, w_011_424);
  and2 I050_102(w_050_102, w_021_007, w_046_029);
  or2  I050_105(w_050_105, w_009_025, w_005_090);
  not1 I050_154(w_050_154, w_035_991);
  not1 I050_155(w_050_155, w_031_1126);
  and2 I050_161(w_050_161, w_047_692, w_026_055);
  not1 I050_162(w_050_162, w_009_076);
  nand2 I050_169(w_050_169, w_012_667, w_012_254);
  not1 I050_174(w_050_174, w_016_033);
  and2 I050_175(w_050_175, w_049_213, w_011_461);
  and2 I050_176(w_050_176, w_024_1383, w_022_009);
  or2  I050_181(w_050_181, w_034_196, w_032_000);
  not1 I050_185(w_050_185, w_037_876);
  nand2 I050_190(w_050_190, w_018_084, w_017_398);
  or2  I050_191(w_050_191, w_006_239, w_021_119);
  nand2 I050_193(w_050_193, w_025_788, w_025_1456);
  or2  I050_197(w_050_197, w_039_133, w_036_1397);
  not1 I050_217(w_050_217, w_000_470);
  nand2 I050_220(w_050_220, w_044_1690, w_007_1420);
  or2  I050_225(w_050_225, w_015_187, w_030_422);
  and2 I050_257(w_050_257, w_035_805, w_033_1077);
  not1 I050_266(w_050_266, w_036_1366);
  or2  I050_275(w_050_275, w_023_449, w_025_837);
  nand2 I050_276(w_050_276, w_018_122, w_021_216);
  nand2 I050_314(w_050_314, w_046_255, w_029_119);
  not1 I050_321(w_050_321, w_019_289);
  or2  I050_322(w_050_322, w_042_000, w_017_333);
  or2  I050_326(w_050_326, w_046_005, w_012_021);
  nand2 I050_342(w_050_342, w_040_1276, w_034_690);
  or2  I050_352(w_050_352, w_017_1439, w_020_1144);
  nand2 I050_353(w_050_353, w_002_103, w_049_700);
  or2  I050_354(w_050_354, w_022_074, w_017_1392);
  not1 I050_362(w_050_362, w_033_672);
  and2 I050_367(w_050_367, w_048_358, w_044_1134);
  nand2 I050_368(w_050_368, w_012_334, w_035_188);
  or2  I050_370(w_050_370, w_039_306, w_003_258);
  not1 I050_380(w_050_380, w_007_561);
  not1 I050_382(w_050_382, w_029_036);
  or2  I050_383(w_050_383, w_048_676, w_014_109);
  and2 I050_393(w_050_393, w_007_534, w_033_195);
  and2 I050_395(w_050_395, w_046_252, w_041_191);
  nand2 I050_406(w_050_406, w_026_723, w_003_188);
  not1 I050_418(w_050_418, w_029_856);
  not1 I050_420(w_050_420, w_012_596);
  and2 I050_435(w_050_435, w_032_233, w_042_074);
  nand2 I050_438(w_050_438, w_006_245, w_002_426);
  and2 I050_448(w_050_448, w_049_1227, w_012_441);
  nand2 I050_462(w_050_462, w_003_158, w_035_036);
  or2  I050_468(w_050_468, w_029_365, w_008_799);
  not1 I050_499(w_050_499, w_030_447);
  nand2 I050_502(w_050_502, w_011_679, w_008_132);
  or2  I050_552(w_050_552, w_011_068, w_047_632);
  or2  I050_556(w_050_556, w_023_1327, w_029_615);
  and2 I050_562(w_050_562, w_030_306, w_009_049);
  nand2 I050_565(w_050_565, w_009_066, w_013_249);
  or2  I050_597(w_050_597, w_008_228, w_035_102);
  or2  I050_610(w_050_610, w_041_022, w_046_259);
  not1 I050_614(w_050_614, w_003_227);
  or2  I050_671(w_050_671, w_015_171, w_012_337);
  not1 I050_683(w_050_683, w_021_079);
  nand2 I050_686(w_050_686, w_040_312, w_033_634);
  nand2 I050_715(w_050_715, w_019_599, w_026_937);
  not1 I050_718(w_050_718, w_043_035);
  nand2 I050_731(w_050_731, w_036_982, w_034_115);
  not1 I050_749(w_050_749, w_049_882);
  not1 I050_751(w_050_751, w_002_266);
  nand2 I050_760(w_050_760, w_012_450, w_025_216);
  or2  I050_764(w_050_764, w_014_296, w_038_304);
  and2 I050_802(w_050_802, w_008_018, w_022_254);
  or2  I050_814(w_050_814, w_016_004, w_015_245);
  nand2 I050_819(w_050_819, w_023_915, w_019_005);
  and2 I050_855(w_050_855, w_031_343, w_017_1077);
  not1 I050_875(w_050_875, w_006_111);
  or2  I050_897(w_050_897, w_041_065, w_013_187);
  or2  I050_961(w_050_961, w_007_061, w_017_622);
  not1 I050_967(w_050_967, w_033_284);
  not1 I050_972(w_050_972, w_035_1391);
  nand2 I050_994(w_050_994, w_027_384, w_046_030);
  and2 I050_1020(w_050_1020, w_023_019, w_005_951);
  not1 I050_1023(w_050_1023, w_020_1038);
  or2  I050_1045(w_050_1045, w_017_018, w_002_182);
  and2 I050_1052(w_050_1052, w_024_790, w_013_313);
  and2 I050_1057(w_050_1057, w_001_325, w_042_017);
  not1 I050_1082(w_050_1082, w_036_319);
  or2  I050_1088(w_050_1088, w_003_098, w_012_042);
  or2  I050_1119(w_050_1119, w_004_1121, w_024_1615);
  not1 I050_1147(w_050_1147, w_008_009);
  or2  I050_1148(w_050_1148, w_016_028, w_011_000);
  nand2 I050_1158(w_050_1158, w_008_580, w_017_1227);
  not1 I050_1164(w_050_1164, w_034_459);
  nand2 I050_1200(w_050_1200, w_041_268, w_029_1074);
  or2  I050_1218(w_050_1218, w_001_1030, w_005_005);
  not1 I050_1224(w_050_1224, w_034_083);
  not1 I050_1231(w_050_1231, w_044_132);
  and2 I050_1239(w_050_1239, w_013_217, w_022_028);
  and2 I050_1244(w_050_1244, w_004_1046, w_034_074);
  not1 I050_1293(w_050_1293, w_034_254);
  and2 I050_1319(w_050_1319, w_042_062, w_026_790);
  and2 I050_1344(w_050_1344, w_049_300, w_006_099);
  nand2 I050_1369(w_050_1369, w_029_720, w_024_761);
  or2  I050_1374(w_050_1374, w_036_337, w_011_031);
  nand2 I050_1379(w_050_1379, w_019_868, w_000_921);
  nand2 I050_1383(w_050_1383, w_048_527, w_024_593);
  and2 I050_1390(w_050_1390, w_035_546, w_006_057);
  nand2 I050_1394(w_050_1394, w_028_102, w_039_595);
  and2 I050_1397(w_050_1397, w_033_1193, w_037_1494);
  and2 I050_1398(w_050_1398, w_016_037, w_012_400);
  not1 I050_1405(w_050_1405, w_020_405);
  not1 I050_1433(w_050_1433, w_028_323);
  not1 I050_1435(w_050_1435, w_013_000);
  not1 I050_1452(w_050_1452, w_020_753);
  or2  I050_1469(w_050_1469, w_030_663, w_009_003);
  not1 I050_1499(w_050_1499, w_000_887);
  and2 I050_1537(w_050_1537, w_022_413, w_001_785);
  nand2 I051_020(w_051_020, w_042_037, w_018_014);
  or2  I051_022(w_051_022, w_039_113, w_027_496);
  or2  I051_023(w_051_023, w_031_051, w_013_102);
  or2  I051_026(w_051_026, w_036_1174, w_030_653);
  nand2 I051_027(w_051_027, w_023_648, w_023_732);
  or2  I051_046(w_051_046, w_049_1136, w_040_390);
  and2 I051_074(w_051_074, w_049_869, w_012_648);
  or2  I051_108(w_051_108, w_039_1726, w_027_183);
  nand2 I051_121(w_051_121, w_017_619, w_003_302);
  or2  I051_126(w_051_126, w_030_105, w_009_106);
  or2  I051_127(w_051_127, w_035_844, w_033_087);
  nand2 I051_143(w_051_143, w_050_1239, w_017_1312);
  and2 I051_149(w_051_149, w_019_290, w_029_502);
  not1 I051_184(w_051_184, w_013_149);
  or2  I051_190(w_051_190, w_050_760, w_008_202);
  nand2 I051_198(w_051_198, w_000_436, w_004_607);
  nand2 I051_202(w_051_202, w_045_524, w_043_089);
  and2 I051_209(w_051_209, w_008_257, w_045_721);
  and2 I051_210(w_051_210, w_049_1167, w_044_1095);
  nand2 I051_230(w_051_230, w_023_1612, w_000_1977);
  and2 I051_246(w_051_246, w_027_344, w_021_153);
  nand2 I051_252(w_051_252, w_038_410, w_038_372);
  not1 I051_265(w_051_265, w_041_004);
  or2  I051_268(w_051_268, w_015_208, w_033_1049);
  nand2 I051_273(w_051_273, w_035_1510, w_023_101);
  or2  I051_274(w_051_274, w_036_123, w_033_1116);
  not1 I051_285(w_051_285, w_000_331);
  and2 I051_290(w_051_290, w_025_1651, w_015_253);
  not1 I051_291(w_051_291, w_015_225);
  nand2 I051_292(w_051_292, w_013_219, w_013_192);
  nand2 I051_294(w_051_294, w_008_079, w_014_614);
  nand2 I051_310(w_051_310, w_007_858, w_021_239);
  not1 I051_347(w_051_347, w_015_020);
  or2  I051_382(w_051_382, w_031_1052, w_047_489);
  and2 I051_407(w_051_407, w_013_252, w_047_434);
  not1 I051_422(w_051_422, w_038_130);
  not1 I051_425(w_051_425, w_012_556);
  nand2 I051_431(w_051_431, w_030_630, w_044_897);
  and2 I051_440(w_051_440, w_033_016, w_007_829);
  nand2 I051_455(w_051_455, w_049_393, w_037_262);
  not1 I051_469(w_051_469, w_011_794);
  not1 I051_480(w_051_480, w_032_154);
  not1 I051_501(w_051_501, w_028_826);
  nand2 I051_559(w_051_559, w_025_1037, w_008_513);
  not1 I051_563(w_051_563, w_050_1405);
  not1 I051_571(w_051_571, w_001_1531);
  and2 I051_576(w_051_576, w_010_159, w_009_023);
  nand2 I051_580(w_051_580, w_024_1563, w_003_297);
  and2 I051_581(w_051_581, w_047_425, w_002_038);
  not1 I051_582(w_051_582, w_042_113);
  not1 I051_595(w_051_595, w_029_377);
  or2  I051_621(w_051_621, w_044_047, w_041_247);
  or2  I051_628(w_051_628, w_013_299, w_008_316);
  and2 I051_633(w_051_633, w_008_067, w_026_843);
  or2  I051_638(w_051_638, w_011_109, w_021_158);
  nand2 I051_640(w_051_640, w_009_094, w_038_438);
  and2 I051_643(w_051_643, w_024_285, w_013_257);
  not1 I051_649(w_051_649, w_042_084);
  and2 I051_653(w_051_653, w_039_142, w_010_357);
  or2  I051_670(w_051_670, w_050_314, w_039_266);
  and2 I051_673(w_051_673, w_032_170, w_000_1924);
  or2  I051_675(w_051_675, w_034_031, w_039_092);
  nand2 I051_701(w_051_701, w_047_241, w_036_1438);
  or2  I051_702(w_051_702, w_040_134, w_030_348);
  or2  I051_703(w_051_703, w_040_1320, w_007_1345);
  and2 I051_710(w_051_710, w_023_204, w_002_432);
  nand2 I051_714(w_051_714, w_026_267, w_026_311);
  or2  I051_735(w_051_735, w_046_087, w_032_208);
  nand2 I051_768(w_051_768, w_014_445, w_027_261);
  or2  I051_773(w_051_773, w_017_1873, w_033_1099);
  not1 I051_777(w_051_777, w_031_057);
  nand2 I051_783(w_051_783, w_001_451, w_004_937);
  and2 I051_804(w_051_804, w_045_1153, w_001_309);
  or2  I051_812(w_051_812, w_005_1408, w_021_034);
  or2  I051_828(w_051_828, w_009_015, w_010_118);
  not1 I051_837(w_051_837, w_011_188);
  and2 I051_847(w_051_847, w_000_1552, w_034_372);
  nand2 I051_849(w_051_849, w_005_508, w_037_541);
  not1 I051_853(w_051_853, w_016_037);
  or2  I051_868(w_051_868, w_010_375, w_044_1383);
  not1 I051_881(w_051_881, w_002_558);
  not1 I051_891(w_051_891, w_033_476);
  not1 I051_939(w_051_939, w_010_066);
  nand2 I051_947(w_051_947, w_006_029, w_018_249);
  nand2 I051_958(w_051_958, w_016_026, w_027_203);
  and2 I051_960(w_051_960, w_018_064, w_001_247);
  or2  I051_982(w_051_982, w_009_001, w_017_005);
  nand2 I051_992(w_051_992, w_019_135, w_038_290);
  not1 I051_996(w_051_996, w_012_186);
  not1 I051_1001(w_051_1001, w_001_344);
  nand2 I051_1012(w_051_1012, w_002_375, w_003_114);
  or2  I051_1015(w_051_1015, w_033_083, w_050_079);
  or2  I051_1022(w_051_1022, w_012_188, w_041_107);
  not1 I051_1023(w_051_1023, w_030_140);
  not1 I051_1044(w_051_1044, w_029_582);
  not1 I051_1064(w_051_1064, w_023_852);
  nand2 I051_1068(w_051_1068, w_039_1227, w_036_1174);
  not1 I051_1073(w_051_1073, w_004_1009);
  not1 I051_1092(w_051_1092, w_022_279);
  or2  I052_011(w_052_011, w_029_220, w_022_408);
  or2  I052_016(w_052_016, w_009_068, w_015_099);
  nand2 I052_017(w_052_017, w_027_220, w_026_1031);
  and2 I052_031(w_052_031, w_047_100, w_033_347);
  or2  I052_034(w_052_034, w_002_442, w_018_267);
  not1 I052_037(w_052_037, w_018_024);
  nand2 I052_042(w_052_042, w_030_345, w_006_316);
  and2 I052_047(w_052_047, w_028_472, w_037_510);
  and2 I052_058(w_052_058, w_017_1383, w_045_662);
  nand2 I052_059(w_052_059, w_002_464, w_031_753);
  nand2 I052_061(w_052_061, w_043_042, w_004_816);
  or2  I052_145(w_052_145, w_024_606, w_043_085);
  not1 I052_166(w_052_166, w_050_855);
  not1 I052_173(w_052_173, w_003_111);
  nand2 I052_185(w_052_185, w_023_1226, w_021_237);
  not1 I052_198(w_052_198, w_034_057);
  nand2 I052_205(w_052_205, w_019_142, w_046_020);
  and2 I052_218(w_052_218, w_005_961, w_034_476);
  and2 I052_242(w_052_242, w_015_044, w_049_1320);
  or2  I052_266(w_052_266, w_009_012, w_037_090);
  or2  I052_309(w_052_309, w_036_149, w_014_537);
  nand2 I052_338(w_052_338, w_011_152, w_043_062);
  or2  I052_382(w_052_382, w_032_005, w_025_1169);
  and2 I052_388(w_052_388, w_014_598, w_034_245);
  not1 I052_391(w_052_391, w_007_931);
  and2 I052_392(w_052_392, w_015_004, w_040_1138);
  or2  I052_405(w_052_405, w_026_1429, w_025_976);
  or2  I052_432(w_052_432, w_034_316, w_000_1696);
  and2 I052_440(w_052_440, w_020_112, w_014_702);
  and2 I052_461(w_052_461, w_020_229, w_029_125);
  or2  I052_465(w_052_465, w_048_436, w_011_107);
  nand2 I052_498(w_052_498, w_047_283, w_048_746);
  or2  I052_503(w_052_503, w_024_998, w_048_204);
  nand2 I052_547(w_052_547, w_022_298, w_030_664);
  and2 I052_566(w_052_566, w_012_044, w_040_869);
  and2 I052_574(w_052_574, w_046_072, w_006_017);
  or2  I052_587(w_052_587, w_016_019, w_009_032);
  and2 I052_640(w_052_640, w_018_233, w_020_312);
  and2 I052_667(w_052_667, w_048_472, w_029_1240);
  or2  I052_711(w_052_711, w_013_163, w_013_077);
  or2  I052_715(w_052_715, w_010_169, w_006_038);
  or2  I052_731(w_052_731, w_046_203, w_038_211);
  not1 I052_733(w_052_733, w_025_389);
  or2  I052_743(w_052_743, w_025_739, w_011_463);
  and2 I052_817(w_052_817, w_048_092, w_048_520);
  not1 I052_825(w_052_825, w_040_037);
  nand2 I052_844(w_052_844, w_014_577, w_048_328);
  not1 I052_853(w_052_853, w_050_1164);
  nand2 I052_857(w_052_857, w_012_657, w_014_644);
  and2 I052_877(w_052_877, w_015_068, w_043_073);
  and2 I052_904(w_052_904, w_040_102, w_014_326);
  nand2 I052_925(w_052_925, w_031_847, w_015_155);
  and2 I052_947(w_052_947, w_049_1359, w_033_1243);
  and2 I052_952(w_052_952, w_001_221, w_050_1224);
  or2  I052_965(w_052_965, w_010_192, w_003_081);
  or2  I052_981(w_052_981, w_044_1427, w_017_644);
  or2  I052_987(w_052_987, w_050_071, w_022_038);
  and2 I052_1001(w_052_1001, w_043_097, w_028_648);
  or2  I052_1038(w_052_1038, w_003_060, w_018_087);
  not1 I052_1058(w_052_1058, w_007_540);
  or2  I052_1072(w_052_1072, w_036_1140, w_045_1242);
  nand2 I052_1104(w_052_1104, w_021_264, w_005_058);
  not1 I052_1110(w_052_1110, w_025_178);
  nand2 I052_1126(w_052_1126, w_024_220, w_043_040);
  and2 I052_1133(w_052_1133, w_050_105, w_042_051);
  and2 I052_1203(w_052_1203, w_001_129, w_017_681);
  not1 I052_1220(w_052_1220, w_021_191);
  not1 I052_1247(w_052_1247, w_020_538);
  and2 I052_1248(w_052_1248, w_026_1304, w_004_628);
  nand2 I052_1264(w_052_1264, w_001_1126, w_043_077);
  not1 I052_1284(w_052_1284, w_050_1398);
  not1 I052_1289(w_052_1289, w_015_046);
  or2  I052_1295(w_052_1295, w_006_331, w_007_1358);
  or2  I052_1299(w_052_1299, w_002_453, w_012_474);
  not1 I052_1301(w_052_1301, w_047_595);
  not1 I052_1304(w_052_1304, w_038_178);
  not1 I052_1323(w_052_1323, w_042_088);
  and2 I052_1331(w_052_1331, w_024_1053, w_040_1291);
  nand2 I052_1340(w_052_1340, w_008_447, w_003_062);
  not1 I052_1341(w_052_1341, w_050_102);
  nand2 I052_1364(w_052_1364, w_015_082, w_017_264);
  not1 I052_1375(w_052_1375, w_017_1797);
  and2 I052_1379(w_052_1379, w_049_370, w_009_047);
  nand2 I052_1394(w_052_1394, w_006_103, w_049_080);
  or2  I052_1396(w_052_1396, w_002_354, w_038_181);
  nand2 I052_1437(w_052_1437, w_002_462, w_018_216);
  not1 I052_1458(w_052_1458, w_011_678);
  or2  I052_1482(w_052_1482, w_018_119, w_019_487);
  nand2 I052_1525(w_052_1525, w_042_100, w_024_132);
  not1 I052_1549(w_052_1549, w_002_165);
  not1 I052_1554(w_052_1554, w_020_1053);
  or2  I052_1564(w_052_1564, w_020_308, w_014_226);
  not1 I052_1566(w_052_1566, w_019_586);
  or2  I052_1573(w_052_1573, w_043_051, w_036_1153);
  nand2 I052_1588(w_052_1588, w_000_147, w_006_193);
  nand2 I052_1598(w_052_1598, w_017_902, w_050_731);
  nand2 I052_1601(w_052_1601, w_030_811, w_046_231);
  not1 I052_1621(w_052_1621, w_010_146);
  or2  I052_1682(w_052_1682, w_048_787, w_000_662);
  and2 I052_1690(w_052_1690, w_002_328, w_028_287);
  and2 I052_1709(w_052_1709, w_045_1622, w_017_1380);
  or2  I052_1721(w_052_1721, w_009_096, w_021_123);
  nand2 I052_1771(w_052_1771, w_016_034, w_013_163);
  or2  I052_1783(w_052_1783, w_018_189, w_014_218);
  and2 I052_1785(w_052_1785, w_040_212, w_051_673);
  and2 I052_1792(w_052_1792, w_040_055, w_003_047);
  not1 I052_1801(w_052_1801, w_020_439);
  nand2 I052_1844(w_052_1844, w_045_163, w_022_184);
  nand2 I052_1856(w_052_1856, w_011_826, w_007_1231);
  nand2 I052_1875(w_052_1875, w_020_929, w_032_232);
  not1 I052_1907(w_052_1907, w_043_055);
  not1 I052_1918(w_052_1918, w_000_1536);
  and2 I053_000(w_053_000, w_026_846, w_032_021);
  or2  I053_001(w_053_001, w_049_095, w_023_023);
  or2  I053_003(w_053_003, w_018_094, w_006_018);
  not1 I053_004(w_053_004, w_028_465);
  not1 I053_005(w_053_005, w_000_1139);
  and2 I053_007(w_053_007, w_012_035, w_031_1129);
  nand2 I053_011(w_053_011, w_044_1230, w_037_161);
  and2 I053_012(w_053_012, w_037_1406, w_050_020);
  nand2 I053_013(w_053_013, w_035_087, w_034_328);
  nand2 I053_014(w_053_014, w_013_174, w_013_084);
  not1 I053_016(w_053_016, w_001_909);
  and2 I053_017(w_053_017, w_000_1939, w_044_156);
  not1 I053_018(w_053_018, w_014_362);
  or2  I053_019(w_053_019, w_032_231, w_036_1049);
  or2  I053_023(w_053_023, w_029_552, w_027_575);
  not1 I053_024(w_053_024, w_050_181);
  not1 I053_028(w_053_028, w_044_1447);
  not1 I053_029(w_053_029, w_039_087);
  nand2 I053_031(w_053_031, w_013_181, w_025_311);
  and2 I053_032(w_053_032, w_014_164, w_024_064);
  or2  I053_033(w_053_033, w_040_048, w_007_272);
  nand2 I053_034(w_053_034, w_013_080, w_030_795);
  not1 I053_035(w_053_035, w_009_099);
  not1 I053_036(w_053_036, w_033_121);
  or2  I053_040(w_053_040, w_005_598, w_044_357);
  or2  I053_042(w_053_042, w_002_442, w_006_275);
  not1 I053_043(w_053_043, w_040_1084);
  not1 I053_044(w_053_044, w_051_563);
  or2  I053_045(w_053_045, w_037_741, w_052_034);
  and2 I053_047(w_053_047, w_021_058, w_020_599);
  not1 I053_048(w_053_048, w_034_199);
  or2  I053_049(w_053_049, w_027_149, w_050_190);
  nand2 I053_050(w_053_050, w_050_010, w_004_980);
  or2  I053_053(w_053_053, w_036_495, w_044_018);
  nand2 I053_060(w_053_060, w_048_908, w_041_055);
  not1 I053_063(w_053_063, w_022_018);
  or2  I053_064(w_053_064, w_027_552, w_035_238);
  not1 I053_068(w_053_068, w_042_134);
  or2  I053_069(w_053_069, w_043_094, w_049_403);
  and2 I053_071(w_053_071, w_010_083, w_031_229);
  and2 I053_073(w_053_073, w_029_557, w_045_170);
  and2 I053_076(w_053_076, w_029_1170, w_021_134);
  or2  I053_077(w_053_077, w_046_008, w_048_561);
  or2  I053_080(w_053_080, w_050_321, w_006_089);
  not1 I053_083(w_053_083, w_040_044);
  nand2 I053_084(w_053_084, w_033_1142, w_015_249);
  or2  I053_085(w_053_085, w_020_469, w_046_237);
  nand2 I053_087(w_053_087, w_048_781, w_036_161);
  or2  I053_089(w_053_089, w_005_1376, w_032_210);
  or2  I053_091(w_053_091, w_032_155, w_043_020);
  not1 I053_092(w_053_092, w_042_036);
  and2 I053_095(w_053_095, w_048_194, w_020_171);
  not1 I053_096(w_053_096, w_006_019);
  or2  I053_098(w_053_098, w_026_466, w_025_247);
  and2 I053_103(w_053_103, w_027_458, w_008_769);
  nand2 I053_104(w_053_104, w_005_544, w_050_193);
  and2 I053_105(w_053_105, w_027_451, w_002_302);
  or2  I053_106(w_053_106, w_015_050, w_020_1084);
  and2 I053_107(w_053_107, w_014_327, w_034_592);
  nand2 I053_108(w_053_108, w_035_433, w_031_647);
  and2 I053_109(w_053_109, w_043_006, w_034_680);
  not1 I053_110(w_053_110, w_012_196);
  or2  I053_114(w_053_114, w_039_1311, w_052_047);
  not1 I053_116(w_053_116, w_024_692);
  or2  I053_117(w_053_117, w_015_283, w_050_468);
  or2  I053_118(w_053_118, w_031_724, w_000_986);
  or2  I053_120(w_053_120, w_019_417, w_027_218);
  or2  I053_121(w_053_121, w_026_265, w_003_312);
  or2  I054_003(w_054_003, w_037_157, w_050_972);
  or2  I054_007(w_054_007, w_044_1769, w_028_197);
  or2  I054_016(w_054_016, w_043_021, w_020_979);
  not1 I054_036(w_054_036, w_038_108);
  nand2 I054_042(w_054_042, w_007_071, w_037_1441);
  or2  I054_052(w_054_052, w_036_481, w_050_1452);
  and2 I054_057(w_054_057, w_041_018, w_013_080);
  not1 I054_060(w_054_060, w_024_462);
  not1 I054_065(w_054_065, w_019_1074);
  nand2 I054_073(w_054_073, w_012_497, w_042_058);
  nand2 I054_079(w_054_079, w_023_487, w_002_169);
  nand2 I054_086(w_054_086, w_022_251, w_004_022);
  or2  I054_095(w_054_095, w_036_1014, w_052_1001);
  and2 I054_102(w_054_102, w_017_921, w_041_201);
  not1 I054_103(w_054_103, w_041_202);
  not1 I054_117(w_054_117, w_050_1469);
  nand2 I054_158(w_054_158, w_021_007, w_048_597);
  or2  I054_166(w_054_166, w_025_021, w_025_116);
  and2 I054_170(w_054_170, w_022_046, w_032_225);
  nand2 I054_172(w_054_172, w_046_202, w_004_1661);
  nand2 I054_180(w_054_180, w_036_452, w_046_060);
  not1 I054_186(w_054_186, w_015_026);
  and2 I054_188(w_054_188, w_053_003, w_000_583);
  and2 I054_193(w_054_193, w_050_105, w_047_480);
  and2 I054_204(w_054_204, w_022_129, w_036_978);
  or2  I054_220(w_054_220, w_028_384, w_052_017);
  or2  I054_233(w_054_233, w_001_1184, w_017_013);
  nand2 I054_238(w_054_238, w_053_095, w_018_204);
  nand2 I054_251(w_054_251, w_012_369, w_039_1836);
  and2 I054_269(w_054_269, w_040_239, w_046_248);
  not1 I054_275(w_054_275, w_046_267);
  not1 I054_286(w_054_286, w_030_670);
  nand2 I054_299(w_054_299, w_037_355, w_043_064);
  not1 I054_300(w_054_300, w_032_103);
  or2  I054_303(w_054_303, w_034_527, w_001_435);
  and2 I054_308(w_054_308, w_010_128, w_025_719);
  nand2 I054_313(w_054_313, w_011_022, w_020_114);
  not1 I054_315(w_054_315, w_022_038);
  not1 I054_320(w_054_320, w_018_142);
  not1 I054_332(w_054_332, w_011_869);
  nand2 I054_334(w_054_334, w_020_032, w_035_111);
  not1 I054_343(w_054_343, w_031_500);
  not1 I054_352(w_054_352, w_010_403);
  not1 I054_353(w_054_353, w_053_118);
  or2  I054_355(w_054_355, w_010_036, w_006_201);
  nand2 I054_365(w_054_365, w_032_058, w_022_042);
  and2 I054_366(w_054_366, w_026_1026, w_021_248);
  and2 I054_382(w_054_382, w_008_032, w_007_503);
  or2  I054_390(w_054_390, w_010_017, w_000_786);
  not1 I054_399(w_054_399, w_027_028);
  not1 I054_401(w_054_401, w_008_319);
  nand2 I054_411(w_054_411, w_014_821, w_034_201);
  and2 I054_413(w_054_413, w_002_474, w_038_327);
  and2 I054_414(w_054_414, w_025_180, w_043_027);
  or2  I054_432(w_054_432, w_051_285, w_033_1647);
  or2  I054_437(w_054_437, w_023_256, w_011_765);
  nand2 I054_440(w_054_440, w_018_269, w_042_073);
  not1 I054_444(w_054_444, w_018_041);
  and2 I054_469(w_054_469, w_049_020, w_024_1539);
  or2  I054_470(w_054_470, w_003_136, w_027_012);
  not1 I054_477(w_054_477, w_039_199);
  or2  I054_479(w_054_479, w_052_031, w_029_1236);
  and2 I054_482(w_054_482, w_000_236, w_031_587);
  and2 I054_492(w_054_492, w_047_345, w_014_717);
  and2 I054_499(w_054_499, w_038_390, w_045_495);
  or2  I054_508(w_054_508, w_015_080, w_012_375);
  or2  I054_509(w_054_509, w_029_1272, w_001_1105);
  not1 I054_518(w_054_518, w_027_114);
  not1 I054_532(w_054_532, w_042_009);
  nand2 I054_535(w_054_535, w_029_628, w_032_234);
  not1 I054_537(w_054_537, w_035_1335);
  nand2 I054_540(w_054_540, w_015_210, w_005_243);
  and2 I054_544(w_054_544, w_036_723, w_018_005);
  and2 I054_546(w_054_546, w_031_456, w_025_592);
  nand2 I054_549(w_054_549, w_053_114, w_012_400);
  and2 I054_553(w_054_553, w_002_226, w_033_294);
  and2 I054_570(w_054_570, w_020_228, w_016_012);
  nand2 I054_572(w_054_572, w_015_041, w_020_278);
  or2  I054_577(w_054_577, w_042_025, w_053_000);
  and2 I054_578(w_054_578, w_017_1351, w_038_181);
  not1 I054_579(w_054_579, w_009_094);
  and2 I054_581(w_054_581, w_050_342, w_035_644);
  and2 I054_592(w_054_592, w_029_273, w_009_088);
  nand2 I054_596(w_054_596, w_022_061, w_046_223);
  nand2 I054_599(w_054_599, w_022_118, w_027_041);
  not1 I054_606(w_054_606, w_011_007);
  nand2 I054_618(w_054_618, w_004_1667, w_031_852);
  not1 I054_620(w_054_620, w_021_221);
  or2  I054_627(w_054_629, w_049_1169, w_054_628);
  nand2 I054_628(w_054_630, w_054_629, w_022_068);
  not1 I054_629(w_054_631, w_054_630);
  or2  I054_630(w_054_632, w_016_013, w_054_631);
  not1 I054_631(w_054_633, w_054_632);
  not1 I054_632(w_054_634, w_054_633);
  not1 I054_633(w_054_635, w_054_634);
  or2  I054_634(w_054_636, w_025_556, w_054_635);
  not1 I054_635(w_054_637, w_054_636);
  or2  I054_636(w_054_628, w_018_276, w_054_637);
  or2  I055_001(w_055_001, w_025_1134, w_050_090);
  and2 I055_005(w_055_005, w_014_171, w_015_264);
  not1 I055_007(w_055_007, w_046_198);
  or2  I055_012(w_055_012, w_030_780, w_028_150);
  or2  I055_021(w_055_021, w_051_026, w_038_391);
  and2 I055_023(w_055_023, w_001_1665, w_012_144);
  or2  I055_036(w_055_036, w_041_201, w_020_430);
  or2  I055_044(w_055_044, w_009_083, w_001_907);
  nand2 I055_053(w_055_053, w_002_351, w_015_040);
  not1 I055_057(w_055_057, w_027_183);
  or2  I055_061(w_055_061, w_032_118, w_022_217);
  not1 I055_076(w_055_076, w_012_357);
  not1 I055_087(w_055_087, w_051_847);
  not1 I055_090(w_055_090, w_054_193);
  or2  I055_094(w_055_094, w_042_100, w_031_349);
  or2  I055_100(w_055_100, w_051_633, w_050_556);
  not1 I055_104(w_055_104, w_017_1449);
  not1 I055_109(w_055_109, w_003_127);
  nand2 I055_111(w_055_111, w_018_194, w_053_085);
  not1 I055_113(w_055_113, w_042_031);
  and2 I055_123(w_055_123, w_035_1227, w_019_317);
  not1 I055_128(w_055_128, w_028_813);
  and2 I055_148(w_055_148, w_054_158, w_047_640);
  not1 I055_149(w_055_149, w_025_914);
  nand2 I055_154(w_055_154, w_007_1605, w_008_821);
  not1 I055_155(w_055_155, w_013_038);
  and2 I055_157(w_055_157, w_047_224, w_009_098);
  or2  I055_160(w_055_160, w_033_221, w_029_332);
  or2  I055_162(w_055_162, w_043_011, w_029_962);
  not1 I055_164(w_055_164, w_041_053);
  or2  I055_167(w_055_167, w_049_620, w_012_567);
  nand2 I055_169(w_055_169, w_043_065, w_001_457);
  not1 I055_170(w_055_170, w_040_673);
  nand2 I055_173(w_055_173, w_042_128, w_049_327);
  or2  I055_181(w_055_181, w_002_327, w_004_491);
  and2 I055_213(w_055_213, w_040_320, w_042_002);
  not1 I055_214(w_055_214, w_022_339);
  not1 I055_216(w_055_216, w_020_784);
  or2  I055_220(w_055_220, w_041_069, w_042_030);
  or2  I055_226(w_055_226, w_050_749, w_022_325);
  nand2 I055_232(w_055_232, w_015_016, w_047_301);
  not1 I055_233(w_055_233, w_031_820);
  not1 I055_242(w_055_242, w_047_251);
  or2  I055_243(w_055_243, w_041_273, w_023_764);
  nand2 I055_245(w_055_245, w_021_275, w_046_052);
  or2  I055_253(w_055_253, w_044_794, w_040_060);
  or2  I055_254(w_055_254, w_035_109, w_050_764);
  not1 I055_259(w_055_259, w_026_993);
  nand2 I055_260(w_055_260, w_002_005, w_049_529);
  and2 I055_261(w_055_261, w_017_432, w_004_1886);
  or2  I055_284(w_055_284, w_054_414, w_038_100);
  nand2 I055_291(w_055_291, w_014_326, w_038_439);
  and2 I055_292(w_055_292, w_034_300, w_023_066);
  nand2 I055_300(w_055_300, w_039_714, w_015_153);
  not1 I055_306(w_055_306, w_001_948);
  not1 I055_311(w_055_311, w_019_757);
  not1 I055_324(w_055_324, w_019_527);
  and2 I055_325(w_055_325, w_014_235, w_011_155);
  not1 I055_327(w_055_327, w_050_101);
  not1 I055_335(w_055_335, w_011_534);
  nand2 I055_339(w_055_339, w_036_025, w_005_722);
  and2 I055_361(w_055_361, w_009_094, w_031_827);
  nand2 I055_363(w_055_363, w_041_249, w_010_057);
  nand2 I055_370(w_055_370, w_050_499, w_042_117);
  or2  I055_373(w_055_373, w_053_098, w_042_128);
  and2 I055_382(w_055_382, w_028_076, w_011_541);
  and2 I055_385(w_055_385, w_050_751, w_031_457);
  and2 I055_389(w_055_389, w_018_128, w_004_862);
  not1 I055_420(w_055_420, w_000_894);
  or2  I055_421(w_055_421, w_046_215, w_025_697);
  not1 I055_422(w_055_422, w_022_030);
  not1 I055_423(w_055_423, w_015_199);
  or2  I055_435(w_055_435, w_009_029, w_018_050);
  or2  I055_443(w_055_443, w_037_085, w_029_718);
  nand2 I055_466(w_055_466, w_051_649, w_051_992);
  nand2 I055_469(w_055_469, w_028_189, w_013_176);
  not1 I055_473(w_055_473, w_005_1160);
  nand2 I055_475(w_055_475, w_030_159, w_042_105);
  not1 I055_494(w_055_494, w_010_117);
  nand2 I055_525(w_055_525, w_014_271, w_048_077);
  and2 I055_526(w_055_526, w_040_030, w_001_209);
  not1 I055_567(w_055_567, w_020_209);
  and2 I055_576(w_055_576, w_021_134, w_024_735);
  and2 I055_590(w_055_590, w_050_015, w_006_151);
  or2  I055_594(w_055_594, w_009_047, w_044_788);
  not1 I055_598(w_055_598, w_021_024);
  nand2 I055_602(w_055_602, w_011_455, w_023_100);
  not1 I055_604(w_055_604, w_053_000);
  not1 I055_610(w_055_610, w_032_158);
  or2  I055_636(w_055_636, w_027_301, w_036_813);
  and2 I055_647(w_055_647, w_006_194, w_048_229);
  and2 I055_650(w_055_650, w_048_447, w_026_467);
  or2  I055_660(w_055_660, w_009_105, w_044_308);
  not1 I055_661(w_055_661, w_011_546);
  nand2 I055_671(w_055_671, w_000_1216, w_048_802);
  and2 I055_672(w_055_672, w_029_133, w_007_208);
  and2 I055_693(w_055_693, w_049_548, w_009_027);
  not1 I055_715(w_055_715, w_012_486);
  and2 I055_716(w_055_716, w_016_033, w_009_071);
  not1 I055_717(w_055_717, w_020_742);
  or2  I055_735(w_055_735, w_021_145, w_004_1562);
  not1 I055_744(w_055_744, w_025_035);
  nand2 I055_750(w_055_750, w_048_054, w_052_1437);
  or2  I055_772(w_055_772, w_024_895, w_032_126);
  or2  I055_775(w_055_775, w_009_055, w_007_1138);
  or2  I055_786(w_055_786, w_005_220, w_017_225);
  or2  I055_821(w_055_821, w_012_304, w_041_049);
  and2 I055_828(w_055_828, w_032_045, w_042_140);
  or2  I055_835(w_055_835, w_032_065, w_010_290);
  not1 I055_852(w_055_852, w_013_179);
  and2 I055_856(w_055_856, w_005_1058, w_024_1640);
  and2 I056_000(w_056_000, w_044_914, w_044_790);
  and2 I056_018(w_056_018, w_019_783, w_023_329);
  or2  I056_020(w_056_020, w_021_049, w_046_219);
  or2  I056_023(w_056_023, w_044_1769, w_007_666);
  and2 I056_033(w_056_033, w_020_983, w_050_1383);
  not1 I056_085(w_056_085, w_054_315);
  and2 I056_086(w_056_086, w_034_330, w_039_835);
  nand2 I056_112(w_056_112, w_052_1299, w_027_417);
  or2  I056_114(w_056_114, w_023_758, w_007_218);
  not1 I056_124(w_056_124, w_010_229);
  and2 I056_125(w_056_125, w_016_037, w_020_007);
  or2  I056_161(w_056_161, w_044_1379, w_021_088);
  nand2 I056_164(w_056_164, w_028_158, w_034_471);
  and2 I056_165(w_056_165, w_014_212, w_014_205);
  not1 I056_178(w_056_178, w_030_065);
  not1 I056_182(w_056_182, w_055_021);
  not1 I056_192(w_056_192, w_010_197);
  or2  I056_193(w_056_193, w_004_115, w_006_163);
  and2 I056_196(w_056_196, w_014_772, w_031_576);
  not1 I056_203(w_056_203, w_032_102);
  or2  I056_211(w_056_211, w_042_130, w_049_043);
  nand2 I056_217(w_056_217, w_046_077, w_007_1097);
  nand2 I056_231(w_056_231, w_050_418, w_051_714);
  not1 I056_233(w_056_233, w_008_352);
  and2 I056_246(w_056_246, w_038_134, w_055_382);
  not1 I056_251(w_056_251, w_055_214);
  or2  I056_254(w_056_254, w_010_163, w_015_073);
  nand2 I056_273(w_056_273, w_029_188, w_024_003);
  nand2 I056_298(w_056_298, w_043_081, w_003_235);
  not1 I056_315(w_056_315, w_052_1682);
  or2  I056_333(w_056_333, w_033_1015, w_006_299);
  or2  I056_382(w_056_382, w_028_847, w_048_884);
  and2 I056_411(w_056_411, w_030_591, w_025_759);
  or2  I056_441(w_056_441, w_034_382, w_045_1104);
  or2  I056_492(w_056_492, w_013_092, w_004_481);
  not1 I056_503(w_056_503, w_040_325);
  nand2 I056_504(w_056_504, w_033_175, w_005_273);
  not1 I056_512(w_056_512, w_037_900);
  and2 I056_519(w_056_519, w_053_117, w_052_1525);
  not1 I056_589(w_056_589, w_031_853);
  or2  I056_615(w_056_615, w_000_079, w_002_001);
  nand2 I056_625(w_056_625, w_006_087, w_028_018);
  not1 I056_637(w_056_637, w_013_127);
  nand2 I056_650(w_056_650, w_000_1700, w_002_206);
  and2 I056_658(w_056_658, w_046_230, w_048_213);
  or2  I056_659(w_056_659, w_024_1466, w_003_225);
  nand2 I056_668(w_056_668, w_004_1302, w_015_019);
  nand2 I056_679(w_056_679, w_008_443, w_052_440);
  or2  I056_717(w_056_717, w_013_172, w_013_107);
  not1 I056_727(w_056_727, w_049_433);
  not1 I056_745(w_056_745, w_044_1116);
  or2  I056_751(w_056_751, w_007_953, w_036_283);
  not1 I056_795(w_056_795, w_017_1240);
  and2 I056_800(w_056_800, w_028_108, w_024_201);
  and2 I056_810(w_056_810, w_040_227, w_043_055);
  nand2 I056_821(w_056_821, w_020_507, w_004_1871);
  not1 I056_830(w_056_830, w_008_720);
  and2 I056_833(w_056_833, w_010_064, w_004_1388);
  and2 I056_835(w_056_835, w_036_207, w_012_105);
  or2  I056_876(w_056_876, w_005_309, w_043_062);
  nand2 I056_890(w_056_890, w_001_1248, w_015_065);
  and2 I056_894(w_056_894, w_025_106, w_013_103);
  nand2 I056_928(w_056_928, w_049_311, w_042_100);
  not1 I056_929(w_056_929, w_009_102);
  or2  I056_936(w_056_936, w_054_186, w_029_133);
  and2 I056_972(w_056_972, w_030_349, w_053_042);
  and2 I056_980(w_056_980, w_053_084, w_047_259);
  and2 I056_1064(w_056_1064, w_039_482, w_002_249);
  nand2 I056_1109(w_056_1109, w_032_180, w_038_058);
  or2  I056_1115(w_056_1115, w_003_084, w_012_620);
  not1 I056_1121(w_056_1121, w_019_968);
  or2  I056_1172(w_056_1172, w_020_288, w_033_845);
  or2  I056_1176(w_056_1176, w_016_011, w_006_125);
  and2 I056_1184(w_056_1184, w_054_275, w_002_344);
  nand2 I056_1223(w_056_1223, w_042_022, w_009_086);
  and2 I056_1229(w_056_1229, w_040_052, w_004_1326);
  or2  I056_1269(w_056_1269, w_006_323, w_013_029);
  not1 I056_1275(w_056_1275, w_012_338);
  not1 I056_1290(w_056_1290, w_038_152);
  nand2 I056_1315(w_056_1315, w_002_558, w_033_323);
  not1 I056_1342(w_056_1342, w_044_1152);
  and2 I056_1363(w_056_1363, w_006_100, w_006_277);
  nand2 I056_1388(w_056_1388, w_025_255, w_000_300);
  nand2 I056_1391(w_056_1391, w_004_1823, w_025_1047);
  and2 I056_1409(w_056_1409, w_020_330, w_009_021);
  not1 I056_1424(w_056_1424, w_052_1690);
  nand2 I056_1446(w_056_1446, w_019_675, w_050_1379);
  and2 I056_1460(w_056_1460, w_008_489, w_007_873);
  nand2 I056_1465(w_056_1465, w_009_091, w_032_066);
  or2  I056_1468(w_056_1468, w_051_621, w_049_542);
  or2  I056_1502(w_056_1502, w_003_190, w_052_1331);
  and2 I056_1511(w_056_1511, w_019_695, w_027_429);
  or2  I056_1534(w_056_1534, w_030_845, w_024_143);
  or2  I056_1537(w_056_1537, w_003_175, w_030_559);
  nand2 I056_1540(w_056_1540, w_012_235, w_041_235);
  nand2 I056_1562(w_056_1562, w_023_1348, w_010_065);
  not1 I056_1615(w_056_1615, w_054_303);
  not1 I056_1623(w_056_1623, w_038_287);
  or2  I056_1651(w_056_1651, w_047_115, w_040_1038);
  or2  I056_1671(w_056_1671, w_043_020, w_033_1409);
  not1 I057_025(w_057_025, w_004_258);
  not1 I057_034(w_057_034, w_053_049);
  and2 I057_037(w_057_037, w_054_413, w_036_1234);
  and2 I057_058(w_057_058, w_042_035, w_011_654);
  and2 I057_105(w_057_105, w_002_509, w_028_140);
  not1 I057_137(w_057_137, w_001_1629);
  or2  I057_145(w_057_145, w_003_279, w_022_135);
  and2 I057_177(w_057_177, w_026_952, w_018_264);
  not1 I057_186(w_057_186, w_034_125);
  not1 I057_190(w_057_190, w_023_1262);
  not1 I057_209(w_057_209, w_013_328);
  nand2 I057_222(w_057_222, w_006_243, w_055_123);
  not1 I057_225(w_057_225, w_009_013);
  or2  I057_228(w_057_228, w_040_020, w_002_428);
  and2 I057_233(w_057_233, w_009_052, w_017_1145);
  and2 I057_239(w_057_239, w_023_227, w_025_1408);
  or2  I057_240(w_057_240, w_001_905, w_003_069);
  or2  I057_250(w_057_250, w_031_260, w_026_567);
  and2 I057_276(w_057_276, w_004_326, w_029_394);
  nand2 I057_277(w_057_277, w_015_198, w_014_172);
  nand2 I057_284(w_057_284, w_052_1792, w_007_518);
  nand2 I057_298(w_057_298, w_029_970, w_028_801);
  and2 I057_330(w_057_330, w_027_482, w_018_153);
  not1 I057_369(w_057_369, w_017_010);
  and2 I057_399(w_057_399, w_031_016, w_039_847);
  and2 I057_413(w_057_413, w_001_1353, w_050_257);
  and2 I057_430(w_057_430, w_029_532, w_027_214);
  not1 I057_454(w_057_454, w_012_635);
  nand2 I057_487(w_057_487, w_005_551, w_056_193);
  or2  I057_516(w_057_516, w_032_073, w_004_1793);
  and2 I057_551(w_057_551, w_008_485, w_002_528);
  or2  I057_592(w_057_592, w_009_006, w_011_273);
  or2  I057_606(w_057_606, w_046_011, w_018_004);
  or2  I057_632(w_057_632, w_025_202, w_047_065);
  or2  I057_645(w_057_645, w_010_098, w_029_756);
  and2 I057_653(w_057_653, w_000_342, w_032_039);
  nand2 I057_660(w_057_660, w_046_216, w_053_005);
  and2 I057_676(w_057_676, w_039_507, w_009_004);
  and2 I057_709(w_057_709, w_056_020, w_019_559);
  nand2 I057_743(w_057_743, w_005_1098, w_009_049);
  not1 I057_790(w_057_790, w_005_123);
  nand2 I057_816(w_057_816, w_013_299, w_022_139);
  not1 I057_828(w_057_828, w_044_1459);
  nand2 I057_829(w_057_829, w_044_1274, w_000_496);
  or2  I057_832(w_057_832, w_037_1320, w_019_505);
  and2 I057_854(w_057_854, w_009_066, w_036_496);
  nand2 I057_857(w_057_857, w_037_160, w_053_045);
  nand2 I057_861(w_057_861, w_027_160, w_050_016);
  not1 I057_883(w_057_883, w_046_014);
  and2 I057_915(w_057_915, w_055_181, w_019_164);
  and2 I057_928(w_057_928, w_008_477, w_022_295);
  nand2 I057_936(w_057_936, w_052_059, w_054_238);
  not1 I057_983(w_057_983, w_033_1489);
  and2 I057_984(w_057_984, w_046_121, w_034_201);
  nand2 I057_1003(w_057_1003, w_054_079, w_005_1106);
  nand2 I057_1031(w_057_1031, w_022_085, w_029_904);
  or2  I057_1038(w_057_1038, w_009_075, w_036_147);
  or2  I057_1047(w_057_1047, w_013_168, w_025_240);
  not1 I057_1060(w_057_1060, w_000_290);
  and2 I057_1103(w_057_1103, w_056_1537, w_031_625);
  not1 I057_1124(w_057_1124, w_031_226);
  or2  I057_1156(w_057_1156, w_032_175, w_043_029);
  and2 I057_1158(w_057_1158, w_037_884, w_000_1560);
  not1 I057_1166(w_057_1166, w_046_238);
  not1 I057_1174(w_057_1174, w_002_505);
  and2 I057_1216(w_057_1216, w_028_022, w_043_056);
  or2  I057_1249(w_057_1249, w_017_234, w_047_606);
  or2  I057_1252(w_057_1252, w_010_324, w_000_1427);
  nand2 I057_1266(w_057_1266, w_008_678, w_029_307);
  or2  I057_1301(w_057_1301, w_015_255, w_025_1161);
  not1 I057_1307(w_057_1307, w_009_031);
  nand2 I057_1337(w_057_1337, w_005_076, w_022_000);
  or2  I057_1351(w_057_1351, w_018_124, w_023_1410);
  and2 I057_1360(w_057_1360, w_027_436, w_042_008);
  nand2 I057_1410(w_057_1410, w_051_202, w_010_291);
  nand2 I057_1414(w_057_1414, w_000_1863, w_041_198);
  and2 I057_1445(w_057_1445, w_047_013, w_048_057);
  nand2 I057_1467(w_057_1467, w_023_211, w_037_535);
  not1 I057_1517(w_057_1517, w_033_1187);
  or2  I057_1525(w_057_1525, w_020_1120, w_006_138);
  or2  I057_1536(w_057_1536, w_003_043, w_026_1357);
  and2 I057_1562(w_057_1562, w_023_255, w_029_715);
  or2  I057_1591(w_057_1591, w_047_545, w_040_495);
  nand2 I057_1599(w_057_1599, w_043_029, w_053_028);
  and2 I057_1600(w_057_1600, w_023_1439, w_013_274);
  not1 I057_1605(w_057_1605, w_026_201);
  and2 I057_1615(w_057_1615, w_027_584, w_027_456);
  or2  I057_1646(w_057_1646, w_043_032, w_044_1630);
  or2  I057_1717(w_057_1717, w_051_812, w_036_114);
  nand2 I057_1740(w_057_1740, w_050_045, w_008_222);
  nand2 I057_1768(w_057_1768, w_004_223, w_056_182);
  and2 I057_1817(w_057_1817, w_056_972, w_049_813);
  not1 I057_1838(w_057_1838, w_041_098);
  nand2 I058_011(w_058_011, w_046_054, w_019_488);
  not1 I058_025(w_058_025, w_047_000);
  or2  I058_034(w_058_034, w_022_327, w_042_052);
  nand2 I058_038(w_058_038, w_051_382, w_016_014);
  or2  I058_041(w_058_041, w_036_199, w_021_155);
  nand2 I058_054(w_058_054, w_002_289, w_047_062);
  nand2 I058_058(w_058_058, w_009_081, w_035_1125);
  and2 I058_064(w_058_064, w_019_625, w_026_331);
  or2  I058_074(w_058_074, w_024_1105, w_005_053);
  nand2 I058_080(w_058_080, w_035_678, w_027_199);
  or2  I058_097(w_058_097, w_021_262, w_019_191);
  not1 I058_108(w_058_108, w_052_1875);
  nand2 I058_125(w_058_125, w_033_1214, w_042_035);
  not1 I058_147(w_058_147, w_039_775);
  not1 I058_174(w_058_174, w_000_687);
  not1 I058_186(w_058_186, w_040_463);
  and2 I058_190(w_058_190, w_045_830, w_047_140);
  nand2 I058_196(w_058_196, w_015_035, w_003_149);
  not1 I058_199(w_058_199, w_023_1607);
  or2  I058_203(w_058_203, w_040_984, w_014_545);
  or2  I058_212(w_058_212, w_054_382, w_004_994);
  or2  I058_220(w_058_220, w_028_189, w_031_306);
  not1 I058_240(w_058_240, w_057_190);
  not1 I058_242(w_058_242, w_019_890);
  nand2 I058_266(w_058_266, w_050_462, w_014_533);
  not1 I058_302(w_058_302, w_032_103);
  nand2 I058_315(w_058_315, w_041_096, w_047_074);
  or2  I058_360(w_058_360, w_028_025, w_016_032);
  or2  I058_367(w_058_367, w_033_103, w_029_187);
  or2  I058_392(w_058_392, w_053_071, w_049_1169);
  and2 I058_403(w_058_403, w_041_205, w_056_717);
  or2  I058_415(w_058_415, w_004_068, w_022_400);
  and2 I058_431(w_058_431, w_027_552, w_042_093);
  or2  I058_436(w_058_436, w_004_545, w_000_1727);
  not1 I058_459(w_058_459, w_028_557);
  and2 I058_481(w_058_481, w_007_258, w_040_324);
  and2 I058_498(w_058_498, w_016_021, w_000_954);
  or2  I058_521(w_058_521, w_029_020, w_018_267);
  or2  I058_531(w_058_531, w_006_087, w_054_269);
  nand2 I058_533(w_058_533, w_033_413, w_026_388);
  and2 I058_553(w_058_553, w_020_397, w_057_1740);
  and2 I058_589(w_058_589, w_046_276, w_021_167);
  nand2 I058_608(w_058_608, w_031_515, w_002_410);
  nand2 I058_616(w_058_616, w_045_1718, w_050_191);
  nand2 I058_625(w_058_625, w_014_129, w_006_132);
  not1 I058_649(w_058_649, w_000_703);
  not1 I058_701(w_058_701, w_046_005);
  and2 I058_732(w_058_732, w_053_023, w_020_464);
  and2 I058_743(w_058_743, w_049_311, w_010_114);
  or2  I058_762(w_058_762, w_035_088, w_017_1588);
  not1 I058_768(w_058_768, w_032_187);
  or2  I058_780(w_058_780, w_018_109, w_039_629);
  not1 I058_794(w_058_794, w_052_1801);
  and2 I058_809(w_058_809, w_013_073, w_032_199);
  not1 I058_814(w_058_814, w_043_036);
  nand2 I058_822(w_058_822, w_018_040, w_036_079);
  or2  I058_828(w_058_828, w_053_121, w_024_830);
  and2 I058_840(w_058_840, w_004_934, w_003_051);
  nand2 I058_843(w_058_843, w_026_785, w_007_1538);
  or2  I058_875(w_058_875, w_014_805, w_018_037);
  and2 I058_885(w_058_885, w_025_289, w_024_1362);
  not1 I058_891(w_058_891, w_018_263);
  nand2 I058_919(w_058_919, w_010_116, w_003_241);
  not1 I058_935(w_058_935, w_010_063);
  and2 I058_938(w_058_938, w_020_183, w_026_065);
  nand2 I058_955(w_058_955, w_015_071, w_051_108);
  nand2 I058_961(w_058_961, w_011_691, w_017_003);
  not1 I058_1006(w_058_1006, w_042_107);
  nand2 I058_1019(w_058_1019, w_009_048, w_012_509);
  nand2 I058_1023(w_058_1023, w_025_1537, w_051_230);
  or2  I058_1027(w_058_1027, w_007_640, w_007_415);
  and2 I058_1033(w_058_1033, w_055_775, w_011_670);
  and2 I058_1040(w_058_1040, w_017_482, w_022_113);
  not1 I058_1050(w_058_1050, w_041_021);
  nand2 I058_1064(w_058_1064, w_051_1023, w_022_311);
  or2  I058_1086(w_058_1086, w_025_592, w_053_114);
  nand2 I058_1121(w_058_1121, w_034_669, w_031_425);
  nand2 I058_1144(w_058_1144, w_022_235, w_026_997);
  not1 I058_1145(w_058_1145, w_047_190);
  nand2 I058_1146(w_058_1146, w_021_223, w_016_031);
  nand2 I058_1160(w_058_1160, w_013_093, w_024_218);
  or2  I058_1169(w_058_1169, w_022_373, w_025_1611);
  or2  I058_1187(w_058_1187, w_031_246, w_055_173);
  not1 I058_1190(w_058_1190, w_031_398);
  or2  I058_1220(w_058_1220, w_031_289, w_000_1725);
  and2 I058_1236(w_058_1236, w_015_186, w_002_032);
  nand2 I058_1255(w_058_1255, w_018_007, w_046_048);
  nand2 I058_1291(w_058_1291, w_039_007, w_026_1126);
  or2  I058_1294(w_058_1294, w_013_031, w_048_487);
  nand2 I058_1300(w_058_1300, w_014_020, w_019_543);
  or2  I058_1346(w_058_1346, w_015_039, w_000_1227);
  not1 I058_1347(w_058_1347, w_007_317);
  or2  I058_1412(w_058_1412, w_022_088, w_014_825);
  nand2 I058_1424(w_058_1424, w_018_141, w_027_288);
  nand2 I058_1469(w_058_1469, w_017_1563, w_020_030);
  and2 I058_1473(w_058_1473, w_048_824, w_041_042);
  nand2 I058_1478(w_058_1478, w_004_1121, w_034_305);
  nand2 I058_1485(w_058_1485, w_037_143, w_037_1625);
  nand2 I058_1500(w_058_1500, w_037_508, w_012_110);
  nand2 I058_1589(w_058_1589, w_021_027, w_039_834);
  or2  I058_1606(w_058_1606, w_053_073, w_052_1601);
  and2 I058_1624(w_058_1624, w_054_353, w_051_670);
  or2  I058_1629(w_058_1629, w_027_578, w_042_063);
  and2 I058_1630(w_058_1630, w_047_073, w_050_175);
  not1 I058_1712(w_058_1712, w_007_283);
  not1 I058_1721(w_058_1721, w_005_811);
  nand2 I058_1743(w_058_1743, w_040_1046, w_023_585);
  not1 I058_1762(w_058_1762, w_010_309);
  not1 I058_1779(w_058_1779, w_012_506);
  and2 I059_008(w_059_008, w_021_225, w_058_481);
  or2  I059_014(w_059_014, w_003_305, w_025_1070);
  nand2 I059_017(w_059_017, w_001_1394, w_041_037);
  or2  I059_020(w_059_020, w_005_269, w_004_1108);
  nand2 I059_023(w_059_023, w_026_423, w_055_245);
  or2  I059_042(w_059_042, w_031_279, w_044_795);
  not1 I059_052(w_059_052, w_054_437);
  nand2 I059_059(w_059_059, w_051_982, w_036_405);
  or2  I059_065(w_059_065, w_010_073, w_027_558);
  not1 I059_080(w_059_080, w_042_079);
  or2  I059_082(w_059_082, w_041_208, w_018_081);
  and2 I059_084(w_059_084, w_048_554, w_039_793);
  not1 I059_093(w_059_093, w_002_043);
  not1 I059_096(w_059_096, w_058_240);
  nand2 I059_113(w_059_113, w_051_628, w_058_935);
  or2  I059_117(w_059_117, w_034_007, w_000_1371);
  and2 I059_125(w_059_125, w_018_056, w_001_827);
  and2 I059_127(w_059_127, w_020_846, w_025_941);
  nand2 I059_139(w_059_139, w_007_525, w_051_837);
  nand2 I059_152(w_059_152, w_047_503, w_043_012);
  nand2 I059_158(w_059_158, w_040_093, w_052_391);
  or2  I059_165(w_059_165, w_038_012, w_042_139);
  not1 I059_172(w_059_172, w_042_051);
  nand2 I059_175(w_059_175, w_033_082, w_056_1409);
  and2 I059_179(w_059_179, w_050_1319, w_033_1291);
  nand2 I059_183(w_059_183, w_016_037, w_004_1798);
  and2 I059_184(w_059_184, w_014_815, w_045_452);
  and2 I059_206(w_059_206, w_049_169, w_000_1250);
  not1 I059_207(w_059_207, w_031_003);
  and2 I059_210(w_059_210, w_053_109, w_028_380);
  nand2 I059_214(w_059_214, w_022_148, w_028_453);
  not1 I059_228(w_059_228, w_021_194);
  not1 I059_229(w_059_229, w_022_392);
  and2 I059_246(w_059_246, w_025_1675, w_029_754);
  nand2 I059_272(w_059_272, w_053_005, w_008_380);
  nand2 I059_278(w_059_278, w_057_225, w_037_812);
  nand2 I059_284(w_059_284, w_023_1037, w_031_116);
  not1 I059_288(w_059_288, w_012_122);
  and2 I059_289(w_059_289, w_020_485, w_058_828);
  and2 I059_293(w_059_293, w_020_422, w_000_1924);
  nand2 I059_296(w_059_296, w_008_449, w_032_126);
  and2 I059_298(w_059_298, w_024_1591, w_048_637);
  and2 I059_303(w_059_303, w_055_420, w_039_1078);
  or2  I059_318(w_059_318, w_056_833, w_037_553);
  or2  I059_333(w_059_333, w_026_148, w_004_254);
  and2 I059_344(w_059_344, w_004_677, w_040_1082);
  not1 I059_346(w_059_346, w_049_315);
  or2  I059_353(w_059_353, w_007_1097, w_017_1814);
  nand2 I059_360(w_059_360, w_007_547, w_044_1580);
  not1 I059_361(w_059_361, w_038_141);
  not1 I059_381(w_059_381, w_015_223);
  or2  I059_383(w_059_383, w_040_539, w_040_1156);
  nand2 I059_395(w_059_395, w_023_262, w_032_029);
  and2 I059_403(w_059_403, w_008_579, w_001_879);
  not1 I059_429(w_059_429, w_037_1554);
  nand2 I059_435(w_059_435, w_000_219, w_022_222);
  or2  I059_445(w_059_445, w_023_956, w_033_018);
  or2  I059_450(w_059_450, w_034_563, w_030_677);
  not1 I059_457(w_059_457, w_037_1309);
  nand2 I059_463(w_059_463, w_048_243, w_042_008);
  and2 I059_478(w_059_478, w_052_1564, w_035_936);
  and2 I059_482(w_059_482, w_046_049, w_058_1473);
  not1 I059_485(w_059_485, w_020_614);
  and2 I059_489(w_059_489, w_029_516, w_008_830);
  or2  I059_492(w_059_492, w_016_014, w_049_013);
  and2 I059_497(w_059_497, w_048_171, w_021_179);
  or2  I059_503(w_059_503, w_049_1006, w_000_627);
  not1 I059_509(w_059_509, w_026_266);
  nand2 I059_518(w_059_518, w_010_045, w_053_080);
  and2 I059_549(w_059_549, w_043_058, w_043_046);
  and2 I059_561(w_059_561, w_050_033, w_021_136);
  and2 I059_565(w_059_565, w_007_785, w_006_315);
  not1 I059_572(w_059_572, w_004_1207);
  or2  I059_573(w_059_573, w_057_413, w_020_138);
  and2 I059_577(w_059_577, w_019_353, w_058_762);
  nand2 I059_597(w_059_597, w_024_260, w_034_089);
  and2 I059_599(w_059_599, w_021_049, w_017_1153);
  nand2 I059_606(w_059_606, w_005_665, w_028_409);
  not1 I059_608(w_059_608, w_028_526);
  and2 I059_619(w_059_619, w_052_877, w_048_799);
  and2 I059_622(w_059_622, w_044_1616, w_030_072);
  and2 I059_632(w_059_632, w_024_336, w_042_121);
  and2 I059_651(w_059_651, w_019_077, w_022_177);
  nand2 I059_653(w_059_653, w_012_435, w_028_516);
  and2 I059_692(w_059_692, w_040_526, w_048_694);
  nand2 I060_003(w_060_003, w_038_158, w_044_907);
  nand2 I060_005(w_060_005, w_053_121, w_035_1621);
  and2 I060_006(w_060_006, w_055_385, w_004_407);
  and2 I060_007(w_060_007, w_021_026, w_034_216);
  nand2 I060_009(w_060_009, w_029_887, w_048_000);
  nand2 I060_010(w_060_010, w_026_1002, w_007_526);
  and2 I060_011(w_060_011, w_050_671, w_047_303);
  not1 I060_012(w_060_012, w_015_276);
  nand2 I060_013(w_060_013, w_010_171, w_011_077);
  not1 I060_016(w_060_016, w_043_098);
  not1 I060_018(w_060_018, w_026_871);
  not1 I060_019(w_060_019, w_001_489);
  or2  I060_020(w_060_020, w_057_1124, w_051_022);
  nand2 I060_022(w_060_022, w_044_1635, w_026_099);
  not1 I060_024(w_060_024, w_059_497);
  and2 I060_025(w_060_025, w_018_162, w_008_444);
  or2  I060_026(w_060_026, w_019_269, w_014_436);
  and2 I060_028(w_060_028, w_023_914, w_048_904);
  or2  I060_029(w_060_029, w_025_171, w_055_604);
  nand2 I060_030(w_060_030, w_038_333, w_021_124);
  nand2 I060_031(w_060_031, w_021_220, w_021_231);
  and2 I060_032(w_060_032, w_034_400, w_015_113);
  and2 I060_033(w_060_033, w_026_175, w_037_1489);
  nand2 I060_034(w_060_034, w_042_068, w_013_242);
  or2  I060_035(w_060_035, w_050_225, w_018_160);
  not1 I060_037(w_060_037, w_015_237);
  not1 I060_038(w_060_038, w_029_1328);
  nand2 I060_039(w_060_039, w_003_080, w_026_366);
  and2 I060_040(w_060_040, w_052_011, w_030_623);
  or2  I060_041(w_060_041, w_004_1485, w_006_322);
  nand2 I060_046(w_060_046, w_033_022, w_055_292);
  and2 I060_047(w_060_047, w_025_999, w_013_161);
  or2  I060_052(w_060_052, w_029_1127, w_048_373);
  not1 I060_053(w_060_053, w_043_032);
  not1 I060_054(w_060_054, w_001_190);
  nand2 I060_055(w_060_055, w_022_278, w_038_170);
  or2  I060_056(w_060_056, w_031_476, w_046_250);
  and2 I060_057(w_060_057, w_001_845, w_001_620);
  not1 I060_058(w_060_058, w_052_1482);
  and2 I060_059(w_060_059, w_030_635, w_037_197);
  nand2 I060_060(w_060_060, w_039_1699, w_058_392);
  or2  I060_062(w_060_062, w_035_996, w_042_054);
  or2  I060_063(w_060_063, w_028_319, w_033_117);
  and2 I060_065(w_060_065, w_019_782, w_036_361);
  not1 I060_066(w_060_066, w_013_058);
  or2  I060_067(w_060_067, w_045_110, w_043_019);
  not1 I060_069(w_060_069, w_023_379);
  and2 I060_070(w_060_070, w_021_154, w_028_829);
  and2 I060_072(w_060_072, w_005_173, w_032_116);
  not1 I060_074(w_060_074, w_003_040);
  not1 I060_076(w_060_076, w_011_079);
  or2  I060_077(w_060_077, w_001_1127, w_002_235);
  nand2 I060_080(w_060_080, w_000_1686, w_037_496);
  not1 I060_081(w_060_081, w_000_1623);
  or2  I060_082(w_060_082, w_052_733, w_032_130);
  nand2 I060_084(w_060_084, w_026_772, w_038_457);
  or2  I060_088(w_060_088, w_037_119, w_002_301);
  or2  I060_091(w_060_091, w_040_856, w_057_592);
  and2 I060_093(w_060_093, w_013_096, w_010_217);
  or2  I060_094(w_060_094, w_040_978, w_031_674);
  nand2 I060_095(w_060_095, w_002_528, w_003_157);
  or2  I060_096(w_060_096, w_024_1188, w_021_075);
  not1 I060_097(w_060_097, w_018_280);
  not1 I060_098(w_060_098, w_015_073);
  not1 I060_100(w_060_100, w_000_1179);
  and2 I060_101(w_060_101, w_017_022, w_057_1166);
  not1 I060_102(w_060_102, w_015_243);
  and2 I060_103(w_060_103, w_034_595, w_048_560);
  or2  I060_104(w_060_104, w_034_494, w_029_987);
  and2 I060_106(w_060_106, w_002_120, w_045_266);
  or2  I061_000(w_061_000, w_013_226, w_010_171);
  and2 I061_009(w_061_009, w_048_276, w_017_251);
  nand2 I061_012(w_061_012, w_005_017, w_014_806);
  nand2 I061_049(w_061_049, w_024_017, w_034_322);
  nand2 I061_055(w_061_055, w_037_1711, w_023_785);
  or2  I061_071(w_061_071, w_043_101, w_049_1140);
  or2  I061_076(w_061_076, w_025_988, w_056_1424);
  or2  I061_084(w_061_084, w_013_173, w_043_022);
  not1 I061_089(w_061_089, w_026_048);
  and2 I061_106(w_061_106, w_015_026, w_018_159);
  or2  I061_108(w_061_108, w_016_008, w_006_021);
  not1 I061_114(w_061_114, w_007_107);
  not1 I061_121(w_061_121, w_020_525);
  or2  I061_151(w_061_151, w_003_068, w_005_379);
  and2 I061_161(w_061_161, w_039_938, w_044_697);
  not1 I061_182(w_061_182, w_059_207);
  nand2 I061_184(w_061_184, w_004_1767, w_013_060);
  or2  I061_201(w_061_201, w_036_1426, w_013_252);
  nand2 I061_212(w_061_212, w_030_126, w_000_272);
  not1 I061_213(w_061_213, w_017_1645);
  not1 I061_216(w_061_216, w_003_177);
  and2 I061_217(w_061_217, w_004_045, w_011_454);
  and2 I061_223(w_061_223, w_002_058, w_008_134);
  or2  I061_232(w_061_232, w_030_019, w_053_104);
  nand2 I061_236(w_061_236, w_046_181, w_043_099);
  or2  I061_240(w_061_240, w_032_086, w_007_213);
  or2  I061_255(w_061_255, w_020_857, w_009_013);
  or2  I061_260(w_061_260, w_039_977, w_049_112);
  and2 I061_263(w_061_263, w_009_030, w_053_105);
  nand2 I061_274(w_061_274, w_049_616, w_005_1381);
  and2 I061_279(w_061_279, w_041_140, w_051_023);
  or2  I061_280(w_061_280, w_058_891, w_020_183);
  or2  I061_293(w_061_293, w_036_1150, w_038_045);
  not1 I061_297(w_061_297, w_058_058);
  or2  I061_300(w_061_300, w_056_246, w_030_426);
  nand2 I061_303(w_061_303, w_027_065, w_047_653);
  nand2 I061_322(w_061_322, w_023_291, w_040_729);
  not1 I061_337(w_061_337, w_037_1488);
  or2  I061_363(w_061_363, w_013_044, w_038_362);
  or2  I061_367(w_061_367, w_031_611, w_006_153);
  or2  I061_373(w_061_373, w_014_273, w_047_384);
  not1 I061_374(w_061_374, w_030_766);
  nand2 I061_375(w_061_375, w_043_067, w_025_017);
  and2 I061_392(w_061_392, w_048_901, w_006_031);
  not1 I061_400(w_061_400, w_042_112);
  not1 I061_404(w_061_404, w_038_150);
  not1 I061_409(w_061_409, w_042_014);
  or2  I061_411(w_061_411, w_001_1123, w_053_118);
  and2 I061_424(w_061_424, w_049_999, w_028_119);
  not1 I061_426(w_061_426, w_035_1203);
  not1 I061_430(w_061_430, w_043_015);
  nand2 I061_435(w_061_435, w_038_451, w_058_1712);
  nand2 I061_437(w_061_437, w_006_196, w_051_581);
  nand2 I061_450(w_061_450, w_039_1643, w_038_136);
  not1 I061_461(w_061_461, w_021_089);
  or2  I061_468(w_061_468, w_032_173, w_055_750);
  or2  I061_473(w_061_473, w_035_1621, w_055_716);
  nand2 I061_479(w_061_479, w_017_491, w_029_541);
  and2 I061_486(w_061_486, w_031_226, w_022_420);
  nand2 I061_497(w_061_497, w_037_1194, w_037_175);
  and2 I061_506(w_061_506, w_042_008, w_022_195);
  not1 I061_513(w_061_513, w_044_1792);
  or2  I061_517(w_061_517, w_028_177, w_036_790);
  or2  I061_535(w_061_535, w_008_009, w_015_110);
  not1 I061_538(w_061_538, w_001_284);
  and2 I061_540(w_061_540, w_046_213, w_015_214);
  not1 I061_546(w_061_546, w_053_019);
  or2  I061_548(w_061_548, w_045_346, w_041_186);
  not1 I061_552(w_061_552, w_007_238);
  not1 I061_560(w_061_560, w_006_313);
  and2 I061_568(w_061_568, w_033_1375, w_043_098);
  and2 I061_582(w_061_582, w_047_028, w_009_076);
  and2 I061_585(w_061_585, w_053_095, w_018_223);
  or2  I061_607(w_061_607, w_028_130, w_056_251);
  or2  I061_622(w_061_622, w_058_080, w_058_875);
  nand2 I061_633(w_061_633, w_051_701, w_000_962);
  nand2 I061_643(w_061_643, w_009_018, w_005_984);
  and2 I061_644(w_061_644, w_019_648, w_010_310);
  not1 I061_663(w_061_663, w_048_677);
  not1 I062_015(w_062_015, w_022_099);
  and2 I062_027(w_062_027, w_006_256, w_047_231);
  and2 I062_032(w_062_032, w_000_1272, w_000_883);
  not1 I062_033(w_062_033, w_022_304);
  not1 I062_063(w_062_063, w_054_332);
  and2 I062_064(w_062_064, w_052_1844, w_003_156);
  not1 I062_071(w_062_071, w_058_1300);
  nand2 I062_072(w_062_072, w_037_355, w_007_1617);
  nand2 I062_077(w_062_077, w_011_406, w_045_1715);
  not1 I062_094(w_062_094, w_024_127);
  or2  I062_097(w_062_097, w_015_279, w_057_983);
  nand2 I062_105(w_062_105, w_004_1365, w_006_191);
  nand2 I062_106(w_062_106, w_035_349, w_019_331);
  not1 I062_127(w_062_127, w_049_309);
  and2 I062_137(w_062_137, w_004_920, w_000_397);
  nand2 I062_140(w_062_140, w_050_353, w_027_493);
  and2 I062_186(w_062_186, w_007_1292, w_054_508);
  or2  I062_196(w_062_196, w_030_112, w_047_606);
  nand2 I062_211(w_062_211, w_050_967, w_038_335);
  not1 I062_240(w_062_240, w_005_430);
  and2 I062_243(w_062_243, w_048_705, w_052_198);
  or2  I062_271(w_062_271, w_053_036, w_027_081);
  and2 I062_286(w_062_286, w_042_051, w_008_089);
  not1 I062_337(w_062_337, w_027_077);
  not1 I062_341(w_062_341, w_051_640);
  nand2 I062_349(w_062_349, w_008_745, w_042_027);
  nand2 I062_362(w_062_362, w_053_121, w_012_524);
  and2 I062_393(w_062_393, w_049_929, w_019_761);
  and2 I062_408(w_062_408, w_055_213, w_035_167);
  not1 I062_418(w_062_418, w_026_1365);
  nand2 I062_433(w_062_433, w_036_018, w_022_181);
  not1 I062_436(w_062_436, w_023_1218);
  and2 I062_447(w_062_447, w_046_233, w_006_134);
  or2  I062_465(w_062_465, w_035_467, w_032_013);
  or2  I062_497(w_062_497, w_049_055, w_033_1112);
  and2 I062_504(w_062_504, w_030_083, w_054_479);
  and2 I062_527(w_062_527, w_046_278, w_040_473);
  or2  I062_544(w_062_544, w_054_499, w_015_237);
  not1 I062_556(w_062_556, w_006_119);
  and2 I062_571(w_062_571, w_055_109, w_027_335);
  not1 I062_587(w_062_587, w_045_1830);
  or2  I062_605(w_062_605, w_050_718, w_012_353);
  or2  I062_608(w_062_608, w_049_260, w_061_373);
  and2 I062_618(w_062_618, w_042_029, w_018_220);
  nand2 I062_689(w_062_689, w_017_300, w_045_331);
  or2  I062_720(w_062_720, w_053_087, w_011_811);
  nand2 I062_732(w_062_732, w_043_022, w_030_055);
  nand2 I062_782(w_062_782, w_005_054, w_031_378);
  and2 I062_783(w_062_783, w_060_100, w_031_054);
  nand2 I062_787(w_062_787, w_024_471, w_016_007);
  or2  I062_805(w_062_805, w_047_056, w_051_958);
  not1 I062_817(w_062_817, w_007_1600);
  nand2 I062_876(w_062_876, w_024_778, w_009_096);
  or2  I062_878(w_062_878, w_046_045, w_032_035);
  or2  I062_887(w_062_887, w_039_1227, w_025_491);
  nand2 I062_900(w_062_900, w_061_089, w_042_031);
  or2  I062_962(w_062_962, w_013_212, w_033_1376);
  or2  I062_972(w_062_972, w_033_1634, w_019_732);
  and2 I062_973(w_062_973, w_006_083, w_051_675);
  not1 I062_998(w_062_998, w_007_247);
  and2 I062_1003(w_062_1003, w_053_029, w_054_399);
  or2  I062_1016(w_062_1016, w_035_028, w_056_830);
  or2  I062_1111(w_062_1111, w_028_267, w_017_798);
  or2  I062_1124(w_062_1124, w_017_003, w_032_160);
  and2 I062_1158(w_062_1158, w_003_173, w_005_115);
  not1 I062_1177(w_062_1177, w_056_659);
  nand2 I062_1180(w_062_1180, w_055_466, w_006_342);
  nand2 I062_1181(w_062_1181, w_060_024, w_004_076);
  not1 I062_1222(w_062_1222, w_022_403);
  not1 I062_1289(w_062_1289, w_002_538);
  nand2 I062_1292(w_062_1292, w_050_1023, w_059_381);
  and2 I062_1296(w_062_1296, w_041_124, w_052_1364);
  nand2 I062_1307(w_062_1307, w_059_478, w_056_125);
  not1 I062_1332(w_062_1332, w_023_1219);
  or2  I063_006(w_063_006, w_021_074, w_034_226);
  and2 I063_016(w_063_016, w_016_033, w_042_027);
  and2 I063_019(w_063_019, w_001_169, w_048_629);
  and2 I063_027(w_063_027, w_004_538, w_039_018);
  nand2 I063_038(w_063_038, w_055_715, w_051_1064);
  and2 I063_041(w_063_041, w_000_903, w_018_225);
  or2  I063_043(w_063_043, w_051_292, w_052_242);
  nand2 I063_049(w_063_049, w_016_034, w_049_651);
  not1 I063_054(w_063_054, w_041_157);
  or2  I063_055(w_063_055, w_000_1598, w_012_607);
  not1 I063_059(w_063_059, w_006_081);
  not1 I063_060(w_063_060, w_059_608);
  or2  I063_093(w_063_093, w_010_058, w_035_1464);
  or2  I063_095(w_063_095, w_014_107, w_057_1410);
  and2 I063_129(w_063_129, w_031_078, w_005_1538);
  not1 I063_137(w_063_137, w_032_119);
  nand2 I063_140(w_063_140, w_013_318, w_039_1392);
  or2  I063_145(w_063_145, w_013_264, w_020_664);
  and2 I063_171(w_063_171, w_050_1244, w_020_989);
  or2  I063_175(w_063_175, w_016_031, w_017_1195);
  not1 I063_183(w_063_183, w_061_400);
  not1 I063_184(w_063_184, w_024_182);
  not1 I063_194(w_063_194, w_035_077);
  and2 I063_255(w_063_255, w_060_039, w_017_335);
  nand2 I063_264(w_063_264, w_030_732, w_029_1276);
  and2 I063_270(w_063_270, w_057_222, w_023_1114);
  or2  I063_283(w_063_283, w_019_1029, w_054_057);
  and2 I063_287(w_063_287, w_042_135, w_001_137);
  and2 I063_289(w_063_289, w_057_743, w_041_206);
  not1 I063_292(w_063_292, w_062_787);
  and2 I063_295(w_063_295, w_033_222, w_041_008);
  and2 I063_312(w_063_312, w_056_231, w_043_040);
  not1 I063_345(w_063_345, w_013_261);
  or2  I063_358(w_063_358, w_051_703, w_031_645);
  or2  I063_373(w_063_373, w_025_150, w_051_1022);
  nand2 I063_375(w_063_375, w_027_414, w_041_250);
  and2 I063_388(w_063_388, w_021_212, w_034_011);
  nand2 I063_392(w_063_392, w_056_211, w_041_152);
  nand2 I063_407(w_063_407, w_036_1440, w_020_557);
  not1 I063_422(w_063_422, w_054_532);
  and2 I063_566(w_063_566, w_033_987, w_003_237);
  or2  I063_572(w_063_572, w_055_154, w_006_127);
  not1 I063_590(w_063_590, w_055_167);
  or2  I063_597(w_063_597, w_004_1062, w_060_010);
  nand2 I063_600(w_063_600, w_031_341, w_051_209);
  nand2 I063_613(w_063_613, w_015_033, w_021_023);
  nand2 I063_618(w_063_618, w_039_429, w_054_606);
  or2  I063_619(w_063_619, w_021_007, w_013_054);
  and2 I063_629(w_063_629, w_060_018, w_038_401);
  and2 I063_695(w_063_695, w_038_136, w_002_552);
  nand2 I063_706(w_063_706, w_039_932, w_028_763);
  and2 I063_722(w_063_722, w_026_984, w_061_114);
  and2 I063_725(w_063_725, w_019_305, w_032_012);
  not1 I063_749(w_063_749, w_005_1588);
  nand2 I063_837(w_063_837, w_021_071, w_045_072);
  or2  I063_909(w_063_909, w_048_567, w_035_209);
  or2  I063_966(w_063_966, w_008_186, w_053_064);
  or2  I063_975(w_063_975, w_052_904, w_017_602);
  or2  I063_1029(w_063_1029, w_019_1026, w_031_925);
  nand2 I063_1040(w_063_1040, w_002_214, w_015_249);
  and2 I063_1059(w_063_1059, w_055_475, w_014_713);
  nand2 I063_1088(w_063_1088, w_060_094, w_005_1222);
  nand2 I063_1094(w_063_1094, w_021_128, w_022_206);
  not1 I063_1100(w_063_1100, w_054_577);
  and2 I063_1122(w_063_1122, w_017_150, w_028_280);
  and2 I063_1140(w_063_1140, w_044_1550, w_036_173);
  nand2 I063_1149(w_063_1149, w_011_260, w_013_281);
  and2 I063_1157(w_063_1157, w_022_064, w_041_084);
  not1 I063_1164(w_063_1164, w_001_1301);
  not1 I063_1171(w_063_1171, w_002_125);
  nand2 I063_1173(w_063_1173, w_001_236, w_053_118);
  not1 I063_1247(w_063_1247, w_050_406);
  nand2 I063_1251(w_063_1251, w_037_046, w_015_048);
  not1 I063_1265(w_063_1265, w_060_012);
  and2 I063_1294(w_063_1294, w_009_028, w_048_159);
  nand2 I063_1297(w_063_1297, w_040_489, w_062_196);
  or2  I063_1311(w_063_1311, w_012_083, w_010_275);
  and2 I063_1336(w_063_1336, w_034_471, w_049_530);
  and2 I063_1337(w_063_1337, w_038_208, w_045_1328);
  and2 I063_1375(w_063_1375, w_055_164, w_028_814);
  nand2 I063_1411(w_063_1411, w_026_396, w_025_825);
  nand2 I063_1422(w_063_1422, w_056_165, w_013_296);
  and2 I063_1429(w_063_1429, w_022_376, w_042_003);
  nand2 I063_1486(w_063_1486, w_039_788, w_016_024);
  or2  I063_1492(w_063_1492, w_007_368, w_011_501);
  not1 I063_1500(w_063_1500, w_032_237);
  nand2 I063_1501(w_063_1501, w_034_404, w_006_148);
  and2 I063_1561(w_063_1561, w_007_074, w_035_228);
  nand2 I063_1578(w_063_1578, w_010_178, w_011_758);
  nand2 I063_1583(w_063_1583, w_059_651, w_022_231);
  and2 I063_1594(w_063_1594, w_004_366, w_003_045);
  nand2 I063_1604(w_063_1604, w_043_081, w_036_222);
  or2  I064_036(w_064_036, w_021_041, w_043_041);
  nand2 I064_039(w_064_039, w_035_003, w_031_485);
  not1 I064_085(w_064_085, w_047_022);
  or2  I064_096(w_064_096, w_053_016, w_063_1311);
  not1 I064_102(w_064_102, w_056_411);
  and2 I064_108(w_064_108, w_034_569, w_008_018);
  not1 I064_115(w_064_115, w_043_013);
  and2 I064_140(w_064_140, w_058_125, w_022_107);
  not1 I064_141(w_064_141, w_036_283);
  or2  I064_145(w_064_145, w_024_949, w_063_049);
  nand2 I064_147(w_064_147, w_014_819, w_013_254);
  not1 I064_156(w_064_156, w_032_045);
  nand2 I064_159(w_064_159, w_020_1255, w_039_250);
  and2 I064_170(w_064_170, w_058_415, w_052_1038);
  or2  I064_179(w_064_179, w_051_773, w_009_041);
  and2 I064_190(w_064_190, w_001_147, w_035_1098);
  or2  I064_193(w_064_193, w_046_232, w_008_242);
  and2 I064_197(w_064_197, w_044_134, w_004_1590);
  or2  I064_210(w_064_210, w_006_230, w_035_037);
  or2  I064_227(w_064_227, w_024_1424, w_054_007);
  nand2 I064_234(w_064_234, w_034_006, w_031_136);
  or2  I064_239(w_064_239, w_013_250, w_007_164);
  and2 I064_252(w_064_252, w_053_047, w_000_1131);
  nand2 I064_254(w_064_254, w_033_457, w_051_1012);
  not1 I064_264(w_064_264, w_051_290);
  or2  I064_266(w_064_266, w_041_121, w_020_416);
  nand2 I064_293(w_064_293, w_010_126, w_051_891);
  nand2 I064_305(w_064_305, w_028_871, w_047_149);
  not1 I064_330(w_064_330, w_013_312);
  or2  I064_364(w_064_364, w_013_016, w_055_242);
  or2  I064_380(w_064_380, w_026_450, w_015_014);
  nand2 I064_396(w_064_396, w_038_485, w_004_1152);
  or2  I064_405(w_064_405, w_062_337, w_010_372);
  nand2 I064_455(w_064_455, w_039_1856, w_030_382);
  not1 I064_474(w_064_474, w_028_062);
  and2 I064_479(w_064_479, w_007_1334, w_056_1511);
  and2 I064_492(w_064_492, w_021_182, w_058_822);
  nand2 I064_563(w_064_563, w_055_007, w_059_303);
  nand2 I064_586(w_064_586, w_030_239, w_058_074);
  nand2 I064_607(w_064_607, w_018_047, w_058_1086);
  or2  I064_609(w_064_609, w_062_349, w_013_156);
  nand2 I064_631(w_064_631, w_054_440, w_000_822);
  and2 I064_636(w_064_636, w_025_082, w_023_1298);
  and2 I064_639(w_064_639, w_034_079, w_043_056);
  not1 I064_666(w_064_666, w_043_092);
  and2 I064_677(w_064_677, w_039_612, w_035_096);
  not1 I064_728(w_064_728, w_063_295);
  or2  I064_749(w_064_749, w_003_143, w_005_1005);
  or2  I064_772(w_064_772, w_023_1115, w_060_038);
  not1 I064_775(w_064_775, w_007_567);
  nand2 I064_790(w_064_790, w_034_498, w_011_170);
  not1 I064_795(w_064_795, w_011_386);
  not1 I064_805(w_064_805, w_063_095);
  nand2 I064_829(w_064_829, w_055_469, w_004_1593);
  nand2 I064_861(w_064_861, w_000_197, w_033_341);
  not1 I064_884(w_064_884, w_012_096);
  or2  I064_889(w_064_889, w_050_686, w_019_771);
  nand2 I064_891(w_064_891, w_057_1252, w_015_039);
  not1 I064_904(w_064_904, w_024_208);
  nand2 I064_912(w_064_912, w_027_150, w_041_267);
  not1 I064_926(w_064_926, w_055_149);
  not1 I064_941(w_064_941, w_052_1375);
  and2 I064_954(w_064_954, w_058_1485, w_031_366);
  and2 I064_996(w_064_996, w_056_512, w_020_1072);
  nand2 I064_999(w_064_999, w_060_101, w_049_031);
  nand2 I064_1012(w_064_1012, w_031_395, w_024_087);
  nand2 I064_1046(w_064_1046, w_048_583, w_060_104);
  not1 I064_1047(w_064_1047, w_025_842);
  nand2 I064_1058(w_064_1058, w_024_812, w_022_370);
  or2  I064_1064(w_064_1064, w_022_410, w_048_751);
  and2 I064_1081(w_064_1081, w_048_117, w_056_519);
  and2 I064_1094(w_064_1094, w_012_175, w_022_171);
  or2  I064_1135(w_064_1135, w_045_288, w_006_244);
  not1 I064_1137(w_064_1137, w_063_1429);
  not1 I064_1140(w_064_1140, w_033_1324);
  nand2 I064_1150(w_064_1150, w_014_015, w_022_023);
  not1 I064_1154(w_064_1154, w_058_1064);
  not1 I064_1161(w_064_1161, w_053_109);
  and2 I064_1186(w_064_1186, w_036_272, w_010_206);
  nand2 I064_1204(w_064_1204, w_017_1888, w_001_687);
  nand2 I064_1225(w_064_1225, w_012_627, w_057_1467);
  not1 I064_1238(w_064_1238, w_052_1295);
  or2  I064_1283(w_064_1283, w_015_172, w_015_038);
  and2 I064_1303(w_064_1303, w_002_188, w_045_1653);
  and2 I064_1323(w_064_1323, w_018_004, w_045_802);
  not1 I064_1337(w_064_1337, w_020_667);
  or2  I064_1362(w_064_1362, w_051_1044, w_041_042);
  and2 I064_1374(w_064_1374, w_037_1259, w_005_160);
  not1 I064_1377(w_064_1377, w_019_405);
  not1 I064_1392(w_064_1392, w_000_1523);
  not1 I064_1433(w_064_1433, w_004_060);
  and2 I064_1435(w_064_1435, w_060_026, w_048_783);
  or2  I064_1438(w_064_1438, w_052_1104, w_037_879);
  and2 I064_1440(w_064_1440, w_024_1622, w_030_078);
  or2  I064_1456(w_064_1456, w_049_013, w_044_1426);
  nand2 I064_1466(w_064_1466, w_062_211, w_001_016);
  nand2 I064_1474(w_064_1474, w_012_655, w_004_897);
  nand2 I064_1509(w_064_1509, w_001_1262, w_025_548);
  or2  I064_1513(w_064_1513, w_033_175, w_013_078);
  or2  I064_1583(w_064_1583, w_058_1779, w_030_570);
  nand2 I064_1594(w_064_1594, w_024_844, w_013_122);
  not1 I064_1602(w_064_1602, w_058_1144);
  or2  I064_1643(w_064_1643, w_035_130, w_018_043);
  or2  I064_1658(w_064_1658, w_061_071, w_034_500);
  not1 I065_000(w_065_000, w_022_312);
  nand2 I065_001(w_065_001, w_006_243, w_043_070);
  or2  I065_002(w_065_002, w_037_629, w_020_289);
  not1 I065_003(w_065_003, w_055_339);
  and2 I065_004(w_065_004, w_010_328, w_050_370);
  not1 I065_005(w_065_005, w_025_137);
  not1 I066_007(w_066_007, w_062_1158);
  nand2 I066_009(w_066_009, w_043_077, w_041_077);
  or2  I066_013(w_066_013, w_008_021, w_054_477);
  or2  I066_016(w_066_016, w_000_1926, w_008_228);
  nand2 I066_022(w_066_022, w_029_283, w_063_283);
  not1 I066_043(w_066_043, w_022_391);
  nand2 I066_047(w_066_047, w_063_572, w_047_501);
  nand2 I066_063(w_066_063, w_055_327, w_031_814);
  or2  I066_066(w_066_066, w_062_127, w_063_749);
  or2  I066_069(w_066_069, w_012_596, w_030_753);
  or2  I066_075(w_066_075, w_006_010, w_044_1146);
  nand2 I066_077(w_066_077, w_003_027, w_047_441);
  not1 I066_086(w_066_086, w_012_058);
  and2 I066_090(w_066_090, w_043_062, w_051_1064);
  and2 I066_116(w_066_116, w_036_1129, w_061_622);
  not1 I066_142(w_066_142, w_003_075);
  not1 I066_154(w_066_154, w_027_460);
  or2  I066_156(w_066_156, w_012_590, w_065_000);
  and2 I066_162(w_066_162, w_045_490, w_051_580);
  not1 I066_188(w_066_188, w_056_1540);
  nand2 I066_213(w_066_213, w_049_1207, w_053_017);
  nand2 I066_222(w_066_222, w_023_459, w_043_030);
  and2 I066_223(w_066_223, w_020_377, w_026_394);
  nand2 I066_282(w_066_282, w_007_232, w_042_096);
  or2  I066_291(w_066_291, w_022_409, w_028_001);
  nand2 I066_307(w_066_307, w_001_1237, w_014_629);
  nand2 I066_324(w_066_324, w_024_1377, w_037_352);
  or2  I066_327(w_066_327, w_020_915, w_023_1199);
  nand2 I066_332(w_066_332, w_035_637, w_042_014);
  not1 I066_355(w_066_355, w_013_223);
  not1 I066_363(w_066_363, w_022_051);
  or2  I066_373(w_066_373, w_062_973, w_055_260);
  not1 I066_378(w_066_378, w_020_1219);
  or2  I066_380(w_066_380, w_037_1432, w_024_1235);
  not1 I066_404(w_066_404, w_011_790);
  and2 I066_412(w_066_412, w_014_058, w_065_000);
  or2  I066_430(w_066_430, w_039_1362, w_052_1709);
  not1 I066_522(w_066_522, w_037_190);
  and2 I066_537(w_066_537, w_044_931, w_055_421);
  nand2 I066_546(w_066_546, w_041_115, w_010_092);
  nand2 I066_558(w_066_558, w_002_425, w_043_089);
  or2  I066_562(w_066_562, w_017_1911, w_060_081);
  and2 I066_574(w_066_574, w_000_573, w_012_165);
  or2  I066_602(w_066_602, w_014_651, w_009_075);
  not1 I066_640(w_066_640, w_041_128);
  not1 I066_702(w_066_702, w_051_268);
  and2 I066_714(w_066_714, w_050_1020, w_016_018);
  nand2 I066_722(w_066_722, w_057_209, w_043_014);
  or2  I066_731(w_066_731, w_045_1333, w_030_273);
  or2  I066_738(w_066_738, w_043_041, w_003_285);
  nand2 I066_753(w_066_753, w_018_149, w_010_333);
  nand2 I066_767(w_066_767, w_030_636, w_033_1032);
  not1 I066_798(w_066_798, w_036_166);
  nand2 I066_823(w_066_823, w_045_1064, w_029_622);
  or2  I066_845(w_066_845, w_019_030, w_056_1315);
  nand2 I066_859(w_066_859, w_037_563, w_028_731);
  nand2 I066_863(w_066_863, w_022_172, w_016_010);
  nand2 I066_870(w_066_870, w_058_1121, w_044_1139);
  or2  I066_889(w_066_889, w_021_009, w_046_075);
  nand2 I066_896(w_066_896, w_049_634, w_049_1057);
  or2  I066_898(w_066_898, w_002_245, w_024_031);
  nand2 I066_900(w_066_900, w_062_465, w_027_334);
  or2  I066_909(w_066_909, w_015_136, w_037_1035);
  and2 I066_930(w_066_930, w_061_479, w_041_150);
  nand2 I066_971(w_066_971, w_004_1039, w_033_055);
  or2  I066_989(w_066_989, w_026_262, w_004_1001);
  not1 I066_1009(w_066_1009, w_000_314);
  not1 I066_1027(w_066_1027, w_046_018);
  or2  I066_1040(w_066_1040, w_009_067, w_024_509);
  not1 I066_1093(w_066_1093, w_042_073);
  not1 I066_1151(w_066_1151, w_051_292);
  and2 I067_017(w_067_017, w_028_247, w_019_1037);
  and2 I067_019(w_067_019, w_047_103, w_028_236);
  not1 I067_048(w_067_048, w_035_240);
  and2 I067_080(w_067_080, w_053_121, w_036_1309);
  and2 I067_105(w_067_105, w_040_148, w_063_629);
  and2 I067_160(w_067_160, w_029_1141, w_008_110);
  or2  I067_179(w_067_179, w_001_864, w_017_935);
  and2 I067_183(w_067_183, w_037_156, w_049_494);
  not1 I067_185(w_067_185, w_002_473);
  not1 I067_200(w_067_200, w_040_380);
  or2  I067_206(w_067_206, w_054_482, w_048_966);
  not1 I067_209(w_067_209, w_052_059);
  and2 I067_225(w_067_225, w_001_130, w_024_924);
  and2 I067_237(w_067_237, w_000_726, w_039_1362);
  and2 I067_258(w_067_258, w_028_181, w_034_134);
  or2  I067_267(w_067_267, w_048_018, w_028_191);
  or2  I067_280(w_067_280, w_031_330, w_046_145);
  nand2 I067_287(w_067_287, w_052_218, w_063_1122);
  nand2 I067_288(w_067_288, w_053_048, w_018_070);
  not1 I067_292(w_067_292, w_005_801);
  nand2 I067_338(w_067_338, w_040_315, w_010_279);
  or2  I067_360(w_067_360, w_038_299, w_055_076);
  not1 I067_376(w_067_376, w_054_102);
  nand2 I067_403(w_067_403, w_036_1237, w_058_768);
  or2  I067_418(w_067_418, w_040_056, w_039_650);
  and2 I067_434(w_067_434, w_046_207, w_033_1295);
  and2 I067_462(w_067_462, w_046_140, w_044_1141);
  nand2 I067_477(w_067_477, w_013_013, w_044_465);
  and2 I067_512(w_067_512, w_003_021, w_053_068);
  nand2 I067_531(w_067_531, w_012_249, w_025_1097);
  nand2 I067_532(w_067_532, w_005_338, w_052_987);
  or2  I067_541(w_067_541, w_050_174, w_000_1729);
  not1 I067_544(w_067_544, w_047_543);
  not1 I067_558(w_067_558, w_034_403);
  not1 I067_582(w_067_582, w_054_170);
  or2  I067_589(w_067_589, w_053_040, w_022_310);
  not1 I067_595(w_067_595, w_002_135);
  not1 I067_603(w_067_603, w_049_220);
  and2 I067_609(w_067_609, w_016_010, w_024_686);
  not1 I067_620(w_067_620, w_017_236);
  not1 I067_639(w_067_639, w_056_161);
  and2 I067_651(w_067_651, w_056_810, w_014_085);
  or2  I067_655(w_067_655, w_014_090, w_028_340);
  and2 I067_665(w_067_665, w_047_391, w_049_347);
  nand2 I067_676(w_067_676, w_051_595, w_042_141);
  not1 I067_682(w_067_682, w_049_345);
  not1 I067_688(w_067_688, w_046_128);
  and2 I067_690(w_067_690, w_019_080, w_037_1083);
  and2 I067_692(w_067_692, w_055_284, w_044_1224);
  nand2 I067_696(w_067_696, w_062_286, w_022_070);
  not1 I067_703(w_067_703, w_013_328);
  not1 I067_727(w_067_727, w_032_227);
  or2  I067_742(w_067_742, w_011_120, w_004_566);
  or2  I067_746(w_067_746, w_034_568, w_052_1072);
  or2  I067_758(w_067_758, w_047_550, w_020_591);
  and2 I067_763(w_067_763, w_061_106, w_000_071);
  nand2 I067_786(w_067_786, w_038_002, w_061_585);
  and2 I067_799(w_067_799, w_033_697, w_035_1431);
  nand2 I067_807(w_067_807, w_041_044, w_021_277);
  or2  I067_871(w_067_871, w_046_012, w_037_705);
  or2  I067_872(w_067_872, w_023_1595, w_028_204);
  and2 I067_896(w_067_896, w_022_085, w_016_013);
  or2  I067_898(w_067_898, w_005_759, w_040_700);
  and2 I067_905(w_067_905, w_037_690, w_002_564);
  and2 I067_912(w_067_912, w_007_014, w_047_340);
  not1 I067_943(w_067_943, w_028_056);
  nand2 I067_961(w_067_961, w_061_300, w_053_098);
  and2 I067_962(w_067_962, w_022_011, w_058_064);
  nand2 I067_965(w_067_965, w_060_093, w_015_150);
  and2 I068_000(w_068_000, w_021_225, w_050_368);
  not1 I068_003(w_068_003, w_066_043);
  and2 I068_011(w_068_011, w_013_029, w_003_195);
  not1 I068_013(w_068_013, w_027_393);
  and2 I068_017(w_068_017, w_009_026, w_007_1160);
  not1 I068_018(w_068_018, w_028_633);
  or2  I068_019(w_068_019, w_039_533, w_013_249);
  nand2 I068_021(w_068_021, w_003_215, w_067_267);
  or2  I068_022(w_068_022, w_001_014, w_042_077);
  or2  I068_026(w_068_026, w_027_249, w_022_277);
  and2 I068_027(w_068_027, w_047_341, w_063_1094);
  and2 I068_029(w_068_029, w_003_059, w_014_252);
  nand2 I068_030(w_068_030, w_063_055, w_055_389);
  nand2 I068_031(w_068_031, w_067_360, w_008_763);
  or2  I068_036(w_068_036, w_003_079, w_012_366);
  and2 I068_037(w_068_037, w_008_444, w_031_619);
  and2 I068_038(w_068_038, w_039_1731, w_004_245);
  and2 I068_041(w_068_041, w_019_877, w_055_717);
  and2 I068_048(w_068_048, w_001_225, w_024_1121);
  nand2 I068_050(w_068_050, w_006_075, w_052_587);
  or2  I068_055(w_068_055, w_058_531, w_008_010);
  or2  I068_059(w_068_059, w_015_001, w_044_112);
  or2  I068_062(w_068_062, w_026_1347, w_042_029);
  and2 I068_073(w_068_073, w_038_150, w_067_651);
  nand2 I068_075(w_068_075, w_056_637, w_017_1563);
  not1 I068_078(w_068_078, w_017_713);
  not1 I068_083(w_068_083, w_059_042);
  nand2 I068_085(w_068_085, w_029_178, w_032_182);
  nand2 I068_086(w_068_086, w_043_092, w_053_043);
  nand2 I068_095(w_068_095, w_067_183, w_021_092);
  not1 I068_097(w_068_097, w_003_111);
  nand2 I068_105(w_068_105, w_038_207, w_009_025);
  not1 I068_106(w_068_106, w_003_219);
  not1 I068_110(w_068_110, w_009_065);
  or2  I068_114(w_068_114, w_005_1258, w_031_357);
  nand2 I068_119(w_068_119, w_045_1071, w_045_1538);
  and2 I068_126(w_068_126, w_029_092, w_009_105);
  nand2 I068_135(w_068_135, w_044_1465, w_067_688);
  not1 I068_140(w_068_140, w_062_243);
  and2 I068_141(w_068_141, w_016_022, w_031_988);
  not1 I068_142(w_068_142, w_020_503);
  or2  I068_151(w_068_151, w_050_1499, w_008_402);
  not1 I068_157(w_068_157, w_039_310);
  and2 I068_160(w_068_160, w_040_979, w_027_297);
  or2  I068_163(w_068_163, w_002_048, w_035_1147);
  not1 I068_164(w_068_164, w_063_1486);
  or2  I068_165(w_068_165, w_014_140, w_028_035);
  or2  I068_166(w_068_166, w_042_027, w_003_140);
  nand2 I068_169(w_068_169, w_029_083, w_019_277);
  or2  I068_171(w_068_171, w_056_1109, w_061_213);
  and2 I068_176(w_068_176, w_000_1220, w_063_619);
  not1 I068_179(w_068_179, w_066_327);
  not1 I068_184(w_068_184, w_005_742);
  not1 I068_189(w_068_189, w_006_137);
  not1 I068_190(w_068_190, w_064_1374);
  nand2 I068_194(w_068_194, w_003_315, w_016_000);
  or2  I068_197(w_068_197, w_006_153, w_018_186);
  or2  I068_200(w_068_200, w_034_570, w_027_366);
  nand2 I068_203(w_068_203, w_017_732, w_028_851);
  nand2 I068_209(w_068_209, w_054_572, w_002_089);
  and2 I068_210(w_068_210, w_030_170, w_037_1656);
  nand2 I068_211(w_068_211, w_035_276, w_015_283);
  or2  I068_216(w_068_216, w_024_939, w_005_490);
  or2  I068_223(w_068_223, w_039_847, w_025_221);
  and2 I068_224(w_068_224, w_019_358, w_011_557);
  nand2 I068_233(w_068_233, w_020_941, w_028_112);
  nand2 I068_234(w_068_234, w_036_1220, w_017_1113);
  and2 I068_236(w_068_236, w_035_941, w_046_195);
  or2  I068_239(w_068_239, w_042_074, w_056_1562);
  nand2 I068_240(w_068_240, w_016_037, w_006_189);
  not1 I068_243(w_068_243, w_066_022);
  and2 I069_001(w_069_001, w_068_038, w_042_035);
  nand2 I069_019(w_069_019, w_043_013, w_035_095);
  or2  I069_021(w_069_021, w_048_135, w_002_417);
  nand2 I069_038(w_069_038, w_045_041, w_025_1134);
  or2  I069_039(w_069_039, w_043_092, w_013_015);
  not1 I069_049(w_069_049, w_023_126);
  not1 I069_053(w_069_053, w_068_236);
  nand2 I069_068(w_069_068, w_061_411, w_002_230);
  nand2 I069_072(w_069_072, w_029_053, w_029_934);
  or2  I069_182(w_069_182, w_011_455, w_005_484);
  and2 I069_188(w_069_188, w_043_043, w_029_1210);
  nand2 I069_283(w_069_283, w_067_965, w_044_665);
  or2  I069_312(w_069_312, w_027_476, w_032_019);
  nand2 I069_331(w_069_331, w_010_114, w_006_333);
  and2 I069_350(w_069_350, w_005_287, w_019_485);
  or2  I069_368(w_069_368, w_033_033, w_056_668);
  nand2 I069_436(w_069_436, w_022_059, w_033_139);
  not1 I069_474(w_069_474, w_041_052);
  not1 I069_479(w_069_479, w_057_1838);
  and2 I069_510(w_069_510, w_002_001, w_022_230);
  nand2 I069_568(w_069_568, w_040_086, w_013_179);
  and2 I069_620(w_069_620, w_047_568, w_046_124);
  and2 I069_681(w_069_681, w_021_102, w_064_1323);
  and2 I069_723(w_069_723, w_048_132, w_047_230);
  and2 I069_760(w_069_760, w_049_1221, w_007_024);
  or2  I069_805(w_069_805, w_000_608, w_012_183);
  and2 I069_828(w_069_828, w_025_848, w_028_798);
  or2  I069_866(w_069_866, w_022_123, w_061_560);
  and2 I069_920(w_069_920, w_018_220, w_027_105);
  nand2 I069_921(w_069_921, w_031_511, w_044_613);
  nand2 I069_970(w_069_970, w_046_056, w_050_275);
  nand2 I069_976(w_069_976, w_015_075, w_013_268);
  or2  I069_980(w_069_980, w_051_828, w_025_1258);
  and2 I069_1167(w_069_1167, w_048_713, w_017_023);
  not1 I069_1270(w_069_1270, w_014_053);
  or2  I069_1276(w_069_1276, w_008_244, w_068_165);
  nand2 I069_1285(w_069_1285, w_052_965, w_045_1414);
  and2 I069_1356(w_069_1356, w_045_1693, w_026_068);
  nand2 I069_1365(w_069_1365, w_034_133, w_068_216);
  nand2 I069_1369(w_069_1369, w_030_042, w_044_129);
  not1 I069_1571(w_069_1571, w_019_569);
  nand2 I069_1600(w_069_1600, w_036_577, w_017_198);
  nand2 I069_1618(w_069_1618, w_023_157, w_040_075);
  nand2 I069_1620(w_069_1620, w_018_269, w_014_082);
  or2  I069_1642(w_069_1642, w_045_599, w_058_302);
  and2 I069_1675(w_069_1675, w_004_1329, w_022_305);
  nand2 I069_1681(w_069_1681, w_024_107, w_054_618);
  not1 I069_1723(w_069_1723, w_065_002);
  and2 I069_1729(w_069_1729, w_000_948, w_005_1605);
  and2 I069_1731(w_069_1731, w_054_581, w_022_163);
  not1 I069_1744(w_069_1744, w_032_075);
  not1 I069_1762(w_069_1762, w_027_229);
  and2 I069_1776(w_069_1776, w_027_398, w_067_943);
  nand2 I069_1807(w_069_1807, w_012_336, w_034_214);
  and2 I069_1818(w_069_1818, w_020_777, w_041_111);
  or2  I070_004(w_070_004, w_019_926, w_028_285);
  nand2 I070_005(w_070_005, w_064_492, w_025_259);
  and2 I070_013(w_070_013, w_036_107, w_042_022);
  not1 I070_014(w_070_014, w_014_509);
  nand2 I070_015(w_070_015, w_027_579, w_016_027);
  not1 I070_022(w_070_022, w_015_280);
  or2  I070_031(w_070_031, w_010_256, w_065_001);
  or2  I070_032(w_070_032, w_047_594, w_016_016);
  not1 I070_034(w_070_034, w_051_996);
  not1 I070_035(w_070_035, w_068_163);
  nand2 I070_045(w_070_045, w_055_311, w_043_026);
  or2  I070_050(w_070_050, w_048_090, w_052_338);
  not1 I070_051(w_070_051, w_023_1313);
  not1 I070_056(w_070_056, w_055_835);
  or2  I070_061(w_070_061, w_045_1756, w_030_783);
  nand2 I070_062(w_070_062, w_045_066, w_019_791);
  not1 I070_077(w_070_077, w_004_016);
  and2 I070_079(w_070_079, w_021_005, w_015_160);
  or2  I070_080(w_070_080, w_018_224, w_037_007);
  or2  I070_093(w_070_093, w_018_069, w_034_578);
  nand2 I070_107(w_070_107, w_055_160, w_006_319);
  nand2 I070_110(w_070_110, w_038_382, w_004_548);
  not1 I070_114(w_070_114, w_052_266);
  and2 I070_120(w_070_120, w_063_145, w_042_121);
  or2  I070_146(w_070_146, w_026_203, w_015_012);
  not1 I070_149(w_070_149, w_019_262);
  not1 I070_150(w_070_150, w_005_1025);
  and2 I070_160(w_070_160, w_017_851, w_037_793);
  nand2 I070_172(w_070_172, w_042_094, w_048_409);
  or2  I070_175(w_070_175, w_022_036, w_032_081);
  or2  I070_177(w_070_177, w_066_142, w_008_674);
  and2 I070_180(w_070_180, w_025_337, w_022_149);
  and2 I070_182(w_070_182, w_012_537, w_062_1181);
  nand2 I070_183(w_070_183, w_021_205, w_001_1571);
  and2 I070_204(w_070_204, w_067_179, w_059_653);
  or2  I070_212(w_070_212, w_032_031, w_048_148);
  and2 I070_213(w_070_213, w_016_015, w_003_142);
  and2 I070_231(w_070_231, w_068_003, w_007_1334);
  and2 I070_244(w_070_244, w_064_405, w_005_1050);
  nand2 I070_250(w_070_250, w_026_345, w_042_104);
  not1 I070_260(w_070_260, w_052_1566);
  not1 I070_270(w_070_270, w_068_031);
  and2 I070_285(w_070_285, w_022_268, w_051_285);
  and2 I070_314(w_070_314, w_007_311, w_044_1752);
  nand2 I070_318(w_070_318, w_065_000, w_028_454);
  nand2 I070_369(w_070_369, w_028_111, w_031_274);
  nand2 I070_371(w_070_371, w_023_939, w_063_264);
  nand2 I070_374(w_070_374, w_039_526, w_046_034);
  nand2 I070_376(w_070_376, w_050_1158, w_051_849);
  nand2 I070_379(w_070_379, w_041_237, w_042_034);
  not1 I070_387(w_070_387, w_057_790);
  and2 I070_391(w_070_391, w_009_105, w_052_1289);
  nand2 I070_401(w_070_401, w_023_491, w_046_140);
  or2  I070_405(w_070_405, w_050_683, w_032_105);
  or2  I070_409(w_070_409, w_043_022, w_045_1646);
  nand2 I070_423(w_070_423, w_024_781, w_036_1306);
  not1 I070_427(w_070_427, w_056_835);
  not1 I070_430(w_070_430, w_007_1493);
  or2  I070_432(w_070_432, w_042_135, w_065_003);
  not1 I070_446(w_070_446, w_017_703);
  and2 I070_448(w_070_448, w_025_1251, w_034_653);
  and2 I070_450(w_070_450, w_027_387, w_020_478);
  or2  I070_455(w_070_455, w_021_060, w_055_671);
  nand2 I070_459(w_070_459, w_033_638, w_000_1268);
  and2 I070_463(w_070_463, w_025_1079, w_034_315);
  and2 I070_471(w_070_471, w_052_1058, w_059_565);
  or2  I070_472(w_070_472, w_020_518, w_004_1699);
  not1 I071_007(w_071_007, w_059_606);
  not1 I071_011(w_071_011, w_013_133);
  or2  I071_012(w_071_012, w_043_050, w_027_421);
  or2  I071_016(w_071_016, w_006_081, w_057_330);
  nand2 I071_018(w_071_018, w_003_257, w_059_096);
  not1 I071_025(w_071_025, w_069_760);
  not1 I071_028(w_071_028, w_062_027);
  not1 I071_033(w_071_033, w_039_1009);
  not1 I071_040(w_071_040, w_060_084);
  not1 I071_043(w_071_043, w_008_707);
  not1 I071_044(w_071_044, w_055_361);
  or2  I071_048(w_071_048, w_061_473, w_043_089);
  not1 I071_052(w_071_052, w_026_1512);
  and2 I071_056(w_071_056, w_029_164, w_068_141);
  not1 I071_061(w_071_061, w_022_197);
  not1 I071_064(w_071_064, w_004_1911);
  not1 I071_066(w_071_066, w_031_619);
  and2 I071_070(w_071_070, w_057_828, w_022_203);
  not1 I071_071(w_071_071, w_039_1611);
  not1 I071_082(w_071_082, w_004_739);
  not1 I071_086(w_071_086, w_004_266);
  nand2 I071_108(w_071_108, w_063_038, w_068_234);
  or2  I071_125(w_071_125, w_031_039, w_057_186);
  nand2 I071_130(w_071_130, w_057_1038, w_037_684);
  not1 I071_151(w_071_151, w_068_166);
  not1 I071_164(w_071_164, w_044_541);
  not1 I071_167(w_071_167, w_041_108);
  nand2 I071_191(w_071_191, w_038_454, w_004_305);
  not1 I071_193(w_071_193, w_034_669);
  and2 I071_202(w_071_202, w_041_254, w_006_227);
  and2 I071_224(w_071_224, w_036_454, w_002_411);
  and2 I071_227(w_071_227, w_064_1466, w_008_602);
  or2  I071_235(w_071_235, w_061_374, w_059_183);
  or2  I071_263(w_071_263, w_044_137, w_041_237);
  and2 I071_274(w_071_274, w_069_1681, w_037_1461);
  not1 I071_289(w_071_289, w_031_449);
  nand2 I071_293(w_071_293, w_052_1396, w_008_673);
  nand2 I071_295(w_071_295, w_068_160, w_029_509);
  or2  I071_303(w_071_303, w_050_562, w_019_097);
  nand2 I071_306(w_071_306, w_060_072, w_004_1778);
  nand2 I071_312(w_071_312, w_055_602, w_016_026);
  nand2 I071_323(w_071_323, w_070_062, w_028_301);
  nand2 I071_339(w_071_339, w_017_214, w_064_140);
  not1 I071_341(w_071_341, w_058_809);
  nand2 I071_355(w_071_355, w_019_222, w_039_313);
  and2 I071_357(w_071_357, w_057_239, w_026_103);
  not1 I071_358(w_071_358, w_057_936);
  not1 I071_361(w_071_361, w_059_296);
  nand2 I071_380(w_071_380, w_003_307, w_021_171);
  not1 I071_385(w_071_385, w_069_1723);
  nand2 I071_406(w_071_406, w_039_631, w_056_894);
  not1 I071_437(w_071_437, w_041_161);
  not1 I071_442(w_071_442, w_043_060);
  not1 I071_457(w_071_457, w_021_144);
  and2 I071_465(w_071_465, w_023_614, w_029_061);
  and2 I071_477(w_071_477, w_026_763, w_043_024);
  or2  I071_481(w_071_481, w_009_026, w_063_375);
  and2 I071_488(w_071_488, w_030_127, w_037_517);
  or2  I071_519(w_071_519, w_067_786, w_053_014);
  or2  I071_522(w_071_522, w_006_069, w_011_617);
  and2 I071_523(w_071_523, w_019_481, w_053_034);
  not1 I071_529(w_071_529, w_009_056);
  nand2 I071_531(w_071_531, w_038_457, w_056_1121);
  not1 I071_550(w_071_550, w_059_573);
  nand2 I072_001(w_072_001, w_044_175, w_034_558);
  nand2 I072_002(w_072_002, w_051_1068, w_046_131);
  nand2 I072_003(w_072_003, w_024_127, w_004_1280);
  and2 I072_005(w_072_005, w_028_266, w_043_011);
  nand2 I072_006(w_072_006, w_019_763, w_005_781);
  not1 I072_007(w_072_007, w_040_225);
  and2 I072_008(w_072_008, w_019_519, w_068_013);
  or2  I072_010(w_072_010, w_035_1267, w_017_1410);
  not1 I072_013(w_072_013, w_052_1549);
  or2  I072_019(w_072_019, w_001_1631, w_031_312);
  and2 I072_022(w_072_022, w_065_003, w_058_1469);
  not1 I072_024(w_072_024, w_066_086);
  nand2 I072_032(w_072_032, w_030_207, w_050_155);
  not1 I072_035(w_072_035, w_067_541);
  and2 I072_038(w_072_038, w_067_692, w_001_173);
  nand2 I072_040(w_072_040, w_015_081, w_048_409);
  or2  I072_042(w_072_042, w_025_209, w_034_066);
  nand2 I072_047(w_072_047, w_012_661, w_039_027);
  and2 I072_048(w_072_048, w_069_1365, w_014_014);
  nand2 I072_049(w_072_049, w_064_912, w_013_172);
  nand2 I072_051(w_072_051, w_068_209, w_032_013);
  and2 I072_052(w_072_052, w_053_116, w_054_620);
  nand2 I072_053(w_072_053, w_001_140, w_032_222);
  not1 I072_054(w_072_054, w_021_066);
  nand2 I072_055(w_072_055, w_051_581, w_034_371);
  nand2 I072_058(w_072_058, w_041_265, w_071_086);
  or2  I072_059(w_072_059, w_069_312, w_021_227);
  nand2 I072_066(w_072_066, w_070_180, w_046_028);
  nand2 I072_067(w_072_067, w_047_400, w_002_116);
  and2 I072_068(w_072_068, w_061_084, w_045_1878);
  nand2 I072_069(w_072_069, w_045_766, w_049_241);
  nand2 I072_070(w_072_070, w_005_770, w_005_1597);
  and2 I072_073(w_072_073, w_046_277, w_015_265);
  and2 I072_074(w_072_074, w_017_158, w_012_599);
  not1 I072_075(w_072_075, w_057_829);
  or2  I072_076(w_072_076, w_030_737, w_059_482);
  not1 I072_077(w_072_077, w_008_739);
  and2 I072_079(w_072_079, w_060_018, w_040_016);
  or2  I072_081(w_072_081, w_051_947, w_031_289);
  and2 I073_003(w_073_003, w_048_250, w_040_585);
  or2  I073_004(w_073_004, w_069_049, w_025_1287);
  and2 I073_005(w_073_005, w_009_075, w_040_365);
  and2 I073_006(w_073_006, w_022_302, w_033_1524);
  nand2 I073_008(w_073_008, w_019_558, w_040_1134);
  nand2 I073_009(w_073_009, w_018_211, w_020_028);
  nand2 I073_010(w_073_010, w_061_240, w_061_223);
  or2  I073_011(w_073_011, w_070_032, w_004_000);
  not1 I073_012(w_073_012, w_028_279);
  and2 I073_016(w_073_016, w_072_008, w_072_049);
  not1 I073_018(w_073_018, w_053_089);
  not1 I073_019(w_073_019, w_018_273);
  not1 I073_021(w_073_021, w_058_961);
  and2 I073_022(w_073_022, w_060_102, w_054_117);
  not1 I073_023(w_073_023, w_029_611);
  or2  I073_029(w_073_029, w_070_472, w_066_355);
  nand2 I073_030(w_073_030, w_038_387, w_067_206);
  and2 I073_031(w_073_031, w_008_407, w_070_387);
  or2  I073_034(w_073_034, w_021_003, w_057_1717);
  and2 I073_036(w_073_036, w_041_098, w_010_406);
  or2  I073_037(w_073_037, w_014_109, w_001_070);
  not1 I073_042(w_073_042, w_056_203);
  not1 I073_043(w_073_043, w_008_330);
  and2 I073_053(w_073_053, w_034_610, w_070_430);
  nand2 I073_059(w_073_059, w_016_002, w_008_143);
  not1 I073_061(w_073_061, w_001_510);
  and2 I073_062(w_073_062, w_015_022, w_028_767);
  not1 I073_063(w_073_063, w_003_126);
  nand2 I073_064(w_073_064, w_016_025, w_071_380);
  nand2 I073_065(w_073_065, w_070_260, w_037_328);
  nand2 I073_066(w_073_066, w_037_594, w_052_388);
  nand2 I073_067(w_073_067, w_022_346, w_028_355);
  nand2 I073_069(w_073_069, w_029_709, w_049_277);
  and2 I073_071(w_073_071, w_041_012, w_043_000);
  and2 I073_072(w_073_072, w_064_254, w_016_007);
  not1 I073_073(w_073_073, w_068_151);
  and2 I073_076(w_073_076, w_024_1133, w_071_061);
  or2  I073_079(w_073_079, w_027_308, w_032_211);
  nand2 I073_082(w_073_082, w_026_1186, w_053_116);
  nand2 I073_083(w_073_083, w_058_403, w_062_393);
  or2  I073_087(w_073_087, w_042_064, w_010_024);
  and2 I073_090(w_073_090, w_040_387, w_060_106);
  not1 I073_091(w_073_091, w_035_352);
  not1 I073_093(w_073_093, w_048_033);
  or2  I073_094(w_073_094, w_009_047, w_031_387);
  not1 I073_096(w_073_096, w_040_577);
  and2 I073_099(w_073_099, w_041_107, w_069_805);
  not1 I073_100(w_073_100, w_065_002);
  and2 I073_101(w_073_101, w_066_889, w_067_807);
  not1 I074_026(w_074_026, w_044_184);
  or2  I074_039(w_074_039, w_009_098, w_044_1446);
  not1 I074_054(w_074_054, w_011_742);
  and2 I074_059(w_074_059, w_059_210, w_032_138);
  or2  I074_080(w_074_080, w_042_046, w_053_091);
  and2 I074_115(w_074_115, w_035_103, w_011_403);
  nand2 I074_128(w_074_128, w_010_111, w_037_1132);
  and2 I074_129(w_074_129, w_067_403, w_027_437);
  nand2 I074_136(w_074_136, w_027_588, w_013_174);
  or2  I074_155(w_074_155, w_070_204, w_056_1615);
  not1 I074_167(w_074_167, w_071_016);
  not1 I074_169(w_074_169, w_014_366);
  nand2 I074_212(w_074_212, w_067_690, w_019_545);
  and2 I074_214(w_074_214, w_016_036, w_022_123);
  and2 I074_215(w_074_215, w_037_1103, w_014_165);
  and2 I074_219(w_074_219, w_033_528, w_030_225);
  and2 I074_231(w_074_231, w_003_263, w_030_313);
  and2 I074_241(w_074_241, w_069_568, w_056_018);
  not1 I074_246(w_074_246, w_063_725);
  and2 I074_262(w_074_262, w_035_050, w_018_139);
  and2 I074_273(w_074_273, w_047_059, w_004_646);
  or2  I074_274(w_074_274, w_018_148, w_026_1470);
  nand2 I074_278(w_074_278, w_003_045, w_018_052);
  or2  I074_295(w_074_295, w_055_233, w_053_063);
  and2 I074_298(w_074_298, w_020_369, w_047_548);
  or2  I074_357(w_074_357, w_005_647, w_022_316);
  or2  I074_422(w_074_422, w_059_403, w_036_880);
  nand2 I074_496(w_074_496, w_000_1914, w_060_058);
  and2 I074_501(w_074_501, w_069_976, w_032_126);
  or2  I074_551(w_074_551, w_018_212, w_060_041);
  not1 I074_557(w_074_557, w_032_051);
  and2 I074_558(w_074_558, w_014_506, w_004_030);
  or2  I074_582(w_074_582, w_038_276, w_055_261);
  and2 I074_583(w_074_583, w_067_080, w_046_074);
  not1 I074_584(w_074_584, w_048_649);
  or2  I074_625(w_074_625, w_035_104, w_040_832);
  not1 I074_658(w_074_658, w_068_018);
  or2  I074_680(w_074_680, w_050_1435, w_033_927);
  not1 I074_690(w_074_690, w_028_137);
  nand2 I074_713(w_074_713, w_017_1333, w_029_685);
  not1 I074_811(w_074_811, w_038_458);
  nand2 I074_869(w_074_869, w_032_231, w_069_1571);
  nand2 I074_954(w_074_954, w_027_308, w_027_007);
  not1 I074_961(w_074_961, w_005_044);
  not1 I074_1006(w_074_1006, w_005_155);
  nand2 I074_1023(w_074_1023, w_069_479, w_031_385);
  and2 I074_1032(w_074_1032, w_028_873, w_015_147);
  not1 I074_1077(w_074_1077, w_023_328);
  and2 I074_1109(w_074_1109, w_059_165, w_048_849);
  not1 I074_1217(w_074_1217, w_045_077);
  nand2 I074_1229(w_074_1229, w_016_015, w_013_052);
  nand2 I074_1230(w_074_1230, w_068_019, w_043_054);
  nand2 I074_1250(w_074_1250, w_037_1451, w_010_264);
  not1 I074_1265(w_074_1265, w_002_334);
  not1 I074_1283(w_074_1283, w_053_063);
  nand2 I074_1310(w_074_1310, w_032_122, w_005_207);
  and2 I074_1335(w_074_1335, w_008_109, w_008_431);
  nand2 I074_1365(w_074_1365, w_010_297, w_048_593);
  and2 I074_1427(w_074_1427, w_043_077, w_056_382);
  nand2 I074_1449(w_074_1449, w_004_846, w_042_141);
  and2 I074_1450(w_074_1450, w_037_446, w_036_435);
  nand2 I074_1467(w_074_1467, w_066_1093, w_072_070);
  or2  I074_1470(w_074_1470, w_057_1266, w_016_019);
  or2  I074_1501(w_074_1501, w_003_063, w_036_778);
  or2  I074_1578(w_074_1578, w_050_197, w_070_213);
  nand2 I074_1647(w_074_1647, w_021_246, w_064_609);
  nand2 I074_1683(w_074_1683, w_042_041, w_007_1269);
  not1 I074_1697(w_074_1697, w_033_805);
  and2 I075_000(w_075_000, w_059_080, w_023_1141);
  and2 I075_001(w_075_001, w_068_110, w_064_1594);
  and2 I075_003(w_075_003, w_038_325, w_043_053);
  not1 I075_005(w_075_005, w_012_008);
  or2  I075_014(w_075_014, w_050_044, w_051_853);
  and2 I075_025(w_075_025, w_014_361, w_008_751);
  and2 I075_037(w_075_037, w_000_537, w_073_037);
  nand2 I075_049(w_075_049, w_058_1762, w_043_057);
  or2  I075_051(w_075_051, w_034_612, w_016_003);
  nand2 I075_054(w_075_054, w_069_182, w_063_1375);
  nand2 I075_055(w_075_055, w_014_104, w_019_573);
  or2  I075_059(w_075_059, w_045_1659, w_062_972);
  not1 I075_061(w_075_061, w_006_014);
  not1 I075_062(w_075_062, w_025_262);
  or2  I075_065(w_075_065, w_056_086, w_007_547);
  and2 I075_071(w_075_071, w_009_000, w_059_289);
  not1 I075_074(w_075_074, w_026_1028);
  and2 I075_082(w_075_082, w_056_1468, w_039_1145);
  or2  I075_087(w_075_087, w_015_005, w_040_737);
  and2 I075_091(w_075_091, w_031_974, w_016_018);
  not1 I075_096(w_075_096, w_004_754);
  and2 I075_097(w_075_097, w_025_565, w_010_025);
  not1 I075_098(w_075_098, w_019_615);
  nand2 I075_105(w_075_105, w_033_245, w_058_919);
  nand2 I075_109(w_075_109, w_063_1604, w_016_006);
  nand2 I075_116(w_075_116, w_054_188, w_030_747);
  nand2 I075_117(w_075_117, w_032_053, w_033_634);
  nand2 I075_118(w_075_118, w_001_371, w_060_070);
  and2 I075_127(w_075_127, w_041_063, w_072_073);
  and2 I075_132(w_075_132, w_004_1133, w_026_325);
  and2 I075_144(w_075_144, w_031_529, w_065_003);
  and2 I075_151(w_075_151, w_003_202, w_055_155);
  or2  I075_152(w_075_152, w_057_1591, w_020_922);
  or2  I075_159(w_075_159, w_023_476, w_055_291);
  and2 I075_167(w_075_167, w_048_473, w_062_1158);
  or2  I075_172(w_075_172, w_013_320, w_010_040);
  not1 I075_173(w_075_173, w_033_283);
  not1 I075_174(w_075_174, w_058_097);
  or2  I075_179(w_075_179, w_047_060, w_042_014);
  or2  I075_184(w_075_184, w_037_713, w_070_004);
  not1 I075_187(w_075_187, w_049_377);
  and2 I075_213(w_075_213, w_025_730, w_004_201);
  not1 I075_214(w_075_214, w_000_1379);
  not1 I075_217(w_075_217, w_061_468);
  nand2 I075_221(w_075_221, w_039_1548, w_064_1238);
  not1 I075_231(w_075_231, w_054_492);
  not1 I075_234(w_075_234, w_038_473);
  nand2 I075_237(w_075_237, w_043_091, w_020_399);
  nand2 I075_238(w_075_238, w_018_248, w_034_410);
  nand2 I075_239(w_075_239, w_021_143, w_036_166);
  and2 I075_241(w_075_241, w_044_414, w_066_282);
  and2 I075_247(w_075_247, w_019_127, w_052_1588);
  and2 I075_249(w_075_249, w_020_843, w_023_266);
  nand2 I075_252(w_075_252, w_067_209, w_018_258);
  nand2 I075_254(w_075_254, w_068_189, w_014_829);
  or2  I075_257(w_075_257, w_059_172, w_012_578);
  or2  I075_261(w_075_261, w_067_512, w_019_800);
  nand2 I075_263(w_075_263, w_018_021, w_017_605);
  not1 I075_264(w_075_264, w_068_073);
  nand2 I075_266(w_075_266, w_015_008, w_052_844);
  or2  I075_282(w_075_282, w_041_037, w_067_962);
  or2  I076_006(w_076_006, w_001_473, w_029_998);
  and2 I076_010(w_076_010, w_052_1785, w_043_083);
  or2  I076_025(w_076_025, w_058_1743, w_072_066);
  nand2 I076_034(w_076_034, w_074_501, w_057_1646);
  not1 I076_039(w_076_039, w_005_1115);
  and2 I076_045(w_076_045, w_041_169, w_038_269);
  not1 I076_046(w_076_046, w_036_071);
  or2  I076_048(w_076_048, w_015_089, w_042_054);
  or2  I076_049(w_076_049, w_070_172, w_059_152);
  nand2 I076_057(w_076_057, w_056_1275, w_013_210);
  not1 I076_058(w_076_058, w_028_064);
  not1 I076_066(w_076_066, w_003_163);
  and2 I076_074(w_076_074, w_025_022, w_044_374);
  nand2 I076_076(w_076_076, w_055_057, w_036_580);
  and2 I076_078(w_076_078, w_041_264, w_013_325);
  nand2 I076_085(w_076_085, w_039_782, w_071_519);
  or2  I076_094(w_076_094, w_013_286, w_015_053);
  or2  I076_103(w_076_103, w_062_732, w_074_273);
  and2 I076_118(w_076_118, w_075_261, w_053_014);
  nand2 I076_119(w_076_119, w_039_1392, w_057_676);
  nand2 I076_120(w_076_120, w_019_397, w_057_709);
  nand2 I076_128(w_076_128, w_011_576, w_071_361);
  not1 I076_138(w_076_138, w_027_460);
  or2  I076_140(w_076_140, w_023_1292, w_048_850);
  or2  I076_146(w_076_146, w_055_828, w_022_233);
  nand2 I076_149(w_076_149, w_008_199, w_019_825);
  nand2 I076_155(w_076_155, w_074_690, w_030_124);
  and2 I076_169(w_076_169, w_035_999, w_052_1379);
  and2 I076_180(w_076_180, w_018_182, w_062_1016);
  and2 I076_200(w_076_200, w_050_161, w_038_196);
  or2  I076_203(w_076_203, w_028_061, w_063_016);
  and2 I076_208(w_076_208, w_043_029, w_008_778);
  and2 I076_209(w_076_209, w_020_572, w_017_804);
  not1 I076_210(w_076_210, w_004_778);
  or2  I076_211(w_076_211, w_037_982, w_007_996);
  and2 I076_215(w_076_215, w_060_060, w_024_186);
  and2 I076_240(w_076_240, w_024_038, w_055_253);
  or2  I076_242(w_076_242, w_034_424, w_061_055);
  nand2 I076_244(w_076_244, w_026_337, w_041_082);
  not1 I076_262(w_076_262, w_029_661);
  or2  I076_267(w_076_267, w_011_780, w_056_503);
  and2 I076_285(w_076_285, w_047_524, w_049_803);
  nand2 I076_288(w_076_288, w_011_353, w_075_062);
  or2  I076_290(w_076_290, w_057_1646, w_063_1088);
  and2 I076_296(w_076_296, w_027_481, w_073_034);
  nand2 I076_311(w_076_311, w_068_055, w_071_066);
  not1 I076_327(w_076_327, w_065_000);
  not1 I076_330(w_076_330, w_032_058);
  nand2 I076_333(w_076_333, w_020_448, w_064_190);
  or2  I076_335(w_076_335, w_002_419, w_025_553);
  or2  I076_338(w_076_338, w_040_813, w_035_908);
  or2  I076_344(w_076_344, w_036_1023, w_074_1023);
  or2  I076_354(w_076_354, w_068_240, w_003_203);
  and2 I076_355(w_076_355, w_066_213, w_018_120);
  or2  I076_356(w_076_356, w_064_1303, w_056_615);
  and2 I077_009(w_077_009, w_039_1600, w_027_287);
  and2 I077_014(w_077_014, w_020_772, w_002_317);
  or2  I077_023(w_077_023, w_044_022, w_045_290);
  and2 I077_034(w_077_034, w_002_224, w_040_165);
  nand2 I077_055(w_077_055, w_008_250, w_054_535);
  not1 I077_134(w_077_134, w_041_258);
  nand2 I077_151(w_077_151, w_013_300, w_012_373);
  or2  I077_153(w_077_153, w_040_938, w_060_094);
  not1 I077_170(w_077_170, w_023_364);
  nand2 I077_174(w_077_174, w_026_170, w_067_582);
  or2  I077_197(w_077_197, w_064_631, w_015_052);
  and2 I077_201(w_077_201, w_068_106, w_046_148);
  and2 I077_209(w_077_209, w_071_011, w_025_1042);
  not1 I077_223(w_077_223, w_048_415);
  or2  I077_232(w_077_232, w_000_1224, w_052_1856);
  not1 I077_238(w_077_238, w_059_360);
  not1 I077_252(w_077_252, w_014_726);
  nand2 I077_310(w_077_310, w_054_086, w_029_837);
  not1 I077_314(w_077_314, w_065_003);
  not1 I077_438(w_077_438, w_075_087);
  and2 I077_439(w_077_439, w_047_419, w_048_326);
  nand2 I077_460(w_077_460, w_050_420, w_065_001);
  or2  I077_490(w_077_490, w_063_1265, w_036_1457);
  nand2 I077_494(w_077_494, w_043_096, w_025_1572);
  not1 I077_526(w_077_526, w_033_1406);
  and2 I077_540(w_077_540, w_047_372, w_064_941);
  not1 I077_568(w_077_568, w_019_516);
  or2  I077_571(w_077_571, w_059_361, w_028_595);
  and2 I077_589(w_077_589, w_035_217, w_064_145);
  not1 I077_596(w_077_596, w_046_124);
  nand2 I077_602(w_077_602, w_016_028, w_010_320);
  nand2 I077_623(w_077_623, w_008_297, w_005_162);
  not1 I077_632(w_077_632, w_052_857);
  and2 I077_642(w_077_642, w_031_752, w_016_028);
  or2  I077_658(w_077_658, w_046_040, w_039_1932);
  and2 I077_664(w_077_664, w_059_206, w_055_598);
  or2  I077_701(w_077_701, w_050_1052, w_013_291);
  not1 I077_702(w_077_702, w_063_1251);
  nand2 I077_709(w_077_709, w_048_440, w_019_287);
  and2 I077_725(w_077_725, w_002_315, w_050_552);
  not1 I077_769(w_077_769, w_004_1566);
  nand2 I077_798(w_077_798, w_029_614, w_036_866);
  nand2 I077_873(w_077_873, w_046_147, w_025_1698);
  nand2 I077_895(w_077_895, w_056_085, w_006_007);
  nand2 I077_903(w_077_903, w_055_128, w_051_559);
  or2  I077_914(w_077_914, w_025_102, w_060_037);
  nand2 I077_927(w_077_927, w_036_939, w_071_052);
  or2  I077_945(w_077_945, w_005_1268, w_070_093);
  and2 I077_997(w_077_997, w_018_165, w_013_226);
  not1 I077_1006(w_077_1006, w_065_005);
  nand2 I077_1084(w_077_1084, w_072_068, w_042_072);
  not1 I077_1107(w_077_1107, w_041_194);
  nand2 I077_1114(w_077_1114, w_043_005, w_054_444);
  and2 I077_1148(w_077_1148, w_060_018, w_009_054);
  not1 I078_019(w_078_019, w_057_1768);
  or2  I078_037(w_078_037, w_055_772, w_001_525);
  or2  I078_048(w_078_048, w_004_362, w_029_193);
  not1 I078_053(w_078_053, w_058_1500);
  not1 I078_055(w_078_055, w_041_118);
  nand2 I078_088(w_078_088, w_037_1528, w_007_272);
  and2 I078_089(w_078_089, w_030_207, w_028_647);
  nand2 I078_092(w_078_092, w_048_554, w_023_937);
  and2 I078_093(w_078_093, w_032_144, w_037_1149);
  nand2 I078_103(w_078_103, w_044_342, w_002_547);
  not1 I078_109(w_078_109, w_068_037);
  not1 I078_113(w_078_113, w_064_193);
  nand2 I078_148(w_078_148, w_072_022, w_068_233);
  nand2 I078_195(w_078_195, w_015_248, w_014_029);
  or2  I078_205(w_078_205, w_049_289, w_028_495);
  nand2 I078_217(w_078_217, w_005_433, w_054_102);
  or2  I078_218(w_078_218, w_058_1629, w_026_771);
  not1 I078_236(w_078_236, w_007_1045);
  or2  I078_252(w_078_252, w_014_214, w_041_232);
  not1 I078_261(w_078_261, w_011_883);
  and2 I078_281(w_078_281, w_062_271, w_039_1213);
  and2 I078_285(w_078_285, w_067_898, w_054_365);
  not1 I078_287(w_078_287, w_003_197);
  nand2 I078_289(w_078_289, w_017_615, w_001_406);
  not1 I078_347(w_078_347, w_045_710);
  not1 I078_349(w_078_349, w_023_1596);
  and2 I078_353(w_078_353, w_005_084, w_031_509);
  nand2 I078_434(w_078_434, w_048_479, w_035_152);
  and2 I078_455(w_078_455, w_075_054, w_071_071);
  or2  I078_479(w_078_479, w_003_101, w_020_582);
  nand2 I078_500(w_078_500, w_008_163, w_003_226);
  not1 I078_538(w_078_538, w_002_217);
  and2 I078_557(w_078_557, w_074_1467, w_010_064);
  nand2 I078_632(w_078_632, w_038_333, w_047_031);
  not1 I078_636(w_078_636, w_045_1488);
  and2 I078_723(w_078_723, w_036_143, w_041_059);
  not1 I078_747(w_078_747, w_050_1147);
  and2 I078_778(w_078_778, w_034_144, w_018_150);
  or2  I078_801(w_078_801, w_061_375, w_070_061);
  not1 I078_829(w_078_829, w_065_000);
  nand2 I078_835(w_078_835, w_020_338, w_005_006);
  not1 I078_854(w_078_854, w_020_292);
  not1 I078_863(w_078_863, w_045_1086);
  nand2 I078_864(w_078_864, w_060_104, w_076_146);
  and2 I078_865(w_078_865, w_018_229, w_019_671);
  not1 I078_872(w_078_872, w_032_086);
  nand2 I078_884(w_078_884, w_058_041, w_012_172);
  or2  I078_937(w_078_937, w_067_418, w_047_558);
  and2 I078_969(w_078_969, w_034_620, w_062_362);
  nand2 I078_995(w_078_995, w_063_706, w_056_589);
  and2 I078_1036(w_078_1036, w_077_602, w_037_901);
  and2 I078_1042(w_078_1042, w_024_342, w_018_138);
  or2  I078_1120(w_078_1120, w_032_164, w_043_034);
  and2 I078_1150(w_078_1150, w_025_099, w_024_559);
  not1 I078_1153(w_078_1153, w_048_974);
  and2 I078_1155(w_078_1155, w_045_1313, w_077_134);
  or2  I078_1184(w_078_1184, w_064_455, w_035_149);
  nand2 I078_1276(w_078_1276, w_008_268, w_044_324);
  and2 I078_1286(w_078_1286, w_002_586, w_026_1297);
  and2 I078_1342(w_078_1342, w_002_246, w_061_538);
  nand2 I078_1347(w_078_1347, w_026_227, w_001_288);
  nand2 I078_1349(w_078_1349, w_032_216, w_003_022);
  nand2 I078_1352(w_078_1352, w_032_056, w_016_034);
  or2  I078_1362(w_078_1362, w_015_205, w_002_130);
  not1 I078_1469(w_078_1469, w_060_033);
  not1 I078_1496(w_078_1496, w_002_281);
  nand2 I078_1506(w_078_1506, w_033_1498, w_018_056);
  or2  I078_1631(w_078_1631, w_046_127, w_044_1781);
  nand2 I078_1664(w_078_1664, w_047_387, w_003_036);
  and2 I078_1688(w_078_1688, w_050_597, w_058_1589);
  not1 I079_005(w_079_005, w_064_210);
  or2  I079_015(w_079_015, w_053_077, w_044_309);
  nand2 I079_018(w_079_018, w_044_908, w_056_800);
  and2 I079_020(w_079_020, w_060_103, w_035_1234);
  or2  I079_030(w_079_030, w_041_171, w_068_059);
  not1 I079_034(w_079_034, w_015_119);
  not1 I079_048(w_079_048, w_014_340);
  not1 I079_078(w_079_078, w_038_339);
  nand2 I079_094(w_079_094, w_065_003, w_035_064);
  nand2 I079_104(w_079_104, w_038_112, w_074_558);
  and2 I079_112(w_079_112, w_030_222, w_044_1639);
  nand2 I079_115(w_079_115, w_033_423, w_052_566);
  and2 I079_126(w_079_126, w_001_282, w_073_009);
  nand2 I079_128(w_079_128, w_008_732, w_029_383);
  not1 I079_134(w_079_134, w_020_423);
  and2 I079_142(w_079_142, w_078_479, w_076_203);
  not1 I079_145(w_079_145, w_002_071);
  nand2 I079_159(w_079_159, w_029_1109, w_000_1760);
  or2  I079_162(w_079_162, w_001_1631, w_078_1631);
  and2 I079_176(w_079_176, w_070_149, w_025_766);
  nand2 I079_202(w_079_202, w_053_116, w_022_206);
  or2  I079_216(w_079_216, w_000_741, w_024_439);
  and2 I079_218(w_079_218, w_046_079, w_014_159);
  nand2 I079_233(w_079_233, w_002_190, w_040_172);
  nand2 I079_261(w_079_261, w_045_1650, w_019_144);
  nand2 I079_270(w_079_270, w_072_003, w_060_088);
  or2  I079_293(w_079_293, w_024_310, w_017_1443);
  and2 I079_321(w_079_321, w_070_448, w_037_028);
  or2  I079_363(w_079_363, w_014_119, w_023_1105);
  and2 I079_374(w_079_374, w_055_162, w_047_500);
  nand2 I079_382(w_079_382, w_030_533, w_069_068);
  or2  I079_395(w_079_395, w_077_914, w_014_442);
  and2 I079_411(w_079_411, w_025_897, w_052_405);
  and2 I079_425(w_079_425, w_001_893, w_045_805);
  and2 I079_463(w_079_463, w_048_551, w_021_148);
  not1 I079_502(w_079_502, w_054_251);
  or2  I079_526(w_079_526, w_019_240, w_017_442);
  or2  I079_536(w_079_536, w_066_574, w_004_1864);
  or2  I079_539(w_079_539, w_054_509, w_004_1746);
  not1 I079_556(w_079_556, w_033_090);
  nand2 I079_564(w_079_564, w_065_002, w_035_976);
  nand2 I079_568(w_079_568, w_049_447, w_005_226);
  and2 I079_573(w_079_573, w_015_010, w_064_889);
  and2 I079_577(w_079_577, w_051_643, w_066_154);
  or2  I079_578(w_079_578, w_034_350, w_065_002);
  not1 I079_588(w_079_588, w_050_1218);
  or2  I079_598(w_079_598, w_026_451, w_034_009);
  or2  I079_612(w_079_612, w_036_1153, w_052_1264);
  not1 I079_622(w_079_622, w_003_140);
  not1 I079_640(w_079_640, w_026_1520);
  not1 I079_649(w_079_649, w_023_702);
  not1 I079_651(w_079_651, w_074_961);
  or2  I079_667(w_079_667, w_042_129, w_075_174);
  nand2 I079_718(w_079_718, w_074_1365, w_021_112);
  or2  I079_721(w_079_721, w_010_203, w_010_003);
  and2 I079_747(w_079_747, w_058_431, w_021_132);
  nand2 I079_748(w_079_748, w_001_032, w_031_292);
  or2  I079_753(w_079_753, w_035_997, w_059_435);
  and2 I079_784(w_079_784, w_010_171, w_025_088);
  not1 I079_789(w_079_789, w_075_071);
  nand2 I079_797(w_079_797, w_031_061, w_016_013);
  and2 I079_819(w_079_819, w_031_842, w_015_034);
  nand2 I079_839(w_079_839, w_003_095, w_021_049);
  or2  I079_847(w_079_847, w_032_090, w_000_1569);
  nand2 I079_848(w_079_848, w_000_1695, w_027_176);
  nand2 I080_000(w_080_000, w_056_727, w_019_597);
  or2  I080_001(w_080_001, w_037_998, w_068_041);
  nand2 I080_007(w_080_007, w_007_1595, w_051_440);
  not1 I080_008(w_080_008, w_008_296);
  not1 I080_010(w_080_010, w_022_150);
  and2 I080_013(w_080_013, w_053_117, w_055_526);
  and2 I080_018(w_080_018, w_065_003, w_067_287);
  and2 I080_019(w_080_019, w_052_1394, w_045_666);
  or2  I080_021(w_080_021, w_038_484, w_057_645);
  nand2 I080_024(w_080_024, w_054_479, w_031_619);
  not1 I080_028(w_080_028, w_074_262);
  or2  I080_030(w_080_030, w_058_1424, w_066_702);
  nand2 I080_034(w_080_034, w_055_300, w_041_010);
  and2 I080_036(w_080_036, w_062_608, w_052_640);
  and2 I080_040(w_080_040, w_014_696, w_002_340);
  and2 I080_048(w_080_048, w_041_155, w_055_660);
  and2 I080_049(w_080_049, w_014_489, w_021_080);
  or2  I080_050(w_080_050, w_026_874, w_079_649);
  or2  I080_051(w_080_051, w_055_852, w_048_567);
  not1 I080_059(w_080_059, w_031_217);
  or2  I080_061(w_080_061, w_051_947, w_000_1279);
  not1 I080_067(w_080_067, w_068_239);
  nand2 I080_068(w_080_068, w_040_411, w_015_195);
  or2  I080_069(w_080_069, w_066_373, w_046_082);
  nand2 I080_070(w_080_070, w_023_527, w_054_518);
  nand2 I080_077(w_080_077, w_040_272, w_039_1551);
  and2 I080_082(w_080_082, w_027_144, w_065_002);
  not1 I080_090(w_080_090, w_049_871);
  or2  I080_095(w_080_095, w_072_003, w_025_1529);
  nand2 I080_096(w_080_096, w_000_155, w_004_292);
  and2 I080_099(w_080_099, w_064_147, w_060_030);
  nand2 I080_102(w_080_102, w_065_005, w_067_905);
  and2 I080_103(w_080_103, w_029_047, w_044_1224);
  or2  I080_105(w_080_105, w_016_003, w_059_577);
  nand2 I080_106(w_080_106, w_075_221, w_067_288);
  nand2 I080_109(w_080_109, w_071_033, w_059_692);
  or2  I080_110(w_080_110, w_055_169, w_000_1064);
  nand2 I080_111(w_080_111, w_009_020, w_025_377);
  not1 I080_112(w_080_112, w_004_955);
  not1 I080_114(w_080_114, w_050_032);
  not1 I080_115(w_080_115, w_073_042);
  not1 I080_118(w_080_118, w_013_162);
  nand2 I080_119(w_080_119, w_013_258, w_051_768);
  not1 I081_028(w_081_028, w_009_070);
  and2 I081_040(w_081_040, w_049_206, w_066_714);
  or2  I081_050(w_081_050, w_023_265, w_056_1184);
  not1 I081_055(w_081_055, w_001_476);
  not1 I081_059(w_081_059, w_062_618);
  not1 I081_077(w_081_077, w_080_114);
  nand2 I081_086(w_081_086, w_074_054, w_043_021);
  nand2 I081_093(w_081_093, w_076_330, w_039_1496);
  or2  I081_095(w_081_095, w_051_939, w_062_587);
  and2 I081_107(w_081_107, w_044_777, w_016_007);
  and2 I081_142(w_081_142, w_016_024, w_065_005);
  and2 I081_162(w_081_162, w_071_263, w_020_821);
  not1 I081_183(w_081_183, w_064_772);
  not1 I081_208(w_081_208, w_036_196);
  or2  I081_221(w_081_221, w_079_115, w_000_1829);
  not1 I081_223(w_081_223, w_011_201);
  not1 I081_242(w_081_242, w_033_067);
  or2  I081_249(w_081_249, w_069_1731, w_004_1511);
  nand2 I081_290(w_081_290, w_075_051, w_000_528);
  not1 I081_311(w_081_311, w_030_491);
  and2 I081_341(w_081_341, w_038_480, w_039_1890);
  and2 I081_354(w_081_354, w_013_059, w_011_224);
  not1 I081_377(w_081_377, w_021_128);
  or2  I081_385(w_081_385, w_045_1833, w_045_065);
  nand2 I081_392(w_081_392, w_068_164, w_026_435);
  and2 I081_407(w_081_407, w_038_181, w_021_159);
  and2 I081_415(w_081_415, w_078_1150, w_014_565);
  or2  I081_416(w_081_416, w_002_539, w_043_103);
  not1 I081_430(w_081_430, w_009_068);
  or2  I081_437(w_081_437, w_047_262, w_014_366);
  not1 I081_447(w_081_447, w_064_1064);
  not1 I081_468(w_081_468, w_049_1033);
  or2  I081_480(w_081_480, w_057_277, w_073_094);
  not1 I081_481(w_081_481, w_022_066);
  nand2 I081_490(w_081_490, w_043_032, w_078_148);
  or2  I081_532(w_081_532, w_067_799, w_064_234);
  or2  I081_539(w_081_539, w_008_316, w_035_1527);
  or2  I081_558(w_081_558, w_056_1223, w_046_017);
  or2  I081_560(w_081_560, w_042_104, w_061_582);
  or2  I081_571(w_081_571, w_005_1300, w_068_011);
  or2  I081_572(w_081_572, w_002_297, w_068_114);
  not1 I081_576(w_081_576, w_022_280);
  and2 I081_578(w_081_578, w_078_037, w_020_355);
  or2  I081_582(w_081_582, w_077_238, w_045_1139);
  nand2 I081_619(w_081_619, w_054_172, w_079_218);
  or2  I081_647(w_081_647, w_028_342, w_045_1551);
  and2 I081_663(w_081_663, w_027_167, w_064_1046);
  not1 I081_665(w_081_665, w_043_019);
  nand2 I081_669(w_081_669, w_009_048, w_053_109);
  or2  I081_678(w_081_678, w_080_040, w_030_042);
  nand2 I082_083(w_082_083, w_005_457, w_018_278);
  and2 I082_092(w_082_092, w_002_567, w_027_186);
  and2 I082_095(w_082_095, w_078_289, w_030_695);
  nand2 I082_099(w_082_099, w_061_546, w_027_159);
  nand2 I082_115(w_082_115, w_070_270, w_015_267);
  not1 I082_120(w_082_120, w_013_230);
  nand2 I082_155(w_082_155, w_069_970, w_026_521);
  not1 I082_179(w_082_179, w_024_297);
  or2  I082_193(w_082_193, w_048_007, w_029_1118);
  nand2 I082_233(w_082_233, w_069_019, w_003_214);
  or2  I082_240(w_082_240, w_035_644, w_029_1091);
  and2 I082_260(w_082_260, w_007_1531, w_060_097);
  nand2 I082_262(w_082_262, w_081_392, w_016_000);
  nand2 I082_265(w_082_265, w_050_1164, w_076_335);
  and2 I082_275(w_082_275, w_005_094, w_023_1398);
  or2  I082_303(w_082_303, w_051_126, w_064_1435);
  not1 I082_314(w_082_314, w_064_039);
  nand2 I082_337(w_082_337, w_070_450, w_048_230);
  and2 I082_341(w_082_341, w_003_158, w_036_813);
  or2  I082_358(w_082_358, w_017_1041, w_030_073);
  nand2 I082_382(w_082_382, w_063_184, w_028_132);
  not1 I082_409(w_082_409, w_007_377);
  not1 I082_414(w_082_414, w_078_865);
  and2 I082_422(w_082_422, w_046_075, w_064_1150);
  nand2 I082_423(w_082_423, w_012_162, w_020_994);
  and2 I082_426(w_082_426, w_072_042, w_034_419);
  not1 I082_431(w_082_431, w_004_1038);
  not1 I082_466(w_082_466, w_043_084);
  nand2 I082_500(w_082_500, w_019_459, w_012_210);
  not1 I082_507(w_082_507, w_077_014);
  and2 I082_510(w_082_510, w_076_242, w_069_053);
  not1 I082_515(w_082_515, w_049_606);
  not1 I082_517(w_082_517, w_040_260);
  not1 I082_527(w_082_527, w_036_179);
  or2  I082_529(w_082_529, w_007_1405, w_080_118);
  not1 I082_549(w_082_549, w_060_003);
  nand2 I082_586(w_082_586, w_020_1225, w_063_1173);
  not1 I082_589(w_082_589, w_010_090);
  not1 I082_593(w_082_593, w_070_014);
  or2  I082_597(w_082_597, w_043_042, w_019_619);
  not1 I082_649(w_082_649, w_035_1513);
  nand2 I082_658(w_082_658, w_034_462, w_040_679);
  not1 I082_688(w_082_688, w_016_026);
  nand2 I082_691(w_082_691, w_010_355, w_034_178);
  and2 I082_698(w_082_698, w_010_308, w_068_135);
  nand2 I082_721(w_082_721, w_056_1064, w_042_102);
  nand2 I082_734(w_082_734, w_076_025, w_027_008);
  and2 I082_745(w_082_745, w_070_455, w_011_135);
  and2 I082_782(w_082_782, w_050_1344, w_017_1400);
  nand2 I082_799(w_082_799, w_063_016, w_023_666);
  or2  I082_808(w_082_808, w_017_1179, w_032_155);
  nand2 I082_813(w_082_813, w_010_110, w_075_214);
  not1 I083_000(w_083_000, w_028_157);
  or2  I083_001(w_083_001, w_001_224, w_022_268);
  nand2 I083_002(w_083_002, w_063_1294, w_037_1108);
  not1 I083_003(w_083_003, w_031_004);
  nand2 I083_004(w_083_004, w_078_1276, w_053_001);
  and2 I083_005(w_083_005, w_082_586, w_022_032);
  and2 I083_006(w_083_006, w_025_061, w_018_213);
  and2 I083_007(w_083_007, w_050_069, w_015_261);
  nand2 I083_008(w_083_008, w_038_486, w_041_152);
  and2 I083_010(w_083_010, w_016_011, w_045_338);
  not1 I083_011(w_083_011, w_062_436);
  not1 I083_013(w_083_013, w_030_172);
  or2  I083_014(w_083_014, w_006_238, w_020_379);
  nand2 I083_015(w_083_015, w_071_341, w_027_044);
  and2 I083_016(w_083_016, w_048_345, w_051_1073);
  nand2 I083_017(w_083_017, w_001_192, w_016_016);
  nand2 I083_019(w_083_019, w_039_135, w_074_1449);
  or2  I083_020(w_083_020, w_044_1386, w_063_373);
  or2  I083_021(w_083_021, w_053_044, w_045_1824);
  not1 I083_022(w_083_022, w_015_152);
  nand2 I083_023(w_083_023, w_070_034, w_011_225);
  or2  I083_024(w_083_024, w_027_507, w_082_698);
  and2 I083_025(w_083_025, w_037_778, w_045_424);
  not1 I083_026(w_083_026, w_037_119);
  and2 I083_028(w_083_028, w_068_078, w_066_162);
  nand2 I083_029(w_083_029, w_001_098, w_017_397);
  and2 I083_030(w_083_030, w_028_622, w_002_546);
  not1 I083_031(w_083_031, w_005_449);
  nand2 I084_012(w_084_012, w_075_214, w_043_039);
  nand2 I084_013(w_084_013, w_059_318, w_082_099);
  not1 I084_016(w_084_016, w_043_010);
  not1 I084_019(w_084_019, w_026_022);
  nand2 I084_036(w_084_036, w_038_239, w_081_354);
  and2 I084_041(w_084_041, w_057_1599, w_042_086);
  or2  I084_050(w_084_050, w_032_152, w_077_540);
  and2 I084_055(w_084_055, w_057_276, w_039_1654);
  and2 I084_058(w_084_058, w_052_825, w_050_1119);
  not1 I084_065(w_084_065, w_079_839);
  or2  I084_070(w_084_070, w_060_094, w_081_050);
  and2 I084_071(w_084_071, w_026_995, w_066_845);
  and2 I084_073(w_084_073, w_007_223, w_053_050);
  and2 I084_079(w_084_079, w_047_226, w_081_480);
  and2 I084_080(w_084_080, w_003_115, w_059_017);
  not1 I084_091(w_084_091, w_019_814);
  not1 I084_123(w_084_123, w_046_226);
  not1 I084_139(w_084_139, w_065_000);
  not1 I084_142(w_084_142, w_081_107);
  nand2 I084_144(w_084_144, w_018_035, w_032_050);
  and2 I084_158(w_084_158, w_024_741, w_080_069);
  or2  I084_164(w_084_164, w_024_1465, w_026_620);
  nand2 I084_168(w_084_168, w_049_1075, w_067_544);
  or2  I084_197(w_084_197, w_006_105, w_021_025);
  and2 I084_207(w_084_207, w_004_544, w_072_048);
  not1 I084_211(w_084_211, w_072_007);
  not1 I084_233(w_084_233, w_073_076);
  not1 I084_260(w_084_260, w_073_062);
  nand2 I084_267(w_084_267, w_072_052, w_038_464);
  not1 I084_270(w_084_270, w_067_185);
  not1 I084_271(w_084_271, w_018_134);
  or2  I084_275(w_084_275, w_062_544, w_035_608);
  and2 I084_304(w_084_304, w_043_088, w_057_854);
  and2 I084_314(w_084_314, w_002_308, w_051_633);
  nand2 I084_315(w_084_315, w_039_1597, w_059_395);
  nand2 I084_317(w_084_317, w_045_213, w_053_033);
  or2  I084_333(w_084_333, w_030_302, w_060_063);
  nand2 I084_334(w_084_334, w_011_550, w_046_014);
  not1 I084_343(w_084_343, w_076_058);
  or2  I084_351(w_084_351, w_066_307, w_012_552);
  and2 I084_362(w_084_362, w_025_580, w_035_1041);
  nand2 I084_364(w_084_364, w_071_358, w_013_109);
  or2  I084_366(w_084_366, w_003_153, w_000_1039);
  nand2 I084_367(w_084_367, w_047_129, w_035_1023);
  or2  I084_375(w_084_375, w_062_106, w_009_070);
  and2 I084_379(w_084_379, w_023_026, w_051_273);
  nand2 I084_385(w_084_385, w_036_713, w_043_013);
  or2  I084_391(w_084_391, w_047_119, w_077_571);
  nand2 I084_405(w_084_405, w_045_023, w_039_805);
  not1 I084_410(w_084_410, w_076_120);
  nand2 I084_418(w_084_418, w_052_058, w_074_214);
  and2 I084_458(w_084_458, w_027_430, w_024_1066);
  not1 I084_470(w_084_470, w_065_003);
  and2 I084_474(w_084_474, w_059_084, w_056_751);
  nand2 I084_481(w_084_481, w_081_490, w_040_1352);
  nand2 I084_483(w_084_483, w_077_1006, w_037_055);
  not1 I085_001(w_085_001, w_026_1289);
  and2 I085_030(w_085_030, w_019_975, w_082_500);
  or2  I085_033(w_085_033, w_008_069, w_013_049);
  nand2 I085_046(w_085_046, w_014_805, w_024_1385);
  or2  I085_058(w_085_058, w_084_270, w_004_047);
  and2 I085_059(w_085_059, w_078_048, w_004_008);
  not1 I085_064(w_085_064, w_006_056);
  and2 I085_071(w_085_071, w_074_219, w_067_531);
  and2 I085_081(w_085_081, w_018_067, w_003_217);
  nand2 I085_098(w_085_098, w_078_863, w_083_006);
  not1 I085_099(w_085_099, w_061_337);
  nand2 I085_108(w_085_108, w_020_465, w_018_275);
  nand2 I085_109(w_085_109, w_026_665, w_003_016);
  and2 I085_111(w_085_111, w_059_184, w_069_723);
  or2  I085_115(w_085_115, w_049_595, w_040_1125);
  and2 I085_122(w_085_122, w_079_789, w_007_1594);
  and2 I085_127(w_085_127, w_019_001, w_082_721);
  or2  I085_134(w_085_134, w_035_052, w_004_488);
  and2 I085_135(w_085_135, w_031_194, w_034_022);
  and2 I085_146(w_085_146, w_034_674, w_060_031);
  not1 I085_153(w_085_153, w_026_1123);
  or2  I085_177(w_085_177, w_055_036, w_031_789);
  and2 I085_181(w_085_181, w_031_658, w_038_021);
  nand2 I085_184(w_085_184, w_081_341, w_045_1467);
  or2  I085_200(w_085_200, w_045_1507, w_082_782);
  and2 I085_201(w_085_201, w_080_077, w_060_097);
  and2 I085_204(w_085_204, w_008_709, w_044_1209);
  not1 I085_221(w_085_221, w_021_277);
  not1 I085_254(w_085_254, w_080_082);
  not1 I085_256(w_085_256, w_045_1538);
  and2 I085_270(w_085_270, w_014_434, w_083_011);
  and2 I085_274(w_085_274, w_055_094, w_047_518);
  or2  I085_302(w_085_302, w_036_137, w_001_1366);
  nand2 I085_314(w_085_314, w_030_239, w_058_1050);
  nand2 I085_355(w_085_355, w_000_627, w_008_538);
  nand2 I085_357(w_085_357, w_050_162, w_041_037);
  or2  I085_363(w_085_363, w_074_1310, w_017_1885);
  nand2 I085_373(w_085_373, w_069_920, w_065_000);
  not1 I085_385(w_085_385, w_082_314);
  and2 I085_388(w_085_388, w_066_332, w_064_1362);
  or2  I085_395(w_085_395, w_036_456, w_033_649);
  nand2 I085_418(w_085_418, w_021_116, w_009_074);
  or2  I085_427(w_085_427, w_004_626, w_008_163);
  or2  I085_439(w_085_439, w_046_136, w_037_1128);
  or2  I085_454(w_085_454, w_029_399, w_032_106);
  not1 I085_486(w_085_486, w_053_042);
  and2 I085_490(w_085_490, w_001_487, w_055_087);
  nand2 I085_496(w_085_496, w_054_073, w_048_553);
  or2  I085_505(w_085_505, w_041_127, w_050_362);
  not1 I085_511(w_085_511, w_069_1167);
  or2  I085_513(w_085_513, w_063_129, w_006_104);
  nand2 I085_522(w_085_522, w_076_076, w_064_1094);
  and2 I085_536(w_085_536, w_046_098, w_016_016);
  not1 I085_568(w_085_568, w_058_034);
  and2 I085_571(w_085_571, w_006_027, w_073_019);
  not1 I085_576(w_085_576, w_036_256);
  and2 I085_593(w_085_593, w_040_307, w_004_1120);
  and2 I085_602(w_085_602, w_045_171, w_002_111);
  and2 I085_607(w_085_607, w_017_666, w_066_324);
  nand2 I085_609(w_085_609, w_029_637, w_055_373);
  or2  I085_653(w_085_653, w_045_1486, w_031_409);
  nand2 I085_660(w_085_660, w_030_745, w_068_027);
  or2  I085_676(w_085_676, w_069_038, w_035_1255);
  or2  I086_025(w_086_025, w_076_180, w_072_032);
  not1 I086_044(w_086_044, w_036_972);
  or2  I086_049(w_086_049, w_027_578, w_081_407);
  nand2 I086_055(w_086_055, w_024_444, w_015_055);
  or2  I086_066(w_086_066, w_059_093, w_033_605);
  or2  I086_095(w_086_095, w_073_063, w_001_1449);
  and2 I086_096(w_086_096, w_063_1583, w_049_1129);
  not1 I086_108(w_086_108, w_032_141);
  nand2 I086_119(w_086_119, w_071_052, w_001_1662);
  and2 I086_160(w_086_160, w_006_260, w_059_492);
  or2  I086_166(w_086_166, w_065_005, w_048_432);
  or2  I086_176(w_086_176, w_026_860, w_071_130);
  not1 I086_178(w_086_178, w_084_385);
  not1 I086_203(w_086_203, w_050_1200);
  not1 I086_235(w_086_235, w_043_043);
  not1 I086_267(w_086_267, w_049_306);
  and2 I086_288(w_086_288, w_048_054, w_076_034);
  and2 I086_291(w_086_291, w_081_571, w_078_1362);
  nand2 I086_301(w_086_301, w_010_212, w_042_060);
  or2  I086_326(w_086_326, w_064_563, w_061_293);
  or2  I086_342(w_086_342, w_030_059, w_003_151);
  or2  I086_370(w_086_370, w_055_443, w_027_143);
  not1 I086_371(w_086_371, w_063_1594);
  or2  I086_402(w_086_402, w_051_501, w_020_546);
  nand2 I086_515(w_086_515, w_056_1269, w_080_102);
  and2 I086_539(w_086_539, w_059_052, w_061_151);
  nand2 I086_555(w_086_555, w_016_009, w_079_622);
  or2  I086_569(w_086_569, w_031_1065, w_076_262);
  nand2 I086_633(w_086_633, w_071_070, w_049_077);
  and2 I086_652(w_086_652, w_026_374, w_017_1448);
  and2 I086_677(w_086_677, w_082_517, w_023_043);
  nand2 I086_742(w_086_742, w_017_171, w_000_916);
  not1 I086_748(w_086_748, w_043_082);
  not1 I086_755(w_086_755, w_056_1671);
  or2  I086_780(w_086_780, w_003_054, w_069_1369);
  or2  I086_812(w_086_812, w_074_026, w_014_167);
  nand2 I086_838(w_086_838, w_073_091, w_036_169);
  nand2 I086_896(w_086_896, w_006_075, w_003_135);
  and2 I086_909(w_086_909, w_032_212, w_048_548);
  and2 I086_923(w_086_923, w_070_285, w_023_154);
  or2  I086_991(w_086_991, w_005_206, w_070_182);
  and2 I086_1093(w_086_1093, w_066_537, w_007_957);
  or2  I086_1118(w_086_1118, w_053_085, w_002_076);
  or2  I086_1168(w_086_1168, w_024_880, w_073_064);
  nand2 I086_1257(w_086_1257, w_011_166, w_026_058);
  nand2 I086_1269(w_086_1269, w_037_219, w_073_018);
  not1 I086_1316(w_086_1316, w_012_307);
  or2  I086_1430(w_086_1430, w_050_354, w_078_884);
  or2  I086_1493(w_086_1493, w_048_598, w_012_573);
  not1 I086_1567(w_086_1567, w_051_252);
  nand2 I086_1569(w_086_1569, w_079_015, w_064_1047);
  or2  I086_1575(w_086_1575, w_042_054, w_022_246);
  nand2 I086_1642(w_086_1642, w_027_469, w_025_570);
  nand2 I087_021(w_087_021, w_059_293, w_048_406);
  nand2 I087_063(w_087_063, w_065_004, w_017_1903);
  and2 I087_110(w_087_110, w_054_579, w_084_142);
  and2 I087_115(w_087_115, w_004_1009, w_074_129);
  or2  I087_146(w_087_146, w_073_096, w_063_388);
  not1 I087_206(w_087_206, w_079_667);
  not1 I087_242(w_087_242, w_032_101);
  not1 I087_289(w_087_289, w_058_1291);
  not1 I087_304(w_087_304, w_042_019);
  and2 I087_347(w_087_347, w_005_864, w_033_370);
  nand2 I087_393(w_087_393, w_010_007, w_036_206);
  not1 I087_462(w_087_462, w_006_130);
  nand2 I087_467(w_087_467, w_084_364, w_032_052);
  not1 I087_524(w_087_524, w_083_006);
  or2  I087_566(w_087_566, w_012_619, w_010_108);
  or2  I087_590(w_087_590, w_068_026, w_053_106);
  or2  I087_607(w_087_607, w_068_031, w_054_300);
  not1 I087_662(w_087_662, w_036_056);
  and2 I087_709(w_087_709, w_082_092, w_086_166);
  and2 I087_772(w_087_772, w_062_556, w_048_383);
  nand2 I087_840(w_087_840, w_054_334, w_073_079);
  nand2 I087_874(w_087_874, w_012_586, w_052_1721);
  and2 I087_971(w_087_971, w_023_1166, w_077_055);
  or2  I087_973(w_087_973, w_074_551, w_069_283);
  not1 I087_978(w_087_978, w_078_995);
  not1 I087_984(w_087_984, w_052_1301);
  nand2 I087_1001(w_087_1001, w_065_005, w_042_009);
  and2 I087_1009(w_087_1009, w_035_1485, w_070_405);
  and2 I087_1021(w_087_1021, w_083_024, w_047_226);
  nand2 I087_1050(w_087_1050, w_040_1178, w_074_274);
  and2 I087_1062(w_087_1062, w_022_294, w_060_096);
  and2 I087_1068(w_087_1068, w_042_001, w_033_307);
  not1 I087_1097(w_087_1097, w_083_002);
  or2  I087_1098(w_087_1098, w_054_592, w_084_158);
  nand2 I087_1104(w_087_1104, w_028_485, w_040_121);
  not1 I087_1123(w_087_1123, w_056_273);
  or2  I087_1173(w_087_1173, w_086_096, w_016_025);
  and2 I087_1211(w_087_1211, w_044_147, w_009_066);
  nand2 I087_1279(w_087_1279, w_056_233, w_066_066);
  nand2 I087_1302(w_087_1302, w_017_307, w_024_065);
  not1 I087_1307(w_087_1307, w_033_058);
  not1 I087_1314(w_087_1314, w_012_107);
  nand2 I087_1366(w_087_1366, w_046_282, w_062_900);
  and2 I087_1383(w_087_1383, w_034_498, w_028_399);
  not1 I087_1426(w_087_1426, w_079_293);
  or2  I087_1451(w_087_1451, w_058_436, w_039_936);
  nand2 I087_1494(w_087_1494, w_052_853, w_009_099);
  or2  I087_1547(w_087_1547, w_013_272, w_073_029);
  nand2 I087_1581(w_087_1581, w_063_255, w_072_038);
  and2 I087_1584(w_087_1584, w_086_569, w_078_285);
  nand2 I087_1603(w_087_1603, w_078_113, w_026_1336);
  nand2 I087_1609(w_087_1609, w_073_016, w_063_171);
  or2  I087_1682(w_087_1682, w_036_1406, w_000_848);
  not1 I088_020(w_088_020, w_071_550);
  or2  I088_030(w_088_030, w_049_971, w_030_067);
  and2 I088_059(w_088_059, w_027_588, w_044_1261);
  not1 I088_067(w_088_067, w_010_403);
  and2 I088_114(w_088_114, w_065_005, w_033_682);
  nand2 I088_118(w_088_118, w_034_161, w_062_527);
  not1 I088_125(w_088_125, w_062_1177);
  not1 I088_139(w_088_139, w_012_621);
  not1 I088_189(w_088_189, w_029_1159);
  not1 I088_210(w_088_210, w_069_039);
  or2  I088_213(w_088_213, w_065_005, w_017_589);
  not1 I088_239(w_088_239, w_058_190);
  and2 I088_258(w_088_258, w_023_040, w_075_179);
  or2  I088_279(w_088_279, w_069_510, w_006_160);
  nand2 I088_286(w_088_286, w_004_1472, w_068_184);
  nand2 I088_291(w_088_291, w_036_764, w_074_155);
  not1 I088_293(w_088_293, w_063_1029);
  not1 I088_326(w_088_326, w_008_119);
  nand2 I088_366(w_088_366, w_071_191, w_011_182);
  and2 I088_421(w_088_421, w_007_568, w_048_668);
  and2 I088_429(w_088_429, w_063_027, w_081_665);
  not1 I088_437(w_088_437, w_007_236);
  nand2 I088_447(w_088_447, w_046_180, w_049_1001);
  nand2 I088_455(w_088_455, w_087_978, w_070_146);
  not1 I088_458(w_088_458, w_034_391);
  or2  I088_467(w_088_467, w_026_660, w_079_526);
  not1 I088_482(w_088_482, w_011_708);
  and2 I088_507(w_088_507, w_001_1362, w_083_002);
  and2 I088_520(w_088_520, w_032_011, w_014_019);
  and2 I088_528(w_088_528, w_041_200, w_085_395);
  nand2 I088_552(w_088_552, w_010_373, w_063_019);
  or2  I088_594(w_088_594, w_019_632, w_064_1140);
  and2 I088_597(w_088_597, w_028_257, w_001_478);
  or2  I088_629(w_088_629, w_081_560, w_074_212);
  or2  I088_642(w_088_642, w_044_954, w_005_487);
  nand2 I088_651(w_088_651, w_065_003, w_007_1103);
  not1 I088_663(w_088_663, w_025_688);
  or2  I088_698(w_088_698, w_019_1021, w_049_543);
  not1 I088_699(w_088_699, w_077_769);
  and2 I088_729(w_088_729, w_012_394, w_000_1909);
  or2  I088_768(w_088_768, w_015_219, w_085_071);
  or2  I088_815(w_088_815, w_083_030, w_018_049);
  and2 I088_900(w_088_900, w_019_858, w_058_498);
  not1 I088_931(w_088_931, w_038_055);
  or2  I088_948(w_088_948, w_067_477, w_005_322);
  not1 I088_1020(w_088_1020, w_066_013);
  nand2 I088_1028(w_088_1028, w_005_675, w_024_1422);
  nand2 I088_1150(w_088_1150, w_060_060, w_061_297);
  or2  I088_1152(w_088_1152, w_080_059, w_033_944);
  and2 I088_1154(w_088_1154, w_071_025, w_000_1356);
  or2  I088_1192(w_088_1192, w_038_473, w_063_1578);
  and2 I088_1214(w_088_1214, w_076_215, w_066_188);
  and2 I088_1239(w_088_1239, w_051_638, w_039_558);
  nand2 I088_1307(w_088_1307, w_034_452, w_014_707);
  nand2 I088_1340(w_088_1340, w_072_076, w_015_081);
  and2 I088_1369(w_088_1369, w_055_567, w_067_676);
  not1 I089_019(w_089_019, w_011_597);
  or2  I089_060(w_089_060, w_020_1147, w_045_1015);
  or2  I089_066(w_089_066, w_088_642, w_002_538);
  not1 I089_067(w_089_067, w_019_908);
  or2  I089_080(w_089_080, w_018_004, w_052_042);
  not1 I089_081(w_089_081, w_067_703);
  or2  I089_101(w_089_101, w_018_216, w_000_1483);
  nand2 I089_107(w_089_107, w_005_080, w_049_541);
  and2 I089_114(w_089_114, w_086_370, w_082_423);
  nand2 I089_127(w_089_127, w_077_873, w_073_065);
  nand2 I089_150(w_089_150, w_085_609, w_038_235);
  and2 I089_155(w_089_155, w_009_108, w_050_1082);
  not1 I089_156(w_089_156, w_018_009);
  and2 I089_179(w_089_179, w_053_004, w_001_487);
  or2  I089_191(w_089_191, w_079_753, w_044_831);
  and2 I089_222(w_089_222, w_056_000, w_081_558);
  not1 I089_282(w_089_282, w_066_859);
  and2 I089_309(w_089_309, w_055_576, w_059_127);
  nand2 I089_328(w_089_328, w_058_367, w_021_189);
  and2 I089_329(w_089_329, w_045_1677, w_061_435);
  not1 I089_340(w_089_340, w_017_1707);
  nand2 I089_360(w_089_360, w_010_097, w_078_632);
  not1 I089_363(w_089_363, w_011_695);
  or2  I089_373(w_089_373, w_085_254, w_005_1429);
  not1 I089_377(w_089_377, w_021_245);
  and2 I089_390(w_089_390, w_057_928, w_007_637);
  not1 I089_402(w_089_402, w_003_029);
  nand2 I089_408(w_089_408, w_066_798, w_005_962);
  or2  I089_419(w_089_419, w_057_1301, w_016_000);
  or2  I089_427(w_089_427, w_075_127, w_031_330);
  and2 I089_438(w_089_438, w_020_979, w_072_059);
  nand2 I089_449(w_089_449, w_067_558, w_063_392);
  nand2 I089_524(w_089_524, w_071_385, w_047_233);
  nand2 I089_547(w_089_547, w_083_005, w_063_175);
  or2  I089_578(w_089_578, w_020_121, w_046_247);
  not1 I089_604(w_089_604, w_087_347);
  nand2 I089_627(w_089_627, w_087_1451, w_041_113);
  not1 I089_629(w_089_629, w_088_1028);
  or2  I089_635(w_089_635, w_077_438, w_064_805);
  and2 I089_647(w_089_647, w_018_128, w_033_1605);
  or2  I089_649(w_089_649, w_036_441, w_040_462);
  not1 I089_679(w_089_679, w_037_1339);
  nand2 I089_688(w_089_688, w_010_317, w_001_661);
  or2  I089_689(w_089_689, w_029_242, w_073_043);
  and2 I089_693(w_089_693, w_062_071, w_032_165);
  nand2 I089_721(w_089_721, w_082_808, w_014_320);
  and2 I089_727(w_089_727, w_014_717, w_081_481);
  nand2 I089_808(w_089_808, w_018_168, w_060_006);
  or2  I089_815(w_089_815, w_080_112, w_054_411);
  and2 I089_832(w_089_832, w_022_067, w_023_780);
  not1 I089_873(w_089_873, w_067_696);
  not1 I089_874(w_089_874, w_024_1244);
  nand2 I089_948(w_089_948, w_087_709, w_045_224);
  not1 I089_951(w_089_951, w_018_230);
  nand2 I089_962(w_089_962, w_051_783, w_037_1210);
  or2  I089_1077(w_089_1077, w_036_953, w_043_073);
  or2  I089_1140(w_089_1140, w_057_233, w_034_273);
  or2  I089_1149(w_089_1149, w_042_122, w_017_804);
  and2 I089_1169(w_089_1169, w_048_918, w_055_053);
  not1 I089_1204(w_089_1204, w_063_618);
  and2 I089_1209(w_089_1209, w_042_063, w_025_458);
  or2  I089_1226(w_089_1226, w_063_287, w_076_118);
  nand2 I089_1242(w_089_1242, w_002_236, w_030_503);
  and2 I089_1252(w_089_1252, w_003_076, w_014_151);
  and2 I089_1258(w_089_1258, w_023_061, w_053_018);
  not1 I089_1266(w_089_1266, w_050_1231);
  not1 I089_1277(w_089_1277, w_042_055);
  nand2 I089_1290(w_089_1290, w_023_1259, w_044_1197);
  and2 I089_1302(w_089_1302, w_083_016, w_013_120);
  not1 I090_015(w_090_015, w_078_747);
  nand2 I090_085(w_090_085, w_016_013, w_009_036);
  or2  I090_095(w_090_095, w_040_1383, w_013_188);
  and2 I090_145(w_090_145, w_079_034, w_089_107);
  and2 I090_146(w_090_146, w_011_129, w_075_187);
  nand2 I090_172(w_090_172, w_016_006, w_030_222);
  nand2 I090_195(w_090_195, w_084_211, w_049_710);
  nand2 I090_196(w_090_196, w_088_520, w_084_315);
  and2 I090_201(w_090_201, w_052_185, w_045_082);
  not1 I090_210(w_090_210, w_081_095);
  or2  I090_223(w_090_223, w_005_131, w_020_961);
  not1 I090_226(w_090_226, w_042_111);
  not1 I090_244(w_090_244, w_083_021);
  and2 I090_250(w_090_250, w_076_327, w_053_110);
  nand2 I090_266(w_090_266, w_065_004, w_067_048);
  nand2 I090_314(w_090_314, w_021_198, w_032_032);
  and2 I090_341(w_090_341, w_064_996, w_053_013);
  or2  I090_363(w_090_363, w_004_1555, w_047_489);
  nand2 I090_384(w_090_384, w_022_324, w_000_055);
  not1 I090_392(w_090_392, w_008_182);
  or2  I090_393(w_090_393, w_020_658, w_037_679);
  and2 I090_413(w_090_413, w_013_099, w_046_020);
  and2 I090_414(w_090_414, w_057_430, w_068_029);
  not1 I090_427(w_090_427, w_006_096);
  and2 I090_457(w_090_457, w_023_1452, w_005_267);
  and2 I090_467(w_090_467, w_085_177, w_043_031);
  nand2 I090_474(w_090_474, w_089_689, w_010_162);
  and2 I090_510(w_090_510, w_005_348, w_007_020);
  not1 I090_553(w_090_553, w_000_701);
  and2 I090_606(w_090_606, w_004_805, w_064_1513);
  not1 I090_615(w_090_615, w_021_163);
  and2 I090_648(w_090_648, w_056_1446, w_053_120);
  or2  I090_663(w_090_663, w_079_145, w_070_423);
  not1 I090_672(w_090_672, w_055_335);
  nand2 I090_696(w_090_696, w_068_190, w_064_1225);
  or2  I090_709(w_090_709, w_079_233, w_030_345);
  and2 I090_716(w_090_716, w_020_431, w_064_227);
  or2  I090_747(w_090_747, w_089_1204, w_032_126);
  nand2 I090_813(w_090_813, w_040_766, w_032_237);
  and2 I090_874(w_090_874, w_038_448, w_059_619);
  and2 I090_875(w_090_875, w_050_1045, w_087_971);
  and2 I090_906(w_090_906, w_004_1562, w_017_707);
  nand2 I090_919(w_090_919, w_015_247, w_071_357);
  nand2 I090_940(w_090_940, w_011_398, w_046_118);
  nand2 I090_984(w_090_984, w_026_1113, w_053_096);
  not1 I090_1067(w_090_1067, w_016_001);
  not1 I090_1125(w_090_1125, w_042_111);
  and2 I090_1139(w_090_1139, w_086_838, w_084_483);
  or2  I090_1154(w_090_1154, w_023_450, w_062_015);
  nand2 I090_1208(w_090_1208, w_058_011, w_055_254);
  not1 I091_003(w_091_003, w_078_349);
  not1 I091_004(w_091_004, w_038_034);
  or2  I091_006(w_091_006, w_077_460, w_004_160);
  and2 I091_008(w_091_008, w_022_234, w_042_142);
  and2 I091_012(w_091_012, w_039_065, w_003_019);
  or2  I091_021(w_091_021, w_066_090, w_015_016);
  not1 I091_022(w_091_022, w_062_271);
  and2 I091_024(w_091_024, w_045_1229, w_027_319);
  or2  I091_025(w_091_025, w_028_639, w_065_004);
  and2 I091_030(w_091_030, w_090_196, w_060_062);
  not1 I091_033(w_091_033, w_070_401);
  not1 I091_039(w_091_039, w_010_322);
  nand2 I091_049(w_091_049, w_006_238, w_022_146);
  or2  I091_052(w_091_052, w_005_140, w_071_018);
  not1 I091_054(w_091_054, w_002_427);
  not1 I091_056(w_091_056, w_065_000);
  or2  I091_059(w_091_059, w_067_532, w_035_894);
  or2  I091_065(w_091_065, w_008_704, w_004_993);
  nand2 I091_069(w_091_069, w_056_217, w_049_087);
  not1 I091_077(w_091_077, w_054_570);
  and2 I091_081(w_091_081, w_082_597, w_043_071);
  or2  I091_088(w_091_088, w_038_198, w_008_065);
  and2 I091_089(w_091_089, w_000_1215, w_052_981);
  or2  I091_090(w_091_090, w_090_553, w_025_032);
  nand2 I091_097(w_091_097, w_079_020, w_061_461);
  nand2 I091_099(w_091_099, w_000_074, w_006_081);
  not1 I091_100(w_091_100, w_086_1257);
  and2 I091_101(w_091_101, w_032_037, w_044_1377);
  not1 I091_105(w_091_105, w_090_648);
  not1 I091_106(w_091_106, w_046_223);
  nand2 I091_107(w_091_107, w_008_112, w_090_146);
  and2 I091_112(w_091_112, w_038_281, w_034_434);
  and2 I091_113(w_091_113, w_080_028, w_035_1102);
  and2 I091_119(w_091_119, w_058_1606, w_062_1289);
  and2 I091_122(w_091_122, w_033_563, w_063_038);
  and2 I091_124(w_091_124, w_010_094, w_049_110);
  not1 I091_125(w_091_125, w_039_721);
  or2  I091_128(w_091_128, w_043_051, w_006_062);
  or2  I091_130(w_091_130, w_066_009, w_084_071);
  not1 I091_132(w_091_132, w_078_1496);
  and2 I091_133(w_091_133, w_068_000, w_057_984);
  not1 I091_140(w_091_140, w_066_896);
  and2 I091_141(w_091_141, w_033_550, w_064_115);
  or2  I091_145(w_091_145, w_050_097, w_003_229);
  and2 I091_150(w_091_150, w_072_040, w_047_057);
  and2 I091_159(w_091_159, w_053_060, w_050_176);
  not1 I091_162(w_091_162, w_000_1486);
  not1 I091_163(w_091_163, w_053_076);
  and2 I091_176(w_091_176, w_061_497, w_087_874);
  or2  I091_177(w_091_177, w_040_854, w_008_431);
  nand2 I091_180(w_091_180, w_000_1654, w_008_368);
  and2 I091_182(w_091_182, w_036_1150, w_014_027);
  and2 I092_004(w_092_004, w_041_111, w_057_240);
  or2  I092_026(w_092_026, w_003_009, w_066_1027);
  nand2 I092_091(w_092_091, w_060_065, w_091_024);
  or2  I092_104(w_092_104, w_085_522, w_024_217);
  and2 I092_107(w_092_107, w_042_089, w_087_206);
  nand2 I092_126(w_092_126, w_052_1110, w_035_1357);
  not1 I092_129(w_092_129, w_002_278);
  nand2 I092_136(w_092_136, w_067_682, w_040_663);
  or2  I092_143(w_092_143, w_015_206, w_037_407);
  nand2 I092_151(w_092_151, w_013_215, w_081_416);
  not1 I092_158(w_092_158, w_090_363);
  not1 I092_163(w_092_163, w_046_140);
  or2  I092_164(w_092_164, w_085_653, w_074_1647);
  nand2 I092_200(w_092_200, w_040_1314, w_039_707);
  nand2 I092_201(w_092_201, w_017_413, w_053_012);
  nand2 I092_204(w_092_204, w_065_002, w_083_029);
  not1 I092_230(w_092_230, w_075_151);
  and2 I092_240(w_092_240, w_079_142, w_080_051);
  or2  I092_281(w_092_281, w_025_059, w_059_497);
  nand2 I092_293(w_092_293, w_003_164, w_038_345);
  nand2 I092_311(w_092_311, w_008_830, w_030_548);
  not1 I092_335(w_092_335, w_003_056);
  nand2 I092_337(w_092_337, w_052_1203, w_012_395);
  not1 I092_367(w_092_367, w_040_297);
  or2  I092_396(w_092_396, w_049_1143, w_019_544);
  or2  I092_426(w_092_426, w_059_503, w_091_159);
  nand2 I092_428(w_092_428, w_044_1077, w_011_715);
  not1 I092_517(w_092_517, w_022_166);
  not1 I092_523(w_092_523, w_062_033);
  not1 I092_526(w_092_526, w_003_031);
  nand2 I092_527(w_092_527, w_055_735, w_019_786);
  not1 I092_540(w_092_540, w_018_218);
  and2 I092_584(w_092_584, w_089_329, w_023_878);
  nand2 I092_591(w_092_591, w_020_176, w_074_1450);
  and2 I092_616(w_092_616, w_048_354, w_052_1598);
  and2 I092_639(w_092_639, w_055_744, w_027_351);
  or2  I092_648(w_092_648, w_082_275, w_032_126);
  or2  I092_651(w_092_651, w_019_416, w_085_388);
  and2 I092_767(w_092_767, w_009_067, w_060_046);
  and2 I092_850(w_092_850, w_068_203, w_035_203);
  not1 I092_881(w_092_881, w_053_073);
  nand2 I092_886(w_092_886, w_030_185, w_013_126);
  nand2 I092_912(w_092_912, w_085_385, w_014_199);
  or2  I092_926(w_092_926, w_064_141, w_045_796);
  or2  I092_943(w_092_943, w_000_488, w_085_200);
  not1 I092_970(w_092_970, w_025_983);
  nand2 I092_1039(w_092_1039, w_037_1520, w_021_020);
  nand2 I092_1156(w_092_1156, w_074_1283, w_040_583);
  not1 I092_1159(w_092_1159, w_021_118);
  nand2 I092_1194(w_092_1194, w_064_264, w_005_1254);
  not1 I093_001(w_093_001, w_032_066);
  and2 I093_004(w_093_004, w_022_341, w_084_314);
  and2 I093_005(w_093_005, w_073_079, w_084_164);
  or2  I093_009(w_093_009, w_003_287, w_004_1699);
  nand2 I093_010(w_093_010, w_045_437, w_023_640);
  nand2 I093_011(w_093_011, w_055_324, w_079_159);
  and2 I093_012(w_093_012, w_056_980, w_078_1347);
  not1 I093_015(w_093_015, w_035_026);
  or2  I093_016(w_093_016, w_035_1471, w_009_005);
  and2 I093_017(w_093_017, w_027_536, w_064_904);
  or2  I093_020(w_093_020, w_037_1357, w_053_050);
  or2  I093_022(w_093_022, w_032_002, w_074_1683);
  nand2 I093_023(w_093_023, w_000_502, w_037_001);
  or2  I093_025(w_093_025, w_039_347, w_074_625);
  or2  I093_034(w_093_034, w_010_311, w_073_087);
  and2 I093_040(w_093_040, w_089_060, w_027_132);
  not1 I093_045(w_093_045, w_056_192);
  and2 I093_048(w_093_048, w_072_077, w_078_538);
  not1 I093_049(w_093_049, w_013_237);
  not1 I093_052(w_093_052, w_068_210);
  or2  I093_054(w_093_054, w_085_204, w_064_102);
  not1 I093_055(w_093_055, w_006_067);
  nand2 I093_059(w_093_059, w_080_082, w_030_625);
  not1 I093_062(w_093_062, w_075_117);
  nand2 I093_063(w_093_063, w_067_280, w_045_398);
  or2  I093_065(w_093_065, w_077_725, w_005_066);
  or2  I093_066(w_093_066, w_083_013, w_076_288);
  and2 I093_068(w_093_068, w_064_1602, w_048_536);
  not1 I093_070(w_093_070, w_065_000);
  or2  I094_002(w_094_002, w_023_1410, w_053_071);
  and2 I094_005(w_094_005, w_050_502, w_052_382);
  or2  I094_006(w_094_006, w_089_832, w_026_817);
  nand2 I094_007(w_094_007, w_080_036, w_034_292);
  not1 I094_008(w_094_008, w_064_293);
  and2 I094_009(w_094_009, w_049_537, w_014_321);
  nand2 I094_011(w_094_011, w_039_1582, w_056_1290);
  not1 I094_012(w_094_012, w_038_144);
  and2 I094_013(w_094_013, w_088_1369, w_054_390);
  nand2 I094_014(w_094_014, w_019_176, w_081_663);
  not1 I094_016(w_094_016, w_037_1422);
  not1 I094_022(w_094_022, w_043_048);
  and2 I094_024(w_094_024, w_014_314, w_084_367);
  or2  I094_036(w_094_036, w_037_1307, w_010_146);
  and2 I094_044(w_094_044, w_037_1278, w_052_947);
  and2 I094_045(w_094_045, w_067_965, w_091_113);
  nand2 I094_046(w_094_046, w_066_971, w_044_176);
  and2 I094_049(w_094_049, w_019_020, w_089_727);
  or2  I094_050(w_094_050, w_036_712, w_037_1054);
  nand2 I094_051(w_094_051, w_089_951, w_015_058);
  and2 I094_053(w_094_053, w_023_969, w_006_226);
  nand2 I094_055(w_094_055, w_077_526, w_003_280);
  not1 I094_056(w_094_056, w_006_334);
  nand2 I094_058(w_094_058, w_059_059, w_051_184);
  not1 I094_061(w_094_061, w_060_038);
  or2  I094_063(w_094_063, w_012_592, w_048_651);
  and2 I094_068(w_094_068, w_023_1140, w_077_310);
  and2 I094_074(w_094_074, w_045_1738, w_016_021);
  and2 I094_076(w_094_076, w_010_346, w_058_608);
  not1 I094_081(w_094_081, w_005_1557);
  and2 I094_083(w_094_083, w_093_045, w_027_182);
  and2 I094_085(w_094_085, w_001_1156, w_017_813);
  not1 I094_087(w_094_087, w_010_048);
  not1 I094_090(w_094_090, w_065_005);
  not1 I094_091(w_094_091, w_052_1248);
  not1 I094_095(w_094_095, w_051_653);
  not1 I094_096(w_094_096, w_073_076);
  not1 I094_098(w_094_098, w_008_064);
  and2 I094_100(w_094_100, w_064_1583, w_082_593);
  and2 I095_020(w_095_020, w_052_711, w_058_220);
  not1 I095_042(w_095_042, w_011_262);
  and2 I095_045(w_095_045, w_081_208, w_007_1574);
  or2  I095_054(w_095_054, w_084_379, w_057_1216);
  nand2 I095_059(w_095_059, w_066_522, w_006_142);
  not1 I095_067(w_095_067, w_036_032);
  not1 I095_068(w_095_068, w_034_363);
  nand2 I095_099(w_095_099, w_048_243, w_080_049);
  nand2 I095_117(w_095_117, w_056_928, w_028_874);
  not1 I095_130(w_095_130, w_072_052);
  not1 I095_148(w_095_148, w_016_030);
  or2  I095_157(w_095_157, w_022_212, w_011_068);
  nand2 I095_167(w_095_167, w_084_267, w_052_715);
  or2  I095_180(w_095_180, w_084_142, w_019_766);
  not1 I095_198(w_095_198, w_006_312);
  not1 I095_233(w_095_233, w_051_198);
  and2 I095_279(w_095_279, w_071_477, w_094_095);
  not1 I095_329(w_095_329, w_094_016);
  nand2 I095_353(w_095_353, w_061_232, w_044_1251);
  nand2 I095_373(w_095_373, w_094_009, w_027_318);
  nand2 I095_387(w_095_387, w_066_016, w_041_152);
  and2 I095_445(w_095_445, w_044_607, w_010_216);
  nand2 I095_468(w_095_468, w_046_138, w_084_418);
  not1 I095_476(w_095_476, w_066_1151);
  or2  I095_479(w_095_479, w_043_101, w_023_822);
  or2  I095_486(w_095_486, w_057_399, w_022_055);
  or2  I095_503(w_095_503, w_076_285, w_050_266);
  and2 I095_506(w_095_506, w_003_290, w_081_040);
  and2 I095_528(w_095_528, w_040_306, w_076_209);
  and2 I095_576(w_095_576, w_023_718, w_028_135);
  and2 I095_580(w_095_580, w_003_084, w_028_118);
  and2 I095_581(w_095_581, w_039_1588, w_074_241);
  or2  I095_639(w_095_639, w_084_123, w_013_186);
  and2 I095_660(w_095_660, w_017_1250, w_011_731);
  and2 I095_675(w_095_675, w_015_108, w_073_099);
  not1 I095_718(w_095_718, w_040_096);
  and2 I095_734(w_095_734, w_093_011, w_090_663);
  not1 I095_736(w_095_736, w_079_030);
  not1 I095_755(w_095_755, w_009_009);
  and2 I095_834(w_095_834, w_061_184, w_043_105);
  and2 I095_836(w_095_836, w_092_527, w_013_280);
  nand2 I095_841(w_095_841, w_086_896, w_057_025);
  or2  I095_845(w_095_845, w_009_015, w_081_669);
  nand2 I095_859(w_095_859, w_026_366, w_011_501);
  not1 I095_884(w_095_884, w_048_551);
  and2 I095_898(w_095_898, w_032_069, w_059_344);
  nand2 I095_900(w_095_900, w_011_735, w_041_081);
  nand2 I096_002(w_096_002, w_044_264, w_017_929);
  nand2 I096_003(w_096_003, w_062_817, w_012_497);
  and2 I096_007(w_096_007, w_072_040, w_047_418);
  or2  I096_012(w_096_012, w_026_190, w_056_1502);
  nand2 I096_027(w_096_027, w_056_196, w_037_111);
  nand2 I096_039(w_096_039, w_067_258, w_089_156);
  not1 I096_042(w_096_042, w_049_786);
  not1 I096_048(w_096_048, w_010_355);
  nand2 I096_054(w_096_054, w_031_1109, w_003_081);
  not1 I096_058(w_096_058, w_003_243);
  not1 I096_073(w_096_073, w_034_599);
  not1 I096_076(w_096_076, w_086_1642);
  or2  I096_085(w_096_085, w_035_029, w_024_114);
  or2  I096_099(w_096_099, w_020_937, w_006_081);
  or2  I096_108(w_096_108, w_049_008, w_079_216);
  and2 I096_109(w_096_109, w_041_074, w_082_341);
  nand2 I096_110(w_096_110, w_078_1352, w_085_418);
  and2 I096_117(w_096_117, w_078_1342, w_074_1335);
  and2 I096_118(w_096_118, w_077_490, w_026_1268);
  or2  I096_134(w_096_134, w_031_465, w_073_083);
  and2 I096_142(w_096_142, w_051_210, w_070_077);
  or2  I096_143(w_096_143, w_059_485, w_037_812);
  not1 I096_144(w_096_144, w_057_1307);
  nand2 I096_147(w_096_147, w_057_058, w_060_098);
  and2 I096_161(w_096_161, w_071_125, w_062_127);
  or2  I096_162(w_096_162, w_039_530, w_063_345);
  nand2 I096_173(w_096_173, w_071_457, w_067_912);
  or2  I096_176(w_096_176, w_011_678, w_091_163);
  or2  I096_183(w_096_183, w_038_065, w_027_059);
  not1 I096_195(w_096_195, w_077_223);
  and2 I096_196(w_096_196, w_015_157, w_060_031);
  not1 I096_201(w_096_201, w_060_028);
  nand2 I096_208(w_096_208, w_034_577, w_047_195);
  and2 I096_218(w_096_218, w_086_176, w_014_205);
  nand2 I096_224(w_096_224, w_078_1036, w_042_060);
  not1 I096_225(w_096_225, w_057_454);
  nand2 I096_227(w_096_227, w_041_180, w_038_397);
  nand2 I096_228(w_096_228, w_036_1139, w_046_070);
  nand2 I097_020(w_097_020, w_033_1635, w_073_030);
  and2 I097_119(w_097_119, w_092_281, w_065_002);
  or2  I097_143(w_097_143, w_013_280, w_045_957);
  not1 I097_239(w_097_239, w_082_426);
  or2  I097_257(w_097_257, w_087_1302, w_033_115);
  not1 I097_266(w_097_266, w_074_1427);
  or2  I097_278(w_097_278, w_020_117, w_096_118);
  not1 I097_279(w_097_279, w_039_025);
  not1 I097_310(w_097_310, w_013_027);
  not1 I097_354(w_097_354, w_046_136);
  or2  I097_370(w_097_370, w_085_058, w_083_007);
  nand2 I097_386(w_097_386, w_021_198, w_061_607);
  or2  I097_390(w_097_390, w_003_051, w_076_140);
  not1 I097_439(w_097_439, w_071_040);
  or2  I097_446(w_097_446, w_003_153, w_088_699);
  and2 I097_456(w_097_456, w_056_745, w_078_854);
  nand2 I097_469(w_097_469, w_009_092, w_044_1176);
  and2 I097_473(w_097_473, w_017_432, w_047_698);
  nand2 I097_489(w_097_489, w_094_061, w_075_118);
  nand2 I097_555(w_097_555, w_085_256, w_061_450);
  not1 I097_556(w_097_556, w_011_290);
  nand2 I097_562(w_097_562, w_062_1180, w_084_055);
  nand2 I097_573(w_097_573, w_015_255, w_015_046);
  and2 I097_579(w_097_579, w_023_622, w_045_209);
  or2  I097_685(w_097_685, w_068_022, w_006_205);
  nand2 I097_704(w_097_704, w_031_111, w_028_420);
  nand2 I097_712(w_097_712, w_089_373, w_080_013);
  nand2 I097_717(w_097_717, w_052_145, w_075_247);
  nand2 I097_718(w_097_718, w_019_130, w_095_859);
  nand2 I097_740(w_097_740, w_038_052, w_008_247);
  nand2 I097_743(w_097_743, w_006_299, w_092_143);
  and2 I097_753(w_097_753, w_091_006, w_086_095);
  not1 I097_761(w_097_761, w_055_157);
  or2  I097_801(w_097_801, w_058_732, w_002_226);
  or2  I097_810(w_097_810, w_080_106, w_040_333);
  nand2 I097_817(w_097_817, w_012_368, w_007_1519);
  or2  I097_882(w_097_882, w_014_070, w_062_571);
  nand2 I097_887(w_097_887, w_089_1149, w_001_982);
  not1 I098_001(w_098_001, w_015_027);
  or2  I098_004(w_098_004, w_012_264, w_027_180);
  not1 I098_010(w_098_010, w_046_258);
  or2  I098_031(w_098_031, w_029_529, w_090_015);
  and2 I098_146(w_098_146, w_050_066, w_078_089);
  not1 I098_197(w_098_197, w_035_139);
  not1 I098_254(w_098_254, w_084_070);
  or2  I098_263(w_098_263, w_077_1114, w_073_021);
  and2 I098_274(w_098_274, w_026_1105, w_011_112);
  not1 I098_276(w_098_276, w_022_266);
  or2  I098_307(w_098_307, w_007_338, w_043_019);
  nand2 I098_333(w_098_333, w_081_077, w_040_1119);
  not1 I098_368(w_098_368, w_097_310);
  and2 I098_370(w_098_370, w_060_056, w_000_1712);
  not1 I098_387(w_098_387, w_058_1033);
  not1 I098_389(w_098_389, w_044_355);
  not1 I098_426(w_098_426, w_043_042);
  and2 I098_432(w_098_432, w_048_416, w_026_007);
  or2  I098_460(w_098_460, w_058_1294, w_009_034);
  and2 I098_494(w_098_494, w_058_1169, w_018_092);
  nand2 I098_498(w_098_498, w_008_589, w_060_040);
  not1 I098_509(w_098_509, w_049_378);
  not1 I098_513(w_098_513, w_071_043);
  nand2 I098_602(w_098_602, w_027_157, w_051_347);
  or2  I098_607(w_098_607, w_014_826, w_002_492);
  nand2 I098_609(w_098_609, w_032_002, w_004_700);
  or2  I098_613(w_098_613, w_056_890, w_036_1210);
  or2  I098_685(w_098_685, w_074_1501, w_017_019);
  or2  I098_698(w_098_698, w_080_110, w_071_235);
  nand2 I098_734(w_098_734, w_002_178, w_070_374);
  not1 I098_740(w_098_740, w_048_405);
  or2  I098_798(w_098_798, w_052_743, w_018_066);
  or2  I098_801(w_098_801, w_034_339, w_060_059);
  and2 I098_803(w_098_803, w_096_007, w_088_467);
  or2  I098_804(w_098_804, w_087_1366, w_007_1455);
  or2  I098_815(w_098_815, w_084_405, w_032_026);
  nand2 I098_836(w_098_836, w_050_052, w_092_367);
  or2  I098_930(w_098_930, w_065_001, w_078_088);
  nand2 I098_977(w_098_977, w_026_216, w_039_1308);
  or2  I098_1010(w_098_1010, w_069_331, w_023_1182);
  or2  I098_1051(w_098_1051, w_021_009, w_094_055);
  not1 I098_1076(w_098_1076, w_045_711);
  or2  I099_036(w_099_036, w_060_032, w_075_061);
  not1 I099_037(w_099_037, w_080_001);
  or2  I099_039(w_099_039, w_003_297, w_004_996);
  nand2 I099_048(w_099_048, w_047_291, w_019_391);
  or2  I099_080(w_099_080, w_097_279, w_012_446);
  nand2 I099_096(w_099_096, w_001_280, w_058_1019);
  and2 I099_136(w_099_136, w_011_005, w_030_424);
  or2  I099_139(w_099_139, w_050_897, w_096_027);
  nand2 I099_140(w_099_140, w_078_1120, w_060_103);
  or2  I099_149(w_099_149, w_034_241, w_088_482);
  not1 I099_161(w_099_161, w_086_160);
  and2 I099_172(w_099_172, w_009_068, w_017_740);
  or2  I099_191(w_099_191, w_043_004, w_055_636);
  not1 I099_211(w_099_211, w_041_021);
  and2 I099_214(w_099_214, w_072_067, w_097_278);
  and2 I099_224(w_099_224, w_007_948, w_032_087);
  and2 I099_282(w_099_282, w_076_211, w_037_675);
  nand2 I099_292(w_099_292, w_076_085, w_070_463);
  nand2 I099_389(w_099_389, w_013_114, w_019_755);
  and2 I099_412(w_099_412, w_089_282, w_019_190);
  and2 I099_429(w_099_429, w_014_517, w_012_500);
  nand2 I099_453(w_099_453, w_087_1581, w_083_014);
  nand2 I099_495(w_099_495, w_022_227, w_076_267);
  nand2 I099_519(w_099_519, w_038_022, w_035_276);
  and2 I099_545(w_099_545, w_000_1522, w_087_1173);
  or2  I099_553(w_099_553, w_017_1860, w_001_242);
  or2  I099_611(w_099_611, w_087_973, w_027_102);
  not1 I099_632(w_099_632, w_042_109);
  not1 I099_677(w_099_677, w_043_035);
  nand2 I099_686(w_099_686, w_078_723, w_064_197);
  and2 I099_691(w_099_691, w_031_744, w_018_064);
  or2  I099_714(w_099_714, w_026_622, w_065_005);
  not1 I099_796(w_099_796, w_077_009);
  not1 I099_816(w_099_816, w_048_827);
  nand2 I099_818(w_099_818, w_047_462, w_084_470);
  and2 I099_837(w_099_837, w_046_087, w_004_810);
  or2  I099_937(w_099_937, w_001_295, w_010_403);
  nand2 I099_994(w_099_994, w_024_098, w_096_227);
  nand2 I099_1076(w_099_1076, w_084_079, w_093_048);
  and2 I099_1080(w_099_1080, w_044_990, w_015_209);
  nand2 I099_1093(w_099_1093, w_037_1000, w_043_095);
  not1 I100_000(w_100_000, w_031_662);
  not1 I100_021(w_100_021, w_095_117);
  or2  I100_082(w_100_082, w_086_291, w_086_1569);
  nand2 I100_147(w_100_147, w_046_180, w_084_013);
  not1 I100_155(w_100_155, w_032_150);
  not1 I100_186(w_100_186, w_033_1205);
  or2  I100_214(w_100_214, w_079_718, w_055_023);
  not1 I100_278(w_100_278, w_065_001);
  and2 I100_298(w_100_298, w_051_1092, w_061_363);
  nand2 I100_323(w_100_323, w_095_042, w_074_215);
  or2  I100_347(w_100_347, w_007_526, w_049_099);
  not1 I100_401(w_100_401, w_088_1152);
  and2 I100_467(w_100_467, w_061_108, w_079_568);
  not1 I100_472(w_100_472, w_064_861);
  and2 I100_494(w_100_494, w_099_611, w_012_041);
  or2  I100_516(w_100_516, w_067_742, w_002_483);
  not1 I100_538(w_100_538, w_062_137);
  or2  I100_550(w_100_550, w_096_224, w_052_432);
  not1 I100_576(w_100_576, w_001_294);
  not1 I100_579(w_100_579, w_033_397);
  nand2 I100_597(w_100_597, w_077_055, w_034_563);
  and2 I100_602(w_100_602, w_062_077, w_072_075);
  or2  I100_610(w_100_610, w_049_454, w_065_001);
  or2  I100_627(w_100_627, w_050_1394, w_034_099);
  nand2 I100_667(w_100_667, w_062_782, w_013_105);
  not1 I100_688(w_100_688, w_002_367);
  nand2 I100_712(w_100_712, w_070_120, w_044_1217);
  and2 I100_770(w_100_770, w_038_263, w_039_198);
  not1 I100_777(w_100_777, w_043_068);
  nand2 I100_900(w_100_900, w_007_245, w_063_1336);
  or2  I100_1069(w_100_1069, w_059_158, w_098_387);
  or2  I100_1090(w_100_1090, w_010_017, w_037_1689);
  or2  I100_1155(w_100_1155, w_066_898, w_058_589);
  or2  I100_1177(w_100_1177, w_085_355, w_049_252);
  not1 I100_1197(w_100_1197, w_069_1618);
  nand2 I100_1259(w_100_1259, w_010_298, w_015_012);
  nand2 I100_1316(w_100_1316, w_078_1469, w_054_578);
  not1 I100_1332(w_100_1332, w_036_1475);
  or2  I100_1363(w_100_1363, w_036_398, w_074_680);
  nand2 I100_1408(w_100_1408, w_029_300, w_066_546);
  nand2 I100_1442(w_100_1442, w_056_1465, w_095_373);
  and2 I100_1550(w_100_1550, w_042_077, w_061_404);
  and2 I100_1567(w_100_1567, w_057_857, w_041_087);
  or2  I100_1601(w_100_1601, w_025_1550, w_005_1102);
  or2  I100_1813(w_100_1813, w_082_515, w_024_1590);
  not1 I101_033(w_101_033, w_035_818);
  or2  I101_079(w_101_079, w_004_1470, w_011_475);
  or2  I101_094(w_101_094, w_078_636, w_095_736);
  or2  I101_120(w_101_120, w_062_362, w_020_1151);
  and2 I101_142(w_101_142, w_056_936, w_073_066);
  nand2 I101_145(w_101_145, w_027_038, w_009_044);
  nand2 I101_154(w_101_154, w_009_049, w_072_051);
  not1 I101_166(w_101_166, w_034_452);
  and2 I101_203(w_101_203, w_036_049, w_041_066);
  nand2 I101_221(w_101_221, w_098_509, w_058_1236);
  and2 I101_227(w_101_227, w_054_401, w_084_379);
  or2  I101_244(w_101_244, w_050_961, w_093_059);
  or2  I101_324(w_101_324, w_098_740, w_057_516);
  not1 I101_354(w_101_354, w_085_593);
  and2 I101_356(w_101_356, w_086_025, w_053_068);
  nand2 I101_367(w_101_367, w_019_614, w_070_035);
  or2  I101_368(w_101_368, w_031_620, w_024_293);
  and2 I101_432(w_101_432, w_096_054, w_040_1304);
  and2 I101_437(w_101_437, w_004_146, w_032_068);
  or2  I101_453(w_101_453, w_053_107, w_029_589);
  and2 I101_496(w_101_496, w_033_999, w_048_317);
  or2  I101_523(w_101_523, w_071_289, w_041_004);
  not1 I101_539(w_101_539, w_034_439);
  nand2 I101_566(w_101_566, w_000_414, w_014_143);
  and2 I101_594(w_101_594, w_059_117, w_042_053);
  or2  I101_615(w_101_615, w_003_111, w_031_750);
  not1 I101_655(w_101_655, w_036_1481);
  or2  I101_661(w_101_661, w_086_044, w_096_117);
  or2  I101_670(w_101_670, w_080_068, w_064_479);
  nand2 I101_672(w_101_672, w_000_762, w_058_533);
  or2  I101_684(w_101_684, w_083_025, w_053_011);
  or2  I101_745(w_101_745, w_078_829, w_040_364);
  not1 I102_010(w_102_010, w_078_1042);
  and2 I102_017(w_102_017, w_002_568, w_069_1675);
  and2 I102_030(w_102_030, w_060_091, w_088_421);
  nand2 I102_072(w_102_072, w_046_020, w_042_100);
  not1 I102_126(w_102_126, w_036_1379);
  and2 I102_130(w_102_130, w_042_025, w_031_091);
  not1 I102_211(w_102_211, w_056_795);
  nand2 I102_294(w_102_294, w_070_432, w_060_019);
  not1 I102_346(w_102_346, w_025_374);
  nand2 I102_363(w_102_363, w_000_739, w_078_019);
  not1 I102_370(w_102_370, w_092_293);
  not1 I102_462(w_102_462, w_005_766);
  nand2 I102_505(w_102_505, w_079_374, w_016_023);
  nand2 I102_507(w_102_507, w_015_103, w_014_093);
  nand2 I102_519(w_102_519, w_050_322, w_053_108);
  nand2 I102_520(w_102_520, w_048_209, w_068_142);
  nand2 I102_594(w_102_594, w_072_024, w_057_1517);
  and2 I102_605(w_102_605, w_020_692, w_031_038);
  nand2 I102_763(w_102_763, w_018_142, w_060_022);
  and2 I102_797(w_102_797, w_089_1252, w_009_047);
  nand2 I102_848(w_102_848, w_014_262, w_058_1721);
  nand2 I102_931(w_102_931, w_079_784, w_009_006);
  nand2 I102_948(w_102_948, w_093_065, w_028_586);
  nand2 I102_1039(w_102_1039, w_068_119, w_056_679);
  and2 I102_1199(w_102_1199, w_016_001, w_029_032);
  not1 I102_1214(w_102_1214, w_060_054);
  nand2 I102_1216(w_102_1216, w_013_235, w_014_640);
  and2 I102_1258(w_102_1260, w_102_1259, w_026_838);
  nand2 I102_1259(w_102_1261, w_058_054, w_102_1260);
  and2 I102_1260(w_102_1262, w_040_724, w_102_1261);
  or2  I102_1261(w_102_1263, w_026_1029, w_102_1262);
  and2 I102_1262(w_102_1264, w_102_1263, w_018_055);
  and2 I102_1263(w_102_1259, w_102_1264, w_102_1278);
  nand2 I102_1264(w_102_1269, w_102_1268, w_045_405);
  nand2 I102_1265(w_102_1270, w_102_1269, w_003_114);
  or2  I102_1266(w_102_1271, w_007_874, w_102_1270);
  and2 I102_1267(w_102_1272, w_076_138, w_102_1271);
  nand2 I102_1268(w_102_1273, w_086_1093, w_102_1272);
  and2 I102_1269(w_102_1274, w_102_1273, w_073_073);
  and2 I102_1270(w_102_1275, w_046_119, w_102_1274);
  not1 I102_1271(w_102_1276, w_102_1275);
  not1 I102_1272(w_102_1268, w_102_1259);
  and2 I102_1273(w_102_1278, w_030_769, w_102_1276);
  nand2 I103_031(w_103_031, w_064_790, w_067_595);
  or2  I103_062(w_103_062, w_021_137, w_016_027);
  not1 I103_064(w_103_064, w_081_539);
  or2  I103_088(w_103_088, w_038_290, w_018_054);
  nand2 I103_098(w_103_098, w_043_084, w_031_762);
  or2  I103_113(w_103_113, w_080_024, w_011_654);
  or2  I103_133(w_103_133, w_009_012, w_061_280);
  not1 I103_146(w_103_146, w_012_412);
  not1 I103_169(w_103_169, w_038_006);
  not1 I103_196(w_103_196, w_021_261);
  and2 I103_232(w_103_232, w_073_008, w_068_194);
  or2  I103_233(w_103_233, w_049_1041, w_091_008);
  or2  I103_237(w_103_237, w_032_163, w_018_145);
  or2  I103_252(w_103_252, w_024_284, w_025_992);
  not1 I103_286(w_103_286, w_026_595);
  nand2 I103_294(w_103_294, w_098_803, w_066_989);
  and2 I103_304(w_103_304, w_038_256, w_052_1220);
  or2  I103_321(w_103_321, w_012_174, w_016_033);
  not1 I103_329(w_103_329, w_012_079);
  nand2 I103_369(w_103_369, w_004_819, w_079_598);
  nand2 I103_375(w_103_375, w_081_162, w_041_107);
  nand2 I103_378(w_103_378, w_067_609, w_092_337);
  not1 I103_445(w_103_445, w_086_812);
  and2 I103_462(w_103_462, w_001_197, w_070_471);
  nand2 I103_523(w_103_523, w_011_814, w_054_042);
  and2 I103_538(w_103_538, w_075_055, w_034_377);
  and2 I103_553(w_103_553, w_007_257, w_066_047);
  and2 I103_554(w_103_554, w_026_360, w_035_1518);
  and2 I103_561(w_103_561, w_039_915, w_096_208);
  not1 I103_590(w_103_590, w_024_1009);
  or2  I103_629(w_103_629, w_017_1802, w_028_566);
  and2 I103_647(w_103_647, w_084_410, w_094_011);
  not1 I103_663(w_103_663, w_093_025);
  or2  I103_692(w_103_692, w_070_079, w_088_326);
  nand2 I103_718(w_103_718, w_072_073, w_057_1414);
  and2 I103_833(w_103_833, w_101_354, w_035_921);
  not1 I103_977(w_103_977, w_005_811);
  not1 I103_994(w_103_994, w_002_046);
  and2 I103_1055(w_103_1055, w_015_176, w_063_722);
  and2 I103_1200(w_103_1200, w_030_368, w_039_272);
  and2 I103_1257(w_103_1257, w_055_423, w_047_675);
  or2  I103_1264(w_103_1264, w_008_408, w_008_312);
  and2 I103_1299(w_103_1299, w_038_221, w_100_597);
  and2 I103_1313(w_103_1313, w_019_090, w_014_093);
  or2  I103_1337(w_103_1337, w_040_848, w_000_042);
  and2 I103_1375(w_103_1375, w_003_125, w_091_125);
  and2 I103_1398(w_103_1398, w_024_177, w_020_219);
  and2 I103_1422(w_103_1422, w_064_156, w_085_111);
  nand2 I104_128(w_104_128, w_073_067, w_052_465);
  or2  I104_176(w_104_176, w_031_333, w_014_208);
  and2 I104_202(w_104_202, w_042_104, w_005_1129);
  or2  I104_233(w_104_233, w_066_1009, w_043_102);
  or2  I104_385(w_104_385, w_085_607, w_023_533);
  nand2 I104_430(w_104_430, w_092_230, w_060_003);
  nand2 I104_529(w_104_529, w_030_444, w_057_1600);
  or2  I104_613(w_104_613, w_057_1605, w_085_108);
  and2 I104_634(w_104_634, w_094_098, w_089_721);
  and2 I104_635(w_104_635, w_024_1498, w_092_163);
  not1 I104_663(w_104_663, w_056_1342);
  and2 I104_684(w_104_684, w_086_119, w_047_577);
  and2 I104_695(w_104_695, w_050_217, w_020_981);
  not1 I104_723(w_104_723, w_051_265);
  not1 I104_759(w_104_759, w_003_288);
  and2 I104_773(w_104_773, w_002_584, w_008_686);
  nand2 I104_776(w_104_776, w_035_1484, w_039_1407);
  not1 I104_784(w_104_784, w_087_1682);
  nand2 I104_800(w_104_800, w_015_163, w_054_003);
  not1 I104_813(w_104_813, w_009_013);
  not1 I104_938(w_104_938, w_063_909);
  not1 I104_1006(w_104_1006, w_069_072);
  and2 I104_1022(w_104_1022, w_094_045, w_040_1263);
  not1 I104_1031(w_104_1031, w_034_354);
  or2  I104_1049(w_104_1049, w_008_543, w_002_343);
  nand2 I104_1173(w_104_1173, w_101_203, w_096_144);
  not1 I104_1248(w_104_1248, w_078_218);
  or2  I104_1263(w_104_1263, w_059_284, w_103_098);
  not1 I104_1410(w_104_1410, w_008_266);
  nand2 I104_1424(w_104_1424, w_095_675, w_009_065);
  nand2 I104_1546(w_104_1546, w_041_025, w_101_684);
  and2 I104_1580(w_104_1580, w_009_014, w_006_064);
  and2 I104_1581(w_104_1581, w_034_369, w_023_1026);
  or2  I104_1647(w_104_1647, w_081_647, w_011_035);
  not1 I104_1651(w_104_1651, w_049_584);
  or2  I104_1694(w_104_1694, w_097_143, w_035_446);
  and2 I104_1704(w_104_1704, w_056_929, w_025_783);
  nand2 I104_1763(w_104_1763, w_094_081, w_094_076);
  nand2 I104_1768(w_104_1768, w_001_639, w_094_036);
  or2  I105_000(w_105_000, w_066_1040, w_046_193);
  nand2 I105_012(w_105_012, w_086_301, w_058_1145);
  or2  I105_043(w_105_043, w_064_1161, w_053_076);
  or2  I105_048(w_105_048, w_058_1412, w_005_1297);
  nand2 I105_063(w_105_063, w_079_819, w_064_1135);
  or2  I105_074(w_105_074, w_082_409, w_087_984);
  and2 I105_090(w_105_090, w_077_174, w_022_316);
  not1 I105_117(w_105_117, w_092_651);
  or2  I105_123(w_105_123, w_103_252, w_085_201);
  and2 I105_126(w_105_126, w_043_093, w_089_627);
  not1 I105_146(w_105_146, w_064_1058);
  and2 I105_297(w_105_297, w_014_086, w_089_1242);
  or2  I105_330(w_105_330, w_029_040, w_078_1155);
  or2  I105_442(w_105_442, w_097_573, w_085_314);
  nand2 I105_458(w_105_458, w_026_258, w_028_704);
  not1 I105_476(w_105_476, w_037_1177);
  nand2 I105_507(w_105_507, w_021_084, w_035_938);
  nand2 I105_552(w_105_552, w_030_767, w_022_075);
  or2  I105_635(w_105_635, w_077_153, w_034_575);
  nand2 I105_636(w_105_636, w_076_119, w_039_599);
  or2  I105_671(w_105_671, w_011_429, w_019_128);
  and2 I105_740(w_105_740, w_036_379, w_061_076);
  and2 I105_819(w_105_819, w_049_076, w_066_722);
  or2  I105_872(w_105_872, w_050_380, w_058_360);
  or2  I105_875(w_105_875, w_085_571, w_019_893);
  or2  I105_956(w_105_956, w_048_446, w_104_634);
  not1 I105_957(w_105_957, w_044_618);
  or2  I105_1029(w_105_1029, w_099_149, w_052_503);
  and2 I105_1042(w_105_1042, w_067_665, w_078_287);
  not1 I105_1050(w_105_1050, w_026_295);
  and2 I105_1105(w_105_1105, w_024_827, w_017_017);
  nand2 I105_1136(w_105_1136, w_064_954, w_046_228);
  or2  I105_1171(w_105_1171, w_081_059, w_078_205);
  not1 I105_1183(w_105_1183, w_036_1346);
  nand2 I105_1248(w_105_1248, w_010_241, w_104_773);
  and2 I105_1249(w_105_1249, w_087_1068, w_005_1572);
  nand2 I105_1352(w_105_1352, w_052_1247, w_038_387);
  nand2 I105_1403(w_105_1403, w_010_173, w_025_601);
  and2 I105_1459(w_105_1459, w_034_608, w_070_448);
  nand2 I105_1472(w_105_1472, w_068_017, w_104_635);
  not1 I105_1578(w_105_1578, w_079_162);
  and2 I105_1716(w_105_1716, w_039_1162, w_019_709);
  and2 I105_1809(w_105_1809, w_094_046, w_007_1347);
  nand2 I105_1812(w_105_1812, w_080_008, w_035_136);
  nand2 I106_037(w_106_037, w_056_625, w_050_1390);
  or2  I106_043(w_106_043, w_005_1628, w_043_043);
  nand2 I106_078(w_106_078, w_058_1630, w_082_799);
  nand2 I106_089(w_106_089, w_044_393, w_095_468);
  and2 I106_090(w_106_090, w_021_107, w_075_005);
  and2 I106_096(w_106_096, w_076_169, w_020_106);
  nand2 I106_148(w_106_148, w_014_609, w_057_228);
  nand2 I106_158(w_106_158, w_001_831, w_028_325);
  and2 I106_172(w_106_172, w_077_034, w_061_274);
  not1 I106_185(w_106_185, w_026_955);
  not1 I106_215(w_106_215, w_058_1220);
  and2 I106_231(w_106_231, w_034_300, w_011_019);
  not1 I106_252(w_106_252, w_091_100);
  nand2 I106_276(w_106_276, w_090_510, w_076_290);
  and2 I106_278(w_106_278, w_094_009, w_007_106);
  nand2 I106_334(w_106_334, w_025_481, w_095_581);
  not1 I106_336(w_106_336, w_031_492);
  nand2 I106_347(w_106_347, w_055_389, w_015_064);
  nand2 I106_355(w_106_355, w_022_224, w_067_200);
  or2  I106_356(w_106_356, w_082_382, w_049_571);
  not1 I106_363(w_106_363, w_008_119);
  or2  I106_370(w_106_370, w_053_091, w_090_1154);
  not1 I106_380(w_106_380, w_024_986);
  not1 I106_424(w_106_424, w_069_1729);
  not1 I106_471(w_106_471, w_020_293);
  not1 I106_479(w_106_479, w_077_702);
  nand2 I106_520(w_106_520, w_043_026, w_036_596);
  or2  I106_524(w_106_524, w_074_1077, w_095_045);
  or2  I106_533(w_106_533, w_094_063, w_001_1573);
  and2 I106_585(w_106_585, w_075_264, w_103_561);
  not1 I106_677(w_106_677, w_100_1363);
  not1 I106_716(w_106_716, w_052_667);
  or2  I106_720(w_106_720, w_026_1366, w_020_752);
  nand2 I106_722(w_106_722, w_021_129, w_074_1470);
  and2 I106_753(w_106_753, w_040_220, w_012_139);
  or2  I106_764(w_106_764, w_091_112, w_035_263);
  nand2 I106_848(w_106_848, w_043_015, w_036_1217);
  and2 I106_854(w_106_854, w_103_1055, w_071_151);
  nand2 I106_902(w_106_902, w_080_096, w_041_180);
  nand2 I106_1034(w_106_1034, w_061_322, w_048_053);
  nand2 I106_1069(w_106_1069, w_074_059, w_045_1349);
  nand2 I106_1199(w_106_1199, w_097_257, w_016_005);
  not1 I106_1235(w_106_1235, w_015_138);
  nand2 I106_1249(w_106_1249, w_092_523, w_019_482);
  not1 I106_1269(w_106_1269, w_089_948);
  nand2 I106_1377(w_106_1377, w_053_016, w_104_1410);
  not1 I107_000(w_107_000, w_079_640);
  and2 I107_007(w_107_007, w_070_177, w_074_167);
  or2  I107_055(w_107_055, w_033_478, w_080_040);
  or2  I107_188(w_107_188, w_076_210, w_083_014);
  and2 I107_211(w_107_211, w_001_845, w_078_937);
  not1 I107_272(w_107_272, w_075_000);
  and2 I107_282(w_107_282, w_032_146, w_045_588);
  not1 I107_286(w_107_286, w_030_253);
  and2 I107_296(w_107_296, w_084_366, w_095_884);
  and2 I107_308(w_107_308, w_058_203, w_075_074);
  or2  I107_332(w_107_332, w_066_738, w_014_079);
  nand2 I107_364(w_107_364, w_089_150, w_021_086);
  not1 I107_398(w_107_398, w_059_445);
  and2 I107_430(w_107_430, w_096_048, w_044_870);
  nand2 I107_432(w_107_432, w_027_587, w_047_415);
  or2  I107_440(w_107_440, w_104_1768, w_106_1034);
  nand2 I107_468(w_107_468, w_037_939, w_039_687);
  nand2 I107_488(w_107_488, w_023_023, w_094_091);
  and2 I107_495(w_107_495, w_018_182, w_000_1603);
  not1 I107_544(w_107_544, w_038_475);
  not1 I107_571(w_107_571, w_026_431);
  nand2 I107_576(w_107_576, w_022_202, w_013_085);
  and2 I107_581(w_107_581, w_052_498, w_049_255);
  nand2 I107_651(w_107_651, w_085_046, w_003_080);
  not1 I107_660(w_107_660, w_064_474);
  nand2 I107_684(w_107_684, w_079_748, w_055_590);
  and2 I107_731(w_107_731, w_056_254, w_003_062);
  or2  I107_821(w_107_821, w_049_521, w_014_299);
  nand2 I107_888(w_107_888, w_106_902, w_010_112);
  nand2 I107_971(w_107_971, w_035_1437, w_073_059);
  and2 I107_995(w_107_995, w_081_086, w_002_151);
  and2 I107_1115(w_107_1115, w_067_655, w_010_087);
  and2 I107_1194(w_107_1194, w_031_100, w_017_205);
  nand2 I107_1322(w_107_1322, w_017_664, w_049_1058);
  not1 I108_007(w_108_007, w_075_144);
  or2  I108_008(w_108_008, w_086_1567, w_051_310);
  and2 I108_009(w_108_009, w_092_1156, w_043_088);
  or2  I108_019(w_108_019, w_082_549, w_064_1012);
  nand2 I108_022(w_108_022, w_091_099, w_044_196);
  and2 I108_054(w_108_054, w_082_688, w_007_233);
  and2 I108_055(w_108_055, w_077_632, w_070_107);
  and2 I108_067(w_108_067, w_065_001, w_050_565);
  and2 I108_076(w_108_076, w_007_1316, w_013_155);
  and2 I108_128(w_108_128, w_046_280, w_105_1472);
  nand2 I108_134(w_108_134, w_076_296, w_011_613);
  and2 I108_149(w_108_149, w_105_507, w_086_203);
  nand2 I108_207(w_108_207, w_023_1431, w_054_355);
  or2  I108_225(w_108_225, w_037_519, w_045_937);
  or2  I108_245(w_108_245, w_048_142, w_042_026);
  and2 I108_251(w_108_251, w_028_000, w_015_166);
  and2 I108_261(w_108_261, w_041_017, w_083_001);
  and2 I108_266(w_108_266, w_099_048, w_005_506);
  or2  I108_277(w_108_277, w_077_903, w_085_418);
  or2  I108_286(w_108_286, w_102_1216, w_024_380);
  not1 I108_309(w_108_309, w_096_173);
  nand2 I108_374(w_108_374, w_057_105, w_063_312);
  or2  I108_381(w_108_381, w_079_048, w_100_1197);
  and2 I108_387(w_108_387, w_019_817, w_000_1396);
  and2 I108_398(w_108_398, w_033_478, w_009_068);
  or2  I108_428(w_108_428, w_002_041, w_083_003);
  or2  I108_467(w_108_467, w_064_607, w_000_1298);
  not1 I108_499(w_108_499, w_060_024);
  or2  I108_500(w_108_500, w_038_392, w_032_201);
  or2  I108_540(w_108_540, w_034_422, w_085_127);
  and2 I108_549(w_108_549, w_031_781, w_010_134);
  not1 I108_591(w_108_591, w_105_1136);
  not1 I108_652(w_108_652, w_103_304);
  and2 I108_673(w_108_673, w_032_244, w_038_049);
  nand2 I108_693(w_108_693, w_016_026, w_096_110);
  and2 I108_705(w_108_705, w_106_356, w_004_102);
  not1 I108_717(w_108_717, w_039_1335);
  nand2 I108_731(w_108_731, w_018_109, w_098_698);
  not1 I108_734(w_108_734, w_041_229);
  or2  I109_030(w_109_030, w_052_061, w_090_341);
  or2  I109_032(w_109_032, w_091_052, w_076_045);
  nand2 I109_039(w_109_039, w_064_1154, w_099_994);
  nand2 I109_046(w_109_046, w_102_030, w_008_538);
  and2 I109_057(w_109_057, w_050_819, w_000_1637);
  and2 I109_073(w_109_073, w_052_1323, w_076_085);
  not1 I109_077(w_109_077, w_060_040);
  nand2 I109_097(w_109_097, w_094_005, w_108_225);
  not1 I109_105(w_109_105, w_030_161);
  or2  I109_143(w_109_143, w_070_045, w_059_597);
  nand2 I109_145(w_109_145, w_104_233, w_074_080);
  or2  I109_162(w_109_162, w_088_118, w_098_333);
  not1 I109_164(w_109_164, w_059_549);
  nand2 I109_167(w_109_167, w_061_232, w_023_834);
  not1 I109_175(w_109_175, w_022_390);
  not1 I109_177(w_109_177, w_048_000);
  not1 I109_180(w_109_180, w_003_212);
  nand2 I109_182(w_109_182, w_090_474, w_006_218);
  or2  I109_184(w_109_184, w_016_037, w_097_489);
  or2  I109_189(w_109_189, w_053_083, w_108_134);
  or2  I109_196(w_109_196, w_085_135, w_105_442);
  not1 I109_206(w_109_206, w_091_024);
  nand2 I109_208(w_109_208, w_094_081, w_082_658);
  not1 I109_222(w_109_222, w_057_034);
  or2  I109_277(w_109_277, w_026_354, w_013_219);
  and2 I109_280(w_109_280, w_012_527, w_071_164);
  not1 I109_296(w_109_296, w_089_1302);
  not1 I109_313(w_109_313, w_064_239);
  nand2 I109_330(w_109_330, w_041_092, w_037_607);
  not1 I109_335(w_109_335, w_093_015);
  nand2 I109_340(w_109_340, w_063_358, w_021_221);
  not1 I109_373(w_109_373, w_025_780);
  and2 I110_026(w_110_026, w_029_113, w_074_1229);
  not1 I110_095(w_110_095, w_032_048);
  and2 I110_168(w_110_168, w_028_209, w_091_077);
  and2 I110_201(w_110_201, w_066_223, w_019_1040);
  and2 I110_216(w_110_216, w_109_105, w_103_321);
  or2  I110_237(w_110_237, w_082_095, w_069_620);
  nand2 I110_254(w_110_254, w_091_039, w_099_816);
  not1 I110_289(w_110_289, w_068_048);
  or2  I110_293(w_110_293, w_075_098, w_091_107);
  or2  I110_297(w_110_297, w_038_015, w_020_830);
  and2 I110_308(w_110_308, w_024_1570, w_090_095);
  nand2 I110_329(w_110_329, w_105_875, w_060_091);
  nand2 I110_340(w_110_340, w_057_1351, w_004_132);
  nand2 I110_430(w_110_430, w_104_202, w_101_661);
  nand2 I110_471(w_110_471, w_055_650, w_025_165);
  not1 I110_529(w_110_529, w_071_293);
  not1 I110_582(w_110_582, w_042_095);
  not1 I110_610(w_110_610, w_080_105);
  or2  I110_625(w_110_625, w_061_644, w_107_272);
  not1 I110_803(w_110_803, w_094_012);
  not1 I110_835(w_110_835, w_093_012);
  and2 I110_857(w_110_857, w_100_347, w_034_621);
  or2  I110_862(w_110_862, w_086_515, w_004_943);
  not1 I110_905(w_110_905, w_021_225);
  or2  I110_914(w_110_914, w_093_054, w_029_638);
  not1 I110_975(w_110_975, w_035_175);
  nand2 I110_981(w_110_981, w_040_593, w_000_1526);
  or2  I110_1010(w_110_1010, w_006_267, w_003_270);
  not1 I110_1241(w_110_1241, w_033_1357);
  nand2 I110_1345(w_110_1345, w_087_1050, w_073_006);
  not1 I110_1372(w_110_1372, w_019_573);
  and2 I110_1446(w_110_1446, w_042_023, w_104_1022);
  or2  I110_1479(w_110_1479, w_055_012, w_047_569);
  nand2 I110_1502(w_110_1502, w_081_468, w_041_157);
  and2 I110_1508(w_110_1508, w_074_496, w_060_069);
  and2 I110_1610(w_110_1612, w_110_1611, w_110_1633);
  and2 I110_1611(w_110_1613, w_110_1612, w_072_010);
  and2 I110_1612(w_110_1614, w_006_208, w_110_1613);
  or2  I110_1613(w_110_1615, w_004_1051, w_110_1614);
  not1 I110_1614(w_110_1616, w_110_1615);
  or2  I110_1615(w_110_1617, w_054_073, w_110_1616);
  and2 I110_1616(w_110_1611, w_095_845, w_110_1617);
  nand2 I110_1617(w_110_1622, w_092_639, w_110_1621);
  or2  I110_1618(w_110_1623, w_110_1622, w_034_460);
  not1 I110_1619(w_110_1624, w_110_1623);
  and2 I110_1620(w_110_1625, w_110_1624, w_067_620);
  and2 I110_1621(w_110_1626, w_003_265, w_110_1625);
  not1 I110_1622(w_110_1627, w_110_1626);
  and2 I110_1623(w_110_1628, w_105_330, w_110_1627);
  nand2 I110_1624(w_110_1629, w_110_1628, w_061_161);
  nand2 I110_1625(w_110_1630, w_110_1629, w_097_562);
  and2 I110_1626(w_110_1631, w_043_050, w_110_1630);
  not1 I110_1627(w_110_1621, w_110_1612);
  and2 I110_1628(w_110_1633, w_043_049, w_110_1631);
  or2  I111_000(w_111_000, w_089_635, w_021_005);
  nand2 I111_029(w_111_029, w_079_134, w_094_087);
  or2  I111_030(w_111_030, w_034_488, w_022_204);
  and2 I111_069(w_111_069, w_078_281, w_093_066);
  and2 I111_080(w_111_080, w_019_512, w_108_076);
  not1 I111_085(w_111_085, w_063_600);
  or2  I111_122(w_111_122, w_066_116, w_069_1744);
  not1 I111_125(w_111_125, w_054_470);
  not1 I111_151(w_111_151, w_093_070);
  not1 I111_153(w_111_153, w_030_154);
  nand2 I111_168(w_111_168, w_020_692, w_070_110);
  nand2 I111_204(w_111_204, w_064_1137, w_032_194);
  nand2 I111_239(w_111_239, w_060_025, w_030_240);
  or2  I111_251(w_111_251, w_100_667, w_038_265);
  not1 I111_256(w_111_256, w_015_257);
  and2 I111_263(w_111_263, w_073_042, w_100_1601);
  and2 I111_264(w_111_264, w_057_660, w_023_1484);
  and2 I111_289(w_111_289, w_027_033, w_010_330);
  not1 I111_292(w_111_292, w_104_695);
  or2  I111_331(w_111_331, w_071_007, w_073_065);
  or2  I111_333(w_111_333, w_084_123, w_099_453);
  nand2 I111_343(w_111_343, w_043_020, w_082_233);
  nand2 I111_352(w_111_352, w_002_040, w_024_617);
  nand2 I111_376(w_111_376, w_034_358, w_038_073);
  not1 I111_383(w_111_383, w_048_652);
  or2  I111_417(w_111_417, w_045_635, w_017_032);
  or2  I111_418(w_111_418, w_039_1600, w_000_1236);
  not1 I111_426(w_111_426, w_036_538);
  nand2 I111_447(w_111_447, w_012_133, w_004_1597);
  not1 I111_482(w_111_482, w_076_338);
  and2 I111_485(w_111_485, w_073_037, w_033_927);
  not1 I111_509(w_111_509, w_003_079);
  and2 I111_604(w_111_604, w_043_040, w_098_613);
  or2  I111_632(w_111_632, w_103_286, w_014_646);
  and2 I111_666(w_111_666, w_034_336, w_038_031);
  not1 I111_679(w_111_679, w_038_155);
  not1 I111_712(w_111_712, w_039_1065);
  or2  I112_022(w_112_022, w_078_103, w_006_208);
  or2  I112_034(w_112_034, w_001_496, w_098_010);
  or2  I112_109(w_112_109, w_040_1195, w_099_837);
  and2 I112_137(w_112_137, w_074_1217, w_087_1009);
  or2  I112_166(w_112_166, w_039_1470, w_099_937);
  nand2 I112_191(w_112_191, w_054_166, w_098_426);
  and2 I112_215(w_112_215, w_009_035, w_060_005);
  or2  I112_254(w_112_254, w_056_492, w_025_1520);
  not1 I112_274(w_112_274, w_051_469);
  and2 I112_279(w_112_279, w_100_494, w_067_237);
  or2  I112_296(w_112_296, w_028_766, w_095_580);
  not1 I112_301(w_112_301, w_048_897);
  and2 I112_350(w_112_350, w_066_714, w_111_030);
  not1 I112_359(w_112_359, w_049_190);
  and2 I112_391(w_112_391, w_025_982, w_009_004);
  not1 I112_416(w_112_416, w_025_1051);
  nand2 I112_465(w_112_465, w_107_364, w_041_254);
  nand2 I112_514(w_112_514, w_041_289, w_092_1159);
  not1 I112_552(w_112_552, w_042_048);
  and2 I112_554(w_112_554, w_008_060, w_085_454);
  or2  I112_596(w_112_596, w_065_005, w_042_130);
  and2 I112_597(w_112_597, w_006_223, w_077_895);
  and2 I112_602(w_112_602, w_105_957, w_045_1066);
  or2  I112_605(w_112_605, w_083_021, w_007_869);
  not1 I112_631(w_112_631, w_055_216);
  nand2 I112_635(w_112_635, w_050_367, w_084_375);
  or2  I112_677(w_112_677, w_051_027, w_043_095);
  and2 I112_707(w_112_707, w_100_1316, w_105_552);
  or2  I112_716(w_112_716, w_012_559, w_083_021);
  not1 I112_756(w_112_756, w_093_009);
  or2  I112_770(w_112_770, w_098_804, w_101_432);
  nand2 I112_804(w_112_804, w_033_574, w_010_027);
  or2  I112_815(w_112_815, w_035_1371, w_003_153);
  and2 I112_831(w_112_831, w_103_369, w_091_105);
  or2  I112_850(w_112_850, w_083_026, w_014_606);
  nand2 I112_865(w_112_865, w_044_107, w_038_160);
  and2 I112_987(w_112_987, w_064_179, w_059_272);
  not1 I113_007(w_113_007, w_109_189);
  nand2 I113_013(w_113_013, w_011_036, w_041_275);
  not1 I113_053(w_113_053, w_095_841);
  not1 I113_093(w_113_093, w_099_136);
  nand2 I113_097(w_113_097, w_025_593, w_016_021);
  nand2 I113_148(w_113_148, w_029_548, w_035_212);
  or2  I113_176(w_113_176, w_053_024, w_095_718);
  or2  I113_293(w_113_293, w_004_476, w_077_709);
  or2  I113_372(w_113_372, w_095_157, w_044_475);
  and2 I113_390(w_113_390, w_063_006, w_029_943);
  and2 I113_432(w_113_432, w_097_753, w_060_067);
  not1 I113_438(w_113_438, w_067_896);
  not1 I113_458(w_113_458, w_046_174);
  not1 I113_464(w_113_464, w_053_106);
  or2  I113_469(w_113_469, w_102_370, w_085_184);
  nand2 I113_526(w_113_526, w_062_962, w_101_745);
  nand2 I113_555(w_113_555, w_040_521, w_105_090);
  and2 I113_575(w_113_575, w_021_006, w_064_252);
  or2  I113_692(w_113_692, w_014_312, w_076_244);
  and2 I113_708(w_113_708, w_047_599, w_075_249);
  nand2 I113_764(w_113_764, w_013_011, w_040_225);
  or2  I113_769(w_113_769, w_030_503, w_009_098);
  or2  I113_771(w_113_771, w_009_065, w_019_369);
  not1 I113_814(w_113_814, w_053_103);
  not1 I113_832(w_113_832, w_072_005);
  or2  I113_869(w_113_869, w_030_266, w_030_250);
  and2 I113_910(w_113_910, w_027_190, w_056_315);
  or2  I113_925(w_113_925, w_091_106, w_020_1215);
  nand2 I113_979(w_113_979, w_078_1688, w_068_083);
  not1 I113_1021(w_113_1021, w_007_741);
  or2  I114_000(w_114_000, w_031_819, w_091_021);
  or2  I114_007(w_114_007, w_098_798, w_001_1022);
  nand2 I114_015(w_114_015, w_099_191, w_010_397);
  nand2 I114_020(w_114_020, w_080_028, w_063_140);
  or2  I114_062(w_114_062, w_056_033, w_009_088);
  nand2 I114_116(w_114_116, w_073_031, w_102_1039);
  and2 I114_126(w_114_126, w_099_519, w_038_367);
  and2 I114_129(w_114_129, w_078_1506, w_048_098);
  and2 I114_161(w_114_161, w_080_021, w_055_005);
  or2  I114_207(w_114_207, w_061_012, w_111_333);
  and2 I114_231(w_114_231, w_095_233, w_036_124);
  or2  I114_252(w_114_252, w_098_836, w_080_090);
  not1 I114_290(w_114_290, w_048_588);
  not1 I114_294(w_114_294, w_112_391);
  not1 I114_302(w_114_302, w_047_532);
  or2  I114_355(w_114_355, w_094_051, w_061_424);
  nand2 I114_435(w_114_435, w_071_442, w_048_783);
  nand2 I114_479(w_114_479, w_085_033, w_000_1489);
  or2  I114_490(w_114_490, w_055_672, w_046_173);
  or2  I114_511(w_114_511, w_018_005, w_050_326);
  or2  I114_541(w_114_541, w_080_109, w_008_635);
  and2 I114_572(w_114_572, w_109_167, w_075_213);
  not1 I114_613(w_114_613, w_111_426);
  or2  I114_627(w_114_627, w_071_048, w_105_872);
  or2  I114_632(w_114_632, w_026_192, w_095_445);
  not1 I114_658(w_114_658, w_052_1341);
  nand2 I114_732(w_114_732, w_099_1093, w_075_105);
  not1 I114_785(w_114_785, w_103_233);
  or2  I114_885(w_114_885, w_057_1249, w_096_201);
  or2  I114_1015(w_114_1015, w_094_002, w_008_039);
  and2 I114_1047(w_114_1047, w_090_427, w_008_044);
  and2 I114_1175(w_114_1175, w_060_011, w_087_467);
  or2  I114_1212(w_114_1212, w_103_1299, w_007_889);
  or2  I114_1247(w_114_1247, w_041_211, w_078_557);
  nand2 I114_1318(w_114_1318, w_038_319, w_060_053);
  and2 I115_014(w_115_014, w_110_216, w_090_392);
  nand2 I115_017(w_115_017, w_028_670, w_017_1370);
  nand2 I115_020(w_115_020, w_027_145, w_046_215);
  not1 I115_066(w_115_066, w_110_340);
  not1 I115_079(w_115_079, w_020_793);
  not1 I115_111(w_115_111, w_083_003);
  not1 I115_112(w_115_112, w_106_424);
  not1 I115_129(w_115_129, w_048_073);
  or2  I115_212(w_115_212, w_082_507, w_059_599);
  and2 I115_286(w_115_286, w_078_252, w_099_691);
  not1 I115_295(w_115_295, w_038_480);
  and2 I115_296(w_115_296, w_114_627, w_064_1377);
  nand2 I115_321(w_115_321, w_110_857, w_109_143);
  or2  I115_333(w_115_333, w_089_419, w_041_146);
  and2 I115_376(w_115_376, w_086_633, w_097_761);
  nand2 I115_388(w_115_388, w_034_189, w_088_059);
  not1 I115_405(w_115_405, w_032_057);
  not1 I115_410(w_115_410, w_106_716);
  and2 I115_413(w_115_413, w_042_003, w_083_023);
  nand2 I115_416(w_115_416, w_106_722, w_021_184);
  not1 I115_420(w_115_420, w_010_018);
  and2 I115_429(w_115_429, w_010_032, w_072_019);
  or2  I115_432(w_115_432, w_035_440, w_074_811);
  or2  I115_434(w_115_434, w_038_068, w_020_886);
  not1 I115_460(w_115_460, w_073_069);
  and2 I115_501(w_115_501, w_035_804, w_108_540);
  or2  I115_508(w_115_508, w_002_192, w_091_119);
  or2  I115_509(w_115_509, w_055_113, w_012_428);
  or2  I115_524(w_115_524, w_000_1380, w_002_447);
  or2  I115_540(w_115_540, w_024_308, w_028_095);
  nand2 I115_559(w_115_559, w_055_306, w_002_302);
  not1 I115_569(w_115_569, w_098_307);
  not1 I115_579(w_115_579, w_075_282);
  and2 I115_598(w_115_598, w_077_1107, w_062_341);
  nand2 I115_603(w_115_603, w_092_886, w_090_085);
  or2  I115_627(w_115_627, w_015_013, w_090_250);
  and2 I116_086(w_116_086, w_059_288, w_026_1415);
  or2  I116_103(w_116_103, w_059_632, w_058_1624);
  and2 I116_115(w_116_115, w_043_005, w_095_067);
  or2  I116_188(w_116_188, w_047_288, w_085_221);
  or2  I116_228(w_116_228, w_065_005, w_066_291);
  or2  I116_359(w_116_359, w_088_125, w_003_096);
  not1 I116_364(w_116_364, w_041_285);
  not1 I116_386(w_116_386, w_055_423);
  or2  I116_390(w_116_390, w_029_1172, w_060_018);
  nand2 I116_395(w_116_395, w_004_488, w_014_663);
  not1 I116_409(w_116_409, w_030_105);
  or2  I116_421(w_116_421, w_050_1397, w_115_112);
  not1 I116_436(w_116_436, w_088_629);
  and2 I116_454(w_116_454, w_051_710, w_087_1211);
  not1 I116_599(w_116_599, w_079_463);
  not1 I116_670(w_116_670, w_048_792);
  not1 I116_730(w_116_730, w_092_026);
  and2 I116_805(w_116_805, w_085_270, w_109_097);
  not1 I116_878(w_116_878, w_027_017);
  not1 I116_901(w_116_901, w_054_432);
  not1 I116_912(w_116_912, w_103_1264);
  nand2 I116_959(w_116_959, w_035_520, w_051_1015);
  not1 I116_1036(w_116_1036, w_032_218);
  nand2 I116_1050(w_116_1050, w_103_113, w_058_199);
  not1 I116_1268(w_116_1268, w_069_368);
  and2 I116_1342(w_116_1342, w_057_137, w_050_041);
  and2 I116_1364(w_116_1364, w_102_211, w_034_584);
  not1 I116_1463(w_116_1463, w_054_308);
  and2 I116_1491(w_116_1491, w_081_430, w_056_1229);
  nand2 I116_1531(w_116_1531, w_060_076, w_047_054);
  or2  I116_1548(w_116_1550, w_116_1574, w_116_1549);
  or2  I116_1549(w_116_1551, w_116_1550, w_060_013);
  and2 I116_1550(w_116_1552, w_009_036, w_116_1551);
  and2 I116_1551(w_116_1553, w_116_1552, w_077_170);
  or2  I116_1552(w_116_1554, w_073_101, w_116_1553);
  and2 I116_1553(w_116_1555, w_059_272, w_116_1554);
  or2  I116_1554(w_116_1556, w_116_1555, w_001_1454);
  nand2 I116_1555(w_116_1557, w_116_1556, w_027_348);
  nand2 I116_1556(w_116_1558, w_116_1557, w_043_059);
  nand2 I116_1557(w_116_1549, w_022_056, w_116_1558);
  or2  I116_1558(w_116_1563, w_116_1562, w_071_531);
  not1 I116_1559(w_116_1564, w_116_1563);
  and2 I116_1560(w_116_1565, w_092_767, w_116_1564);
  not1 I116_1561(w_116_1566, w_116_1565);
  nand2 I116_1562(w_116_1567, w_116_1566, w_095_279);
  nand2 I116_1563(w_116_1568, w_039_1509, w_116_1567);
  not1 I116_1564(w_116_1569, w_116_1568);
  and2 I116_1565(w_116_1570, w_116_1569, w_063_590);
  and2 I116_1566(w_116_1571, w_029_547, w_116_1570);
  nand2 I116_1567(w_116_1572, w_115_559, w_116_1571);
  not1 I116_1568(w_116_1562, w_116_1550);
  and2 I116_1569(w_116_1574, w_039_1457, w_116_1572);
  not1 I117_012(w_117_012, w_053_069);
  nand2 I117_017(w_117_017, w_027_509, w_076_200);
  not1 I117_028(w_117_028, w_098_146);
  not1 I117_052(w_117_052, w_048_134);
  nand2 I117_099(w_117_099, w_043_052, w_008_765);
  not1 I117_142(w_117_142, w_029_151);
  not1 I117_148(w_117_148, w_076_356);
  or2  I117_179(w_117_179, w_077_1084, w_011_098);
  and2 I117_353(w_117_353, w_039_1919, w_017_858);
  or2  I117_365(w_117_365, w_016_011, w_011_775);
  not1 I117_394(w_117_394, w_041_107);
  not1 I117_412(w_117_412, w_023_348);
  and2 I117_428(w_117_428, w_007_839, w_109_030);
  and2 I117_474(w_117_474, w_003_013, w_066_537);
  not1 I117_492(w_117_492, w_079_094);
  or2  I117_498(w_117_498, w_100_688, w_081_249);
  not1 I117_499(w_117_499, w_005_248);
  not1 I117_532(w_117_532, w_102_505);
  and2 I117_539(w_117_539, w_046_266, w_089_340);
  not1 I117_559(w_117_559, w_091_130);
  and2 I117_570(w_117_570, w_020_039, w_083_030);
  or2  I117_589(w_117_589, w_034_016, w_077_589);
  nand2 I117_633(w_117_633, w_058_174, w_064_108);
  nand2 I117_651(w_117_651, w_095_639, w_085_098);
  and2 I117_762(w_117_762, w_089_402, w_012_430);
  and2 I117_767(w_117_767, w_086_176, w_050_052);
  nand2 I117_827(w_117_827, w_061_437, w_024_1098);
  or2  I117_844(w_117_844, w_089_309, w_098_368);
  nand2 I117_872(w_117_872, w_000_808, w_016_020);
  nand2 I117_997(w_117_997, w_087_709, w_114_207);
  nand2 I117_1219(w_117_1219, w_063_1492, w_095_486);
  and2 I117_1471(w_117_1471, w_017_1104, w_045_1231);
  or2  I118_004(w_118_004, w_085_486, w_058_955);
  nand2 I118_125(w_118_125, w_041_188, w_027_481);
  not1 I118_129(w_118_129, w_044_142);
  not1 I118_143(w_118_143, w_025_1317);
  not1 I118_152(w_118_152, w_079_128);
  nand2 I118_222(w_118_222, w_095_068, w_004_1074);
  and2 I118_228(w_118_228, w_100_627, w_045_009);
  not1 I118_232(w_118_232, w_090_875);
  not1 I118_233(w_118_233, w_111_085);
  nand2 I118_264(w_118_264, w_089_815, w_050_994);
  or2  I118_268(w_118_268, w_086_539, w_111_712);
  or2  I118_342(w_118_342, w_019_980, w_063_289);
  not1 I118_360(w_118_360, w_089_449);
  nand2 I118_465(w_118_465, w_076_048, w_054_180);
  nand2 I118_481(w_118_481, w_016_036, w_047_338);
  not1 I118_540(w_118_540, w_075_221);
  and2 I118_650(w_118_650, w_064_999, w_035_772);
  or2  I118_651(w_118_651, w_067_105, w_048_762);
  or2  I118_664(w_118_664, w_023_994, w_031_1054);
  and2 I118_692(w_118_692, w_022_083, w_051_881);
  and2 I118_710(w_118_710, w_062_094, w_005_259);
  nand2 I118_721(w_118_721, w_035_1017, w_017_743);
  or2  I118_784(w_118_784, w_085_373, w_018_139);
  nand2 I118_795(w_118_795, w_077_798, w_071_202);
  not1 I118_921(w_118_921, w_078_093);
  nand2 I118_923(w_118_923, w_105_123, w_068_179);
  and2 I118_945(w_118_945, w_025_1529, w_034_072);
  or2  I118_1006(w_118_1006, w_061_263, w_107_495);
  nand2 I118_1036(w_118_1036, w_109_296, w_085_099);
  or2  I118_1079(w_118_1079, w_044_724, w_094_053);
  nand2 I118_1137(w_118_1137, w_064_775, w_094_049);
  or2  I118_1139(w_118_1139, w_046_195, w_023_1163);
  nand2 I119_026(w_119_026, w_011_586, w_043_001);
  or2  I119_078(w_119_078, w_060_007, w_043_036);
  nand2 I119_276(w_119_276, w_099_1076, w_109_280);
  nand2 I119_341(w_119_341, w_006_321, w_096_142);
  nand2 I119_395(w_119_395, w_058_1027, w_005_036);
  not1 I119_400(w_119_400, w_114_435);
  nand2 I119_410(w_119_410, w_062_097, w_101_227);
  or2  I119_440(w_119_440, w_088_1239, w_016_004);
  or2  I119_455(w_119_455, w_048_881, w_019_629);
  or2  I119_483(w_119_483, w_067_338, w_013_156);
  not1 I119_536(w_119_536, w_107_684);
  not1 I119_587(w_119_587, w_038_136);
  and2 I119_616(w_119_616, w_012_449, w_048_909);
  nand2 I119_642(w_119_642, w_072_074, w_090_1208);
  or2  I119_783(w_119_783, w_050_1293, w_068_211);
  or2  I119_797(w_119_797, w_062_1332, w_049_272);
  and2 I119_798(w_119_798, w_037_1679, w_031_092);
  or2  I119_815(w_119_815, w_082_115, w_114_1247);
  not1 I119_894(w_119_894, w_083_011);
  or2  I119_924(w_119_924, w_015_206, w_075_252);
  nand2 I119_989(w_119_989, w_095_898, w_033_1638);
  nand2 I119_1092(w_119_1092, w_016_030, w_079_411);
  and2 I119_1112(w_119_1112, w_100_214, w_034_582);
  nand2 I119_1202(w_119_1202, w_045_578, w_013_134);
  or2  I119_1223(w_119_1223, w_092_281, w_029_594);
  not1 I119_1278(w_119_1278, w_020_117);
  and2 I119_1282(w_119_1282, w_083_017, w_070_077);
  and2 I119_1318(w_119_1318, w_077_568, w_104_1581);
  and2 I119_1341(w_119_1341, w_038_027, w_066_870);
  or2  I119_1484(w_119_1484, w_091_122, w_115_296);
  or2  I119_1518(w_119_1518, w_024_018, w_006_210);
  not1 I120_000(w_120_000, w_049_488);
  not1 I120_002(w_120_002, w_115_429);
  or2  I120_010(w_120_010, w_033_1307, w_044_199);
  nand2 I120_032(w_120_032, w_011_852, w_043_050);
  or2  I120_035(w_120_035, w_118_1137, w_010_158);
  not1 I120_037(w_120_037, w_007_283);
  and2 I120_041(w_120_041, w_056_1363, w_050_814);
  and2 I120_043(w_120_043, w_112_716, w_068_223);
  and2 I120_047(w_120_047, w_080_095, w_114_015);
  and2 I120_051(w_120_051, w_046_236, w_030_467);
  nand2 I120_057(w_120_057, w_021_117, w_067_872);
  and2 I120_085(w_120_085, w_079_382, w_070_160);
  not1 I120_086(w_120_086, w_108_591);
  and2 I120_094(w_120_094, w_073_061, w_011_515);
  and2 I120_104(w_120_104, w_048_758, w_115_416);
  nand2 I120_109(w_120_109, w_092_104, w_037_1292);
  not1 I120_111(w_120_111, w_114_541);
  or2  I120_116(w_120_116, w_099_139, w_070_114);
  or2  I120_117(w_120_117, w_016_011, w_028_722);
  not1 I120_118(w_120_118, w_029_568);
  or2  I120_127(w_120_127, w_008_011, w_102_1214);
  and2 I120_128(w_120_128, w_106_037, w_056_1269);
  or2  I120_133(w_120_133, w_080_010, w_050_382);
  and2 I120_141(w_120_141, w_116_188, w_040_239);
  and2 I120_152(w_120_152, w_110_1479, w_090_195);
  nand2 I120_156(w_120_156, w_094_016, w_003_012);
  and2 I120_165(w_120_165, w_009_101, w_042_115);
  not1 I120_168(w_120_168, w_041_193);
  nand2 I120_172(w_120_172, w_031_1037, w_107_576);
  not1 I121_053(w_121_053, w_103_538);
  or2  I121_092(w_121_092, w_052_016, w_058_885);
  nand2 I121_102(w_121_102, w_009_053, w_014_080);
  nand2 I121_103(w_121_103, w_083_020, w_065_005);
  not1 I121_114(w_121_114, w_102_605);
  not1 I121_154(w_121_154, w_040_1028);
  or2  I121_202(w_121_202, w_020_041, w_080_118);
  not1 I121_216(w_121_216, w_027_552);
  or2  I121_231(w_121_231, w_033_498, w_006_325);
  nand2 I121_240(w_121_240, w_098_602, w_000_467);
  and2 I121_339(w_121_339, w_069_1620, w_019_721);
  nand2 I121_356(w_121_356, w_015_181, w_002_378);
  or2  I121_390(w_121_390, w_008_809, w_046_168);
  or2  I121_417(w_121_417, w_012_106, w_081_028);
  and2 I121_422(w_121_422, w_060_076, w_023_514);
  nand2 I121_486(w_121_486, w_072_032, w_039_842);
  and2 I121_501(w_121_501, w_108_008, w_042_093);
  nand2 I121_517(w_121_517, w_012_109, w_119_1484);
  or2  I121_524(w_121_524, w_087_662, w_023_906);
  nand2 I121_656(w_121_656, w_110_803, w_048_584);
  not1 I121_697(w_121_697, w_094_022);
  or2  I121_704(w_121_704, w_111_000, w_031_201);
  or2  I121_710(w_121_710, w_057_298, w_030_799);
  nand2 I121_711(w_121_711, w_015_036, w_074_1250);
  and2 I121_723(w_121_723, w_032_098, w_069_866);
  or2  I121_744(w_121_744, w_105_1050, w_060_029);
  nand2 I121_779(w_121_779, w_057_1103, w_112_605);
  and2 I122_002(w_122_002, w_061_663, w_059_289);
  or2  I122_018(w_122_018, w_049_311, w_069_828);
  not1 I122_063(w_122_063, w_097_801);
  nand2 I122_082(w_122_082, w_009_025, w_078_217);
  and2 I122_088(w_122_088, w_113_764, w_065_004);
  or2  I122_098(w_122_098, w_115_286, w_052_1554);
  and2 I122_102(w_122_102, w_034_281, w_083_021);
  nand2 I122_127(w_122_127, w_008_372, w_090_940);
  and2 I122_129(w_122_129, w_087_1314, w_022_338);
  nand2 I122_175(w_122_175, w_112_109, w_051_149);
  not1 I122_177(w_122_177, w_056_876);
  or2  I122_202(w_122_202, w_063_054, w_089_363);
  or2  I122_259(w_122_259, w_010_419, w_009_020);
  not1 I122_274(w_122_274, w_109_196);
  or2  I122_327(w_122_327, w_089_873, w_093_054);
  nand2 I122_331(w_122_331, w_034_323, w_088_1154);
  or2  I122_364(w_122_364, w_025_119, w_026_236);
  and2 I122_390(w_122_390, w_029_243, w_077_1148);
  not1 I122_399(w_122_399, w_007_002);
  not1 I122_410(w_122_410, w_035_815);
  not1 I122_436(w_122_436, w_026_056);
  nand2 I122_478(w_122_478, w_077_314, w_114_007);
  nand2 I122_532(w_122_532, w_100_1332, w_062_1124);
  and2 I122_556(w_122_556, w_063_1337, w_117_012);
  nand2 I122_570(w_122_570, w_102_363, w_022_268);
  or2  I122_572(w_122_572, w_117_570, w_054_352);
  and2 I122_601(w_122_601, w_008_459, w_102_848);
  not1 I122_605(w_122_605, w_024_1393);
  not1 I123_000(w_123_000, w_017_773);
  not1 I123_004(w_123_004, w_011_685);
  and2 I123_063(w_123_063, w_073_003, w_114_062);
  not1 I123_088(w_123_088, w_018_158);
  not1 I123_134(w_123_134, w_091_150);
  not1 I123_182(w_123_182, w_054_007);
  or2  I123_237(w_123_237, w_078_1664, w_072_081);
  or2  I123_334(w_123_334, w_028_557, w_082_466);
  nand2 I123_346(w_123_346, w_049_1111, w_004_1850);
  and2 I123_374(w_123_374, w_001_1013, w_020_354);
  not1 I123_399(w_123_399, w_060_034);
  nand2 I123_400(w_123_400, w_110_582, w_031_052);
  not1 I123_428(w_123_428, w_043_058);
  not1 I123_455(w_123_455, w_075_234);
  nand2 I123_478(w_123_478, w_106_1069, w_068_075);
  or2  I123_494(w_123_494, w_034_420, w_068_140);
  and2 I123_508(w_123_508, w_077_701, w_059_463);
  nand2 I123_518(w_123_518, w_075_241, w_004_515);
  not1 I123_590(w_123_590, w_099_172);
  and2 I123_615(w_123_615, w_097_740, w_034_329);
  not1 I123_616(w_123_616, w_117_872);
  nand2 I123_618(w_123_618, w_074_136, w_046_171);
  or2  I123_627(w_123_627, w_117_633, w_014_145);
  not1 I123_668(w_123_668, w_039_351);
  not1 I123_792(w_123_792, w_108_499);
  nand2 I123_832(w_123_832, w_099_039, w_063_837);
  or2  I123_865(w_123_865, w_098_001, w_053_092);
  or2  I123_970(w_123_970, w_029_277, w_005_296);
  or2  I123_984(w_123_984, w_026_1126, w_108_009);
  or2  I123_990(w_123_990, w_008_547, w_071_406);
  and2 I123_1084(w_123_1084, w_045_1189, w_005_1664);
  nand2 I123_1098(w_123_1098, w_033_1411, w_088_286);
  not1 I123_1121(w_123_1121, w_024_679);
  nand2 I123_1173(w_123_1173, w_113_869, w_077_232);
  nand2 I123_1252(w_123_1252, w_101_145, w_008_084);
  or2  I124_046(w_124_046, w_044_035, w_080_000);
  or2  I124_048(w_124_048, w_037_372, w_015_034);
  or2  I124_061(w_124_061, w_066_640, w_098_930);
  or2  I124_064(w_124_064, w_091_059, w_123_970);
  and2 I124_083(w_124_083, w_046_134, w_020_243);
  nand2 I124_111(w_124_111, w_034_506, w_029_582);
  or2  I124_112(w_124_112, w_037_745, w_022_413);
  or2  I124_135(w_124_135, w_074_1697, w_022_322);
  or2  I124_142(w_124_142, w_051_407, w_096_218);
  and2 I124_152(w_124_152, w_079_104, w_031_575);
  nand2 I124_155(w_124_155, w_009_010, w_089_874);
  and2 I124_165(w_124_165, w_108_277, w_082_260);
  and2 I124_223(w_124_223, w_058_843, w_117_353);
  not1 I124_260(w_124_260, w_046_149);
  and2 I124_274(w_124_274, w_068_243, w_075_217);
  or2  I124_280(w_124_280, w_083_002, w_075_237);
  or2  I124_377(w_124_377, w_101_033, w_016_025);
  not1 I124_381(w_124_381, w_115_432);
  and2 I124_387(w_124_387, w_111_632, w_050_715);
  and2 I124_393(w_124_393, w_098_513, w_048_623);
  or2  I124_457(w_124_457, w_022_298, w_069_1642);
  not1 I124_466(w_124_466, w_054_007);
  and2 I124_488(w_124_488, w_122_274, w_109_177);
  and2 I124_489(w_124_489, w_086_923, w_110_975);
  and2 I124_662(w_124_662, w_047_552, w_088_931);
  and2 I124_740(w_124_740, w_005_954, w_004_1310);
  not1 I125_047(w_125_047, w_084_351);
  and2 I125_095(w_125_095, w_018_024, w_005_252);
  and2 I125_105(w_125_105, w_009_069, w_118_1006);
  nand2 I125_175(w_125_175, w_100_1069, w_103_977);
  and2 I125_221(w_125_221, w_085_490, w_077_023);
  nand2 I125_252(w_125_252, w_064_829, w_122_364);
  or2  I125_354(w_125_354, w_071_295, w_119_783);
  or2  I125_362(w_125_362, w_087_1098, w_027_006);
  and2 I125_394(w_125_394, w_089_679, w_035_1646);
  or2  I125_397(w_125_397, w_015_011, w_016_027);
  and2 I125_448(w_125_448, w_068_022, w_033_1507);
  nand2 I125_526(w_125_526, w_025_1615, w_064_1440);
  nand2 I125_545(w_125_545, w_070_409, w_061_513);
  not1 I125_560(w_125_560, w_042_104);
  and2 I125_683(w_125_683, w_045_082, w_104_784);
  and2 I125_733(w_125_733, w_099_389, w_080_049);
  not1 I125_811(w_125_811, w_121_697);
  or2  I125_840(w_125_840, w_053_053, w_027_513);
  or2  I125_887(w_125_887, w_106_479, w_015_185);
  or2  I125_956(w_125_956, w_004_173, w_075_087);
  and2 I125_981(w_125_981, w_020_366, w_042_028);
  or2  I125_1050(w_125_1050, w_032_108, w_025_1164);
  not1 I125_1055(w_125_1055, w_116_670);
  and2 I125_1126(w_125_1126, w_108_549, w_003_245);
  or2  I125_1201(w_125_1201, w_101_368, w_028_049);
  not1 I125_1361(w_125_1361, w_008_301);
  nand2 I125_1449(w_125_1449, w_004_524, w_073_036);
  or2  I126_001(w_126_001, w_078_1153, w_085_115);
  not1 I126_004(w_126_004, w_081_678);
  nand2 I126_039(w_126_039, w_042_037, w_061_411);
  nand2 I126_083(w_126_083, w_062_186, w_098_607);
  and2 I126_105(w_126_105, w_018_138, w_005_202);
  or2  I126_106(w_126_106, w_113_293, w_057_037);
  or2  I126_111(w_126_111, w_096_228, w_065_002);
  nand2 I126_122(w_126_122, w_114_020, w_062_1003);
  nand2 I126_138(w_126_138, w_109_330, w_035_213);
  nand2 I126_139(w_126_139, w_076_354, w_070_446);
  or2  I126_165(w_126_165, w_069_188, w_029_213);
  nand2 I126_173(w_126_173, w_106_276, w_099_211);
  and2 I126_177(w_126_177, w_008_610, w_097_266);
  not1 I126_181(w_126_181, w_090_813);
  and2 I126_199(w_126_199, w_124_489, w_022_369);
  or2  I126_220(w_126_220, w_026_010, w_045_962);
  nand2 I126_243(w_126_243, w_007_482, w_015_116);
  and2 I126_256(w_126_256, w_123_000, w_085_001);
  or2  I126_270(w_126_270, w_002_544, w_092_428);
  and2 I126_284(w_126_284, w_025_738, w_103_833);
  not1 I126_295(w_126_295, w_107_731);
  or2  I126_305(w_126_305, w_022_309, w_006_009);
  and2 I126_330(w_126_330, w_102_763, w_092_136);
  and2 I126_344(w_126_344, w_063_1501, w_007_1488);
  or2  I126_363(w_126_363, w_000_1057, w_051_868);
  not1 I126_389(w_126_389, w_055_100);
  or2  I126_403(w_126_403, w_098_815, w_041_219);
  and2 I126_420(w_126_420, w_008_025, w_093_066);
  and2 I127_186(w_127_186, w_031_610, w_119_1223);
  nand2 I127_251(w_127_251, w_005_128, w_032_206);
  nand2 I127_298(w_127_298, w_070_376, w_114_129);
  nand2 I127_307(w_127_307, w_021_077, w_080_048);
  nand2 I127_372(w_127_372, w_081_142, w_099_632);
  or2  I127_399(w_127_399, w_091_180, w_061_303);
  or2  I127_426(w_127_426, w_123_618, w_019_062);
  or2  I127_476(w_127_476, w_019_188, w_113_093);
  not1 I127_482(w_127_482, w_094_007);
  and2 I127_516(w_127_516, w_038_412, w_116_436);
  nand2 I127_624(w_127_624, w_049_519, w_062_504);
  not1 I127_697(w_127_697, w_054_204);
  and2 I127_734(w_127_734, w_121_339, w_020_295);
  and2 I127_783(w_127_783, w_074_231, w_092_943);
  or2  I127_802(w_127_802, w_011_552, w_063_975);
  nand2 I127_807(w_127_807, w_104_1763, w_087_772);
  nand2 I127_866(w_127_866, w_045_607, w_090_874);
  or2  I127_889(w_127_889, w_064_795, w_107_007);
  nand2 I127_932(w_127_932, w_117_767, w_115_295);
  and2 I127_1024(w_127_1024, w_091_025, w_070_050);
  nand2 I128_002(w_128_002, w_084_481, w_017_059);
  and2 I128_008(w_128_008, w_044_972, w_006_237);
  or2  I128_012(w_128_012, w_007_1462, w_030_615);
  not1 I128_031(w_128_031, w_095_198);
  not1 I128_033(w_128_033, w_020_652);
  and2 I128_038(w_128_038, w_071_224, w_083_028);
  not1 I128_058(w_128_058, w_066_363);
  not1 I128_061(w_128_061, w_063_183);
  not1 I128_083(w_128_083, w_006_250);
  not1 I128_084(w_128_084, w_099_282);
  nand2 I128_091(w_128_091, w_079_612, w_094_024);
  or2  I128_109(w_128_109, w_071_355, w_121_053);
  nand2 I128_112(w_128_112, w_071_465, w_115_066);
  not1 I128_116(w_128_116, w_094_090);
  not1 I128_133(w_128_133, w_056_1115);
  or2  I128_168(w_128_168, w_119_587, w_044_1344);
  not1 I128_170(w_128_170, w_123_668);
  and2 I128_176(w_128_176, w_032_234, w_114_572);
  not1 I128_191(w_128_191, w_110_1345);
  and2 I128_197(w_128_197, w_110_168, w_042_103);
  and2 I128_207(w_128_207, w_091_056, w_025_420);
  and2 I128_222(w_128_222, w_115_388, w_103_169);
  nand2 I128_242(w_128_242, w_106_355, w_012_022);
  and2 I128_243(w_128_243, w_041_230, w_062_805);
  nand2 I128_246(w_128_246, w_067_758, w_002_064);
  not1 I128_258(w_128_258, w_022_114);
  and2 I128_259(w_128_259, w_022_235, w_081_221);
  not1 I128_264(w_128_264, w_107_1115);
  not1 I129_010(w_129_010, w_010_056);
  or2  I129_041(w_129_041, w_047_235, w_113_692);
  or2  I129_066(w_129_066, w_088_729, w_122_088);
  not1 I129_090(w_129_090, w_091_119);
  or2  I129_245(w_129_245, w_064_1435, w_002_289);
  not1 I129_332(w_129_332, w_047_320);
  and2 I129_368(w_129_368, w_121_779, w_079_395);
  or2  I129_429(w_129_429, w_039_618, w_050_1088);
  and2 I129_518(w_129_518, w_091_049, w_092_584);
  nand2 I129_607(w_129_607, w_016_010, w_090_201);
  or2  I129_608(w_129_608, w_034_649, w_044_147);
  not1 I129_648(w_129_648, w_094_056);
  and2 I129_675(w_129_675, w_094_050, w_059_622);
  or2  I129_681(w_129_681, w_126_083, w_068_197);
  nand2 I129_744(w_129_744, w_022_293, w_072_066);
  or2  I129_747(w_129_747, w_011_876, w_014_613);
  and2 I129_783(w_129_783, w_074_557, w_042_027);
  not1 I129_795(w_129_795, w_053_047);
  and2 I129_808(w_129_808, w_100_1155, w_085_568);
  and2 I129_877(w_129_877, w_013_336, w_113_555);
  or2  I130_000(w_130_000, w_061_506, w_116_409);
  nand2 I130_029(w_130_029, w_019_350, w_068_200);
  and2 I130_035(w_130_035, w_085_660, w_011_474);
  or2  I130_055(w_130_055, w_034_254, w_102_948);
  nand2 I130_110(w_130_110, w_033_970, w_003_164);
  or2  I130_143(w_130_143, w_038_400, w_038_063);
  not1 I130_152(w_130_152, w_010_215);
  and2 I130_195(w_130_195, w_110_289, w_068_036);
  and2 I130_212(w_130_212, w_051_576, w_043_062);
  nand2 I130_221(w_130_221, w_005_1115, w_113_464);
  and2 I130_259(w_130_259, w_032_111, w_037_114);
  nand2 I130_333(w_130_333, w_106_471, w_085_122);
  and2 I130_347(w_130_347, w_076_074, w_107_308);
  and2 I130_499(w_130_499, w_086_1575, w_009_103);
  or2  I130_508(w_130_508, w_028_671, w_023_502);
  or2  I130_562(w_130_562, w_026_691, w_068_203);
  not1 I130_648(w_130_648, w_009_068);
  nand2 I130_696(w_130_696, w_029_233, w_076_094);
  nand2 I130_700(w_130_700, w_120_086, w_004_1161);
  and2 I130_707(w_130_707, w_128_112, w_035_998);
  and2 I130_721(w_130_721, w_114_355, w_058_840);
  or2  I130_977(w_130_977, w_093_068, w_027_043);
  nand2 I131_011(w_131_011, w_003_256, w_074_583);
  not1 I131_031(w_131_031, w_074_1006);
  not1 I131_038(w_131_038, w_072_069);
  and2 I131_070(w_131_070, w_097_685, w_096_002);
  not1 I131_071(w_131_071, w_046_114);
  or2  I131_127(w_131_127, w_033_949, w_035_1546);
  not1 I131_169(w_131_169, w_069_436);
  and2 I131_311(w_131_311, w_036_085, w_130_696);
  nand2 I131_329(w_131_329, w_091_101, w_025_092);
  nand2 I131_345(w_131_345, w_064_1186, w_057_1536);
  nand2 I131_370(w_131_370, w_068_243, w_077_927);
  nand2 I131_374(w_131_374, w_034_140, w_068_029);
  nand2 I131_376(w_131_376, w_088_366, w_046_099);
  not1 I131_405(w_131_405, w_000_1969);
  and2 I131_410(w_131_410, w_007_1378, w_115_212);
  nand2 I131_440(w_131_440, w_050_383, w_113_469);
  not1 I131_538(w_131_538, w_053_092);
  not1 I131_539(w_131_539, w_113_769);
  nand2 I131_562(w_131_562, w_049_554, w_095_180);
  not1 I131_592(w_131_592, w_108_286);
  and2 I131_634(w_131_634, w_085_064, w_085_046);
  or2  I131_766(w_131_766, w_040_314, w_111_679);
  or2  I131_803(w_131_803, w_026_224, w_030_154);
  nand2 I131_847(w_131_847, w_038_233, w_124_048);
  or2  I131_901(w_131_901, w_014_599, w_124_152);
  or2  I131_968(w_131_968, w_060_028, w_002_102);
  nand2 I131_981(w_131_981, w_001_290, w_021_037);
  nand2 I131_1014(w_131_1014, w_022_104, w_120_156);
  not1 I132_001(w_132_001, w_020_135);
  not1 I132_004(w_132_004, w_046_121);
  nand2 I132_007(w_132_007, w_042_040, w_047_107);
  nand2 I132_009(w_132_009, w_018_232, w_039_665);
  and2 I132_011(w_132_011, w_014_154, w_061_535);
  nand2 I132_012(w_132_012, w_105_1105, w_022_401);
  and2 I132_013(w_132_013, w_075_025, w_016_022);
  or2  I132_015(w_132_015, w_029_077, w_092_107);
  not1 I132_017(w_132_017, w_090_709);
  or2  I132_021(w_132_021, w_104_1651, w_114_885);
  not1 I132_025(w_132_025, w_050_435);
  or2  I132_028(w_132_028, w_010_096, w_008_346);
  not1 I132_029(w_132_029, w_079_556);
  or2  I132_031(w_132_031, w_058_1255, w_092_850);
  or2  I132_032(w_132_032, w_011_295, w_098_460);
  and2 I132_033(w_132_033, w_104_1006, w_029_1129);
  not1 I132_034(w_132_034, w_067_639);
  and2 I132_039(w_132_039, w_002_138, w_064_1154);
  or2  I132_042(w_132_042, w_130_143, w_057_369);
  not1 I132_043(w_132_043, w_089_1290);
  not1 I132_046(w_132_046, w_031_983);
  nand2 I132_051(w_132_051, w_122_532, w_088_651);
  not1 I132_055(w_132_055, w_126_295);
  or2  I132_057(w_132_057, w_086_371, w_105_1352);
  and2 I132_063(w_132_063, w_104_1031, w_051_074);
  not1 I132_065(w_132_065, w_043_034);
  nand2 I132_068(w_132_068, w_018_196, w_095_660);
  not1 I132_072(w_132_072, w_031_704);
  nand2 I132_079(w_132_079, w_009_067, w_114_126);
  nand2 I132_085(w_132_085, w_010_370, w_038_155);
  not1 I132_087(w_132_087, w_096_196);
  nand2 I132_089(w_132_089, w_036_071, w_076_128);
  not1 I132_096(w_132_096, w_007_1338);
  not1 I132_104(w_132_104, w_127_307);
  nand2 I133_036(w_133_036, w_031_296, w_132_028);
  and2 I133_042(w_133_042, w_115_420, w_101_539);
  or2  I133_081(w_133_081, w_075_037, w_031_217);
  nand2 I133_138(w_133_138, w_087_393, w_130_721);
  or2  I133_147(w_133_147, w_064_396, w_008_252);
  and2 I133_170(w_133_170, w_075_254, w_018_098);
  and2 I133_214(w_133_214, w_095_353, w_124_280);
  nand2 I133_267(w_133_267, w_020_776, w_036_273);
  not1 I133_293(w_133_293, w_093_040);
  or2  I133_303(w_133_303, w_079_270, w_058_1146);
  and2 I133_320(w_133_320, w_111_168, w_103_647);
  and2 I133_345(w_133_345, w_017_809, w_071_193);
  and2 I133_374(w_133_374, w_132_013, w_110_1372);
  and2 I133_392(w_133_392, w_132_096, w_045_310);
  not1 I133_411(w_133_411, w_054_016);
  nand2 I133_475(w_133_475, w_073_043, w_017_1101);
  nand2 I133_543(w_133_543, w_065_005, w_005_594);
  nand2 I133_656(w_133_656, w_114_732, w_075_266);
  and2 I133_657(w_133_657, w_029_003, w_039_597);
  not1 I133_719(w_133_719, w_021_250);
  not1 I133_737(w_133_737, w_007_1137);
  nand2 I133_739(w_133_739, w_007_729, w_120_118);
  or2  I133_761(w_133_761, w_068_171, w_131_968);
  or2  I133_813(w_133_813, w_061_540, w_000_973);
  nand2 I133_853(w_133_853, w_088_429, w_065_004);
  not1 I133_907(w_133_907, w_125_105);
  or2  I134_006(w_134_006, w_115_413, w_110_430);
  nand2 I134_012(w_134_012, w_028_223, w_068_176);
  not1 I134_019(w_134_019, w_094_006);
  or2  I134_096(w_134_096, w_031_658, w_092_200);
  nand2 I134_097(w_134_097, w_088_1307, w_058_147);
  and2 I134_135(w_134_135, w_004_406, w_053_108);
  and2 I134_150(w_134_150, w_117_498, w_018_012);
  not1 I134_254(w_134_254, w_005_643);
  nand2 I134_295(w_134_295, w_086_055, w_106_278);
  nand2 I134_321(w_134_321, w_130_055, w_025_1341);
  nand2 I134_352(w_134_352, w_072_059, w_114_479);
  and2 I134_375(w_134_375, w_028_116, w_011_361);
  nand2 I134_414(w_134_414, w_056_833, w_073_008);
  not1 I134_430(w_134_430, w_128_258);
  or2  I134_468(w_134_468, w_112_815, w_073_064);
  nand2 I134_477(w_134_477, w_111_509, w_132_087);
  and2 I134_487(w_134_487, w_027_583, w_054_343);
  not1 I134_804(w_134_804, w_071_306);
  nand2 I134_828(w_134_828, w_113_832, w_120_127);
  or2  I134_893(w_134_893, w_045_1102, w_064_1283);
  or2  I134_944(w_134_944, w_066_380, w_089_808);
  not1 I134_1109(w_134_1109, w_078_864);
  or2  I134_1192(w_134_1192, w_062_504, w_088_020);
  nand2 I134_1230(w_134_1230, w_078_353, w_091_090);
  nand2 I135_004(w_135_004, w_069_921, w_104_759);
  or2  I135_018(w_135_018, w_129_368, w_059_429);
  nand2 I135_073(w_135_073, w_063_422, w_132_063);
  not1 I135_078(w_135_078, w_124_155);
  and2 I135_103(w_135_103, w_080_070, w_129_648);
  or2  I135_114(w_135_114, w_045_070, w_121_202);
  not1 I135_145(w_135_145, w_028_087);
  or2  I135_160(w_135_160, w_064_666, w_002_319);
  and2 I135_182(w_135_182, w_109_073, w_066_930);
  not1 I135_221(w_135_221, w_130_347);
  nand2 I135_226(w_135_226, w_081_183, w_133_320);
  or2  I135_258(w_135_258, w_043_023, w_063_597);
  and2 I135_304(w_135_304, w_131_329, w_092_591);
  or2  I135_336(w_135_336, w_049_1303, w_011_328);
  nand2 I135_346(w_135_346, w_099_686, w_052_1573);
  nand2 I135_378(w_135_378, w_010_303, w_023_355);
  or2  I135_385(w_135_385, w_016_013, w_092_912);
  or2  I135_387(w_135_387, w_057_1031, w_027_590);
  and2 I135_459(w_135_459, w_000_160, w_012_266);
  or2  I135_482(w_135_482, w_102_126, w_089_019);
  or2  I135_506(w_135_506, w_038_113, w_052_1340);
  not1 I135_553(w_135_553, w_095_479);
  and2 I135_570(w_135_570, w_075_014, w_123_627);
  nand2 I135_601(w_135_601, w_011_881, w_004_1120);
  not1 I135_606(w_135_606, w_058_701);
  and2 I136_049(w_136_049, w_037_1678, w_014_624);
  not1 I136_080(w_136_080, w_030_470);
  and2 I136_086(w_136_086, w_097_439, w_017_1051);
  nand2 I136_160(w_136_160, w_055_220, w_126_284);
  or2  I136_168(w_136_168, w_116_1050, w_103_252);
  nand2 I136_223(w_136_223, w_088_948, w_038_258);
  and2 I136_321(w_136_321, w_134_135, w_102_072);
  or2  I136_402(w_136_402, w_112_756, w_025_456);
  or2  I136_458(w_136_458, w_047_046, w_122_129);
  and2 I136_501(w_136_501, w_028_149, w_080_067);
  and2 I136_504(w_136_504, w_073_082, w_080_095);
  not1 I136_511(w_136_511, w_101_142);
  not1 I136_629(w_136_629, w_031_292);
  nand2 I136_661(w_136_661, w_079_112, w_080_018);
  or2  I136_665(w_136_665, w_046_123, w_002_293);
  and2 I136_769(w_136_769, w_088_213, w_034_555);
  nand2 I136_806(w_136_806, w_037_1076, w_071_522);
  not1 I136_823(w_136_823, w_107_660);
  nand2 I136_898(w_136_898, w_063_137, w_069_019);
  not1 I137_007(w_137_007, w_097_446);
  and2 I137_012(w_137_012, w_129_808, w_071_274);
  not1 I137_039(w_137_039, w_055_821);
  not1 I137_112(w_137_112, w_058_315);
  nand2 I137_146(w_137_146, w_052_1918, w_099_545);
  nand2 I137_178(w_137_178, w_047_475, w_107_821);
  or2  I137_239(w_137_239, w_118_125, w_108_207);
  not1 I137_276(w_137_276, w_111_485);
  or2  I137_339(w_137_339, w_118_222, w_039_915);
  nand2 I137_344(w_137_344, w_047_329, w_055_148);
  and2 I137_355(w_137_355, w_133_813, w_039_1869);
  or2  I137_379(w_137_379, w_042_076, w_106_148);
  and2 I137_389(w_137_389, w_006_341, w_001_219);
  or2  I137_399(w_137_399, w_124_083, w_043_098);
  and2 I137_417(w_137_417, w_089_114, w_013_035);
  not1 I137_449(w_137_449, w_114_658);
  or2  I137_463(w_137_463, w_068_048, w_056_1460);
  or2  I137_507(w_137_507, w_107_1194, w_122_478);
  nand2 I137_514(w_137_514, w_047_196, w_020_020);
  not1 I137_653(w_137_653, w_101_120);
  and2 I137_735(w_137_735, w_034_416, w_047_570);
  and2 I137_871(w_137_871, w_045_093, w_099_096);
  or2  I137_952(w_137_952, w_003_243, w_125_1449);
  not1 I138_004(w_138_004, w_026_1274);
  or2  I138_005(w_138_005, w_028_172, w_097_239);
  not1 I138_007(w_138_007, w_049_594);
  nand2 I138_008(w_138_008, w_004_201, w_112_191);
  not1 I138_010(w_138_010, w_107_188);
  and2 I138_013(w_138_013, w_097_579, w_083_010);
  and2 I138_017(w_138_017, w_085_302, w_069_681);
  and2 I138_031(w_138_031, w_133_657, w_023_060);
  nand2 I138_040(w_138_040, w_132_072, w_044_030);
  not1 I138_041(w_138_041, w_042_007);
  not1 I138_044(w_138_044, w_006_196);
  or2  I138_049(w_138_049, w_011_037, w_120_109);
  not1 I138_058(w_138_058, w_100_516);
  or2  I138_064(w_138_064, w_057_1562, w_078_236);
  and2 I138_067(w_138_067, w_120_043, w_124_223);
  or2  I138_100(w_138_100, w_106_078, w_081_576);
  and2 I138_101(w_138_101, w_115_434, w_090_906);
  nand2 I138_106(w_138_106, w_023_929, w_001_184);
  or2  I138_109(w_138_109, w_072_006, w_108_149);
  not1 I138_111(w_138_111, w_006_262);
  nand2 I138_132(w_138_132, w_126_111, w_035_217);
  nand2 I138_135(w_138_135, w_039_018, w_075_263);
  and2 I138_142(w_138_142, w_114_613, w_057_177);
  not1 I138_151(w_138_151, w_120_116);
  nand2 I138_160(w_138_160, w_044_1327, w_123_518);
  or2  I138_172(w_138_172, w_058_1187, w_015_184);
  and2 I139_001(w_139_001, w_130_499, w_071_108);
  not1 I139_066(w_139_066, w_071_167);
  or2  I139_069(w_139_069, w_064_1081, w_104_1424);
  nand2 I139_070(w_139_070, w_107_282, w_136_501);
  nand2 I139_076(w_139_076, w_051_702, w_119_341);
  or2  I139_102(w_139_102, w_032_131, w_027_063);
  and2 I139_120(w_139_120, w_006_212, w_062_063);
  and2 I139_129(w_139_129, w_129_010, w_110_1446);
  not1 I139_156(w_139_156, w_077_197);
  nand2 I139_244(w_139_244, w_043_081, w_009_036);
  nand2 I139_283(w_139_283, w_036_297, w_028_251);
  not1 I139_348(w_139_348, w_061_049);
  or2  I139_404(w_139_404, w_125_840, w_035_642);
  nand2 I139_516(w_139_516, w_090_244, w_103_663);
  not1 I139_580(w_139_580, w_119_1112);
  or2  I139_697(w_139_697, w_022_090, w_119_440);
  or2  I139_715(w_139_715, w_085_357, w_053_035);
  nand2 I139_942(w_139_942, w_110_471, w_077_439);
  and2 I139_952(w_139_952, w_075_231, w_102_346);
  and2 I139_1104(w_139_1104, w_086_555, w_022_414);
  nand2 I139_1263(w_139_1263, w_097_704, w_028_430);
  not1 I139_1326(w_139_1326, w_118_232);
  not1 I139_1379(w_139_1379, w_098_1051);
  or2  I139_1455(w_139_1455, w_005_052, w_084_019);
  nand2 I139_1525(w_139_1525, w_105_1578, w_034_314);
  or2  I139_1723(w_139_1723, w_034_376, w_038_255);
  nand2 I139_1735(w_139_1735, w_027_059, w_132_025);
  or2  I140_045(w_140_045, w_018_191, w_063_059);
  nand2 I140_067(w_140_067, w_102_017, w_072_022);
  and2 I140_100(w_140_100, w_015_017, w_020_784);
  and2 I140_212(w_140_212, w_041_246, w_103_088);
  or2  I140_267(w_140_267, w_059_113, w_065_004);
  nand2 I140_376(w_140_376, w_040_183, w_100_538);
  and2 I140_406(w_140_406, w_110_329, w_037_1602);
  or2  I140_442(w_140_442, w_026_1012, w_077_945);
  nand2 I140_483(w_140_483, w_084_012, w_044_1751);
  not1 I140_529(w_140_529, w_131_440);
  and2 I140_548(w_140_548, w_031_861, w_016_022);
  nand2 I140_570(w_140_570, w_070_175, w_021_088);
  nand2 I140_691(w_140_691, w_125_354, w_028_194);
  not1 I140_745(w_140_745, w_036_486);
  or2  I140_799(w_140_799, w_136_160, w_040_019);
  and2 I140_948(w_140_948, w_052_034, w_090_1139);
  nand2 I140_1319(w_140_1319, w_015_013, w_108_673);
  nand2 I140_1423(w_140_1423, w_026_467, w_021_112);
  not1 I140_1554(w_140_1554, w_097_020);
  not1 I140_1596(w_140_1596, w_010_215);
  and2 I141_004(w_141_004, w_108_128, w_100_147);
  nand2 I141_009(w_141_009, w_132_021, w_025_1529);
  not1 I141_024(w_141_024, w_088_507);
  not1 I141_046(w_141_046, w_050_438);
  and2 I141_060(w_141_060, w_083_030, w_050_1057);
  or2  I141_070(w_141_070, w_061_435, w_070_318);
  nand2 I141_073(w_141_073, w_074_295, w_094_074);
  and2 I141_076(w_141_076, w_097_456, w_090_223);
  nand2 I141_077(w_141_077, w_029_300, w_097_718);
  and2 I141_106(w_141_106, w_100_712, w_126_330);
  not1 I141_123(w_141_123, w_106_185);
  nand2 I141_140(w_141_140, w_082_262, w_082_260);
  not1 I141_148(w_141_148, w_100_1259);
  and2 I141_180(w_141_180, w_012_109, w_089_390);
  and2 I141_255(w_141_255, w_023_065, w_126_173);
  and2 I141_261(w_141_261, w_138_067, w_088_768);
  nand2 I141_267(w_141_267, w_006_089, w_086_742);
  nand2 I141_297(w_141_297, w_131_370, w_036_194);
  and2 I141_328(w_141_328, w_105_043, w_083_003);
  or2  I141_336(w_141_336, w_057_1174, w_119_894);
  and2 I141_369(w_141_369, w_051_274, w_000_844);
  not1 I141_495(w_141_495, w_101_094);
  or2  I141_542(w_141_542, w_006_008, w_039_1295);
  and2 I141_591(w_141_591, w_001_1677, w_042_001);
  nand2 I141_606(w_141_606, w_030_648, w_139_952);
  or2  I141_636(w_141_636, w_077_252, w_015_010);
  or2  I141_720(w_141_720, w_059_278, w_027_246);
  not1 I142_022(w_142_022, w_072_019);
  not1 I142_050(w_142_050, w_061_217);
  or2  I142_140(w_142_140, w_023_1043, w_000_1862);
  nand2 I142_170(w_142_170, w_050_610, w_085_602);
  and2 I142_237(w_142_237, w_117_428, w_133_656);
  or2  I142_279(w_142_279, w_031_684, w_061_000);
  or2  I142_340(w_142_340, w_019_474, w_066_909);
  or2  I142_350(w_142_350, w_104_529, w_100_082);
  or2  I142_457(w_142_457, w_096_085, w_068_105);
  nand2 I142_544(w_142_544, w_018_033, w_067_462);
  and2 I142_557(w_142_557, w_061_486, w_046_170);
  nand2 I142_565(w_142_565, w_139_1104, w_060_095);
  not1 I142_644(w_142_644, w_058_625);
  or2  I142_649(w_142_649, w_130_110, w_076_344);
  not1 I142_697(w_142_697, w_045_548);
  nand2 I142_752(w_142_752, w_056_821, w_031_1026);
  or2  I142_776(w_142_776, w_021_013, w_126_199);
  and2 I142_945(w_142_945, w_032_052, w_026_901);
  nand2 I142_1185(w_142_1185, w_079_176, w_004_050);
  nand2 I143_056(w_143_056, w_119_395, w_045_303);
  or2  I143_098(w_143_098, w_134_295, w_110_308);
  or2  I143_103(w_143_103, w_028_414, w_034_061);
  not1 I143_109(w_143_109, w_118_465);
  and2 I143_110(w_143_110, w_128_207, w_056_1534);
  and2 I143_116(w_143_116, w_075_173, w_117_539);
  nand2 I143_323(w_143_323, w_136_504, w_036_1076);
  nand2 I143_328(w_143_328, w_108_019, w_103_294);
  or2  I143_347(w_143_347, w_088_1020, w_103_629);
  or2  I143_363(w_143_363, w_137_653, w_126_305);
  nand2 I143_370(w_143_370, w_120_128, w_135_073);
  and2 I143_404(w_143_404, w_001_732, w_060_018);
  and2 I143_466(w_143_466, w_023_679, w_029_328);
  and2 I143_515(w_143_515, w_014_280, w_134_944);
  not1 I143_753(w_143_753, w_016_014);
  nand2 I143_941(w_143_941, w_004_1615, w_131_374);
  nand2 I143_988(w_143_988, w_106_090, w_068_165);
  not1 I143_1303(w_143_1303, w_062_072);
  or2  I143_1344(w_143_1344, w_027_076, w_072_047);
  nand2 I143_1469(w_143_1469, w_136_049, w_099_292);
  not1 I143_1478(w_143_1478, w_042_132);
  nand2 I143_1529(w_143_1529, w_104_784, w_137_379);
  nand2 I144_014(w_144_014, w_083_003, w_072_003);
  nand2 I144_044(w_144_044, w_039_1835, w_067_746);
  not1 I144_058(w_144_058, w_125_526);
  or2  I144_077(w_144_077, w_000_783, w_064_1392);
  nand2 I144_139(w_144_139, w_014_295, w_099_161);
  not1 I144_147(w_144_147, w_035_1510);
  and2 I144_197(w_144_197, w_011_034, w_000_1197);
  nand2 I144_271(w_144_271, w_007_442, w_043_014);
  or2  I144_274(w_144_274, w_066_156, w_100_602);
  not1 I144_352(w_144_352, w_141_606);
  nand2 I144_511(w_144_511, w_079_018, w_063_292);
  and2 I144_609(w_144_609, w_020_1166, w_132_009);
  or2  I144_688(w_144_688, w_106_231, w_090_696);
  or2  I144_703(w_144_703, w_046_181, w_123_615);
  not1 I144_704(w_144_704, w_079_573);
  and2 I144_726(w_144_726, w_054_596, w_093_010);
  and2 I144_763(w_144_763, w_055_259, w_030_167);
  and2 I144_874(w_144_874, w_045_747, w_134_254);
  nand2 I144_965(w_144_965, w_071_082, w_086_066);
  nand2 I144_993(w_144_993, w_025_082, w_115_014);
  and2 I144_1040(w_144_1040, w_087_1609, w_029_982);
  and2 I144_1102(w_144_1102, w_046_279, w_116_103);
  and2 I144_1115(w_144_1115, w_103_553, w_124_111);
  or2  I144_1212(w_144_1212, w_061_236, w_028_529);
  or2  I144_1226(w_144_1226, w_123_990, w_108_693);
  nand2 I144_1387(w_144_1387, w_001_1613, w_125_1055);
  or2  I144_1570(w_144_1570, w_120_035, w_018_233);
  and2 I145_005(w_145_005, w_139_102, w_031_697);
  not1 I145_006(w_145_006, w_069_021);
  not1 I145_007(w_145_007, w_087_1001);
  or2  I145_009(w_145_009, w_118_784, w_061_409);
  not1 I145_012(w_145_012, w_035_1673);
  nand2 I145_013(w_145_013, w_046_192, w_116_1463);
  or2  I145_015(w_145_015, w_093_022, w_127_426);
  or2  I145_016(w_145_016, w_093_063, w_101_453);
  nand2 I145_017(w_145_017, w_056_1651, w_054_299);
  nand2 I145_020(w_145_020, w_085_134, w_071_007);
  and2 I145_023(w_145_023, w_099_036, w_051_431);
  not1 I145_024(w_145_024, w_135_103);
  or2  I145_027(w_145_027, w_012_445, w_001_1335);
  nand2 I145_032(w_145_032, w_053_024, w_088_458);
  not1 I145_033(w_145_033, w_060_009);
  nand2 I145_034(w_145_034, w_061_201, w_128_168);
  and2 I145_035(w_145_035, w_093_016, w_074_169);
  and2 I145_036(w_145_036, w_144_077, w_022_225);
  not1 I145_037(w_145_037, w_133_081);
  or2  I145_038(w_145_038, w_055_594, w_137_399);
  not1 I145_040(w_145_040, w_143_056);
  not1 I146_007(w_146_007, w_079_078);
  and2 I146_028(w_146_028, w_031_404, w_015_071);
  and2 I146_055(w_146_055, w_006_197, w_022_111);
  not1 I146_057(w_146_057, w_142_565);
  or2  I146_071(w_146_071, w_023_1544, w_114_1318);
  nand2 I146_075(w_146_075, w_075_003, w_090_393);
  not1 I146_115(w_146_115, w_142_279);
  not1 I146_120(w_146_120, w_118_921);
  and2 I146_134(w_146_134, w_112_514, w_020_734);
  and2 I146_191(w_146_191, w_110_237, w_008_567);
  not1 I146_199(w_146_199, w_089_547);
  and2 I146_202(w_146_202, w_129_675, w_131_901);
  and2 I146_220(w_146_220, w_015_080, w_000_695);
  and2 I146_232(w_146_232, w_051_735, w_081_560);
  not1 I146_234(w_146_234, w_131_562);
  not1 I146_260(w_146_260, w_062_1292);
  or2  I146_297(w_146_297, w_056_178, w_049_1243);
  not1 I146_335(w_146_335, w_125_1201);
  and2 I146_366(w_146_366, w_090_716, w_037_670);
  and2 I146_375(w_146_375, w_075_172, w_135_004);
  not1 I146_395(w_146_395, w_058_025);
  or2  I146_401(w_146_401, w_083_017, w_104_1173);
  not1 I146_403(w_146_403, w_054_233);
  nand2 I146_407(w_146_407, w_016_007, w_042_085);
  not1 I146_418(w_146_418, w_054_036);
  and2 I146_424(w_146_424, w_098_609, w_082_649);
  or2  I147_008(w_147_008, w_141_495, w_011_867);
  nand2 I147_030(w_147_030, w_115_017, w_073_076);
  not1 I147_036(w_147_036, w_085_427);
  or2  I147_040(w_147_040, w_052_817, w_030_067);
  nand2 I147_041(w_147_041, w_093_034, w_113_526);
  not1 I147_049(w_147_049, w_076_066);
  and2 I147_053(w_147_053, w_004_108, w_048_236);
  nand2 I147_066(w_147_066, w_033_1277, w_138_106);
  not1 I147_074(w_147_074, w_074_1230);
  or2  I147_076(w_147_076, w_023_071, w_117_844);
  and2 I147_080(w_147_080, w_114_231, w_026_1325);
  or2  I147_093(w_147_093, w_082_155, w_069_1762);
  not1 I147_105(w_147_105, w_016_030);
  and2 I147_126(w_147_126, w_024_262, w_105_458);
  nand2 I147_153(w_147_153, w_145_015, w_060_013);
  and2 I147_156(w_147_156, w_138_172, w_000_801);
  nand2 I147_159(w_147_159, w_103_378, w_041_007);
  not1 I147_176(w_147_176, w_128_259);
  nand2 I147_189(w_147_189, w_063_1297, w_031_134);
  and2 I147_190(w_147_190, w_096_099, w_078_195);
  not1 I147_198(w_147_198, w_107_440);
  or2  I148_120(w_148_120, w_114_290, w_015_104);
  not1 I148_274(w_148_274, w_035_840);
  nand2 I148_490(w_148_490, w_013_024, w_018_006);
  not1 I148_530(w_148_530, w_027_145);
  nand2 I148_715(w_148_715, w_116_1342, w_075_059);
  not1 I148_806(w_148_806, w_001_042);
  and2 I148_903(w_148_903, w_117_412, w_002_280);
  nand2 I148_932(w_148_932, w_054_286, w_021_122);
  and2 I148_1020(w_148_1020, w_132_085, w_008_525);
  or2  I148_1416(w_148_1416, w_041_253, w_123_346);
  or2  I148_1503(w_148_1503, w_123_792, w_052_1304);
  and2 I148_1730(w_148_1730, w_138_135, w_078_835);
  not1 I148_1796(w_148_1796, w_121_154);
  nand2 I148_1819(w_148_1819, w_066_404, w_094_083);
  or2  I148_1863(w_148_1863, w_079_321, w_035_1010);
  not1 I148_1903(w_148_1903, w_046_218);
  not1 I148_1914(w_148_1916, w_148_1915);
  not1 I148_1915(w_148_1917, w_148_1916);
  or2  I148_1916(w_148_1918, w_148_1917, w_041_110);
  nand2 I148_1917(w_148_1919, w_137_417, w_148_1918);
  not1 I148_1918(w_148_1920, w_148_1919);
  or2  I148_1919(w_148_1921, w_148_1920, w_058_1347);
  nand2 I148_1920(w_148_1922, w_148_1921, w_139_1723);
  nand2 I148_1921(w_148_1923, w_075_187, w_148_1922);
  not1 I148_1922(w_148_1924, w_148_1923);
  and2 I148_1923(w_148_1925, w_148_1924, w_041_288);
  and2 I148_1924(w_148_1915, w_110_905, w_148_1925);
  nand2 I149_028(w_149_028, w_139_066, w_024_965);
  not1 I149_076(w_149_076, w_061_121);
  nand2 I149_090(w_149_090, w_062_433, w_147_189);
  nand2 I149_093(w_149_093, w_091_012, w_135_018);
  not1 I149_095(w_149_095, w_075_257);
  or2  I149_218(w_149_218, w_139_1455, w_005_680);
  or2  I149_252(w_149_252, w_063_043, w_043_078);
  or2  I149_309(w_149_309, w_040_632, w_028_473);
  not1 I149_329(w_149_329, w_001_1641);
  nand2 I149_381(w_149_381, w_029_539, w_055_693);
  and2 I149_489(w_149_489, w_115_509, w_103_133);
  not1 I149_580(w_149_580, w_067_603);
  nand2 I149_581(w_149_581, w_064_1474, w_136_086);
  nand2 I149_590(w_149_590, w_137_735, w_064_1509);
  nand2 I149_594(w_149_594, w_077_623, w_080_099);
  and2 I149_805(w_149_805, w_058_266, w_100_1442);
  not1 I149_1027(w_149_1027, w_123_494);
  nand2 I149_1111(w_149_1111, w_053_063, w_090_1125);
  or2  I149_1125(w_149_1125, w_108_387, w_136_223);
  not1 I149_1158(w_149_1158, w_105_636);
  or2  I150_006(w_150_006, w_063_1140, w_087_1584);
  not1 I150_016(w_150_016, w_107_1322);
  not1 I150_106(w_150_106, w_019_058);
  not1 I150_128(w_150_128, w_114_785);
  or2  I150_144(w_150_144, w_010_129, w_114_161);
  and2 I150_229(w_150_229, w_004_1727, w_054_095);
  or2  I150_421(w_150_421, w_057_861, w_075_071);
  not1 I150_493(w_150_493, w_007_001);
  nand2 I150_654(w_150_654, w_101_079, w_120_051);
  and2 I150_715(w_150_715, w_096_076, w_133_036);
  not1 I150_768(w_150_768, w_120_037);
  and2 I150_817(w_150_817, w_126_177, w_125_095);
  nand2 I150_849(w_150_849, w_106_1377, w_010_200);
  nand2 I150_894(w_150_894, w_097_810, w_051_777);
  or2  I150_1118(w_150_1118, w_144_139, w_036_589);
  and2 I150_1283(w_150_1283, w_128_083, w_140_376);
  not1 I150_1395(w_150_1395, w_127_1024);
  nand2 I150_1409(w_150_1409, w_064_586, w_058_1190);
  nand2 I150_1570(w_150_1570, w_146_199, w_132_065);
  nand2 I150_1648(w_150_1648, w_131_592, w_085_274);
  and2 I150_1721(w_150_1721, w_112_416, w_022_058);
  or2  I150_1759(w_150_1759, w_027_498, w_121_656);
  nand2 I150_1761(w_150_1761, w_082_193, w_123_1121);
  not1 I151_097(w_151_097, w_014_390);
  nand2 I151_103(w_151_103, w_110_095, w_132_004);
  not1 I151_165(w_151_165, w_021_235);
  and2 I151_179(w_151_179, w_013_259, w_132_104);
  nand2 I151_190(w_151_190, w_032_057, w_007_817);
  nand2 I151_350(w_151_350, w_123_004, w_061_568);
  not1 I151_370(w_151_370, w_051_783);
  nand2 I151_380(w_151_380, w_149_1111, w_132_063);
  not1 I151_434(w_151_434, w_064_170);
  not1 I151_454(w_151_454, w_019_415);
  and2 I151_553(w_151_553, w_041_114, w_018_236);
  not1 I151_587(w_151_587, w_097_882);
  nand2 I151_595(w_151_595, w_041_181, w_122_390);
  not1 I151_694(w_151_694, w_127_186);
  nand2 I151_765(w_151_765, w_091_004, w_113_458);
  nand2 I151_834(w_151_834, w_084_065, w_026_1048);
  not1 I151_922(w_151_922, w_020_528);
  nand2 I151_1014(w_151_1014, w_001_006, w_052_392);
  not1 I151_1043(w_151_1043, w_107_571);
  not1 I151_1090(w_151_1090, w_060_038);
  or2  I151_1109(w_151_1109, w_058_459, w_091_162);
  nand2 I151_1182(w_151_1182, w_109_164, w_086_652);
  and2 I151_1310(w_151_1310, w_049_1067, w_133_543);
  or2  I151_1378(w_151_1378, w_027_565, w_017_020);
  and2 I152_031(w_152_031, w_111_263, w_083_029);
  or2  I152_039(w_152_039, w_043_052, w_150_654);
  or2  I152_045(w_152_045, w_035_061, w_048_724);
  and2 I152_065(w_152_065, w_089_649, w_094_096);
  and2 I152_081(w_152_081, w_076_010, w_020_193);
  and2 I152_120(w_152_120, w_138_160, w_116_1364);
  or2  I152_142(w_152_142, w_026_949, w_013_215);
  or2  I152_169(w_152_169, w_010_284, w_001_1303);
  not1 I152_176(w_152_176, w_029_042);
  and2 I152_177(w_152_177, w_034_433, w_003_114);
  not1 I152_216(w_152_216, w_042_110);
  nand2 I152_220(w_152_220, w_089_101, w_074_658);
  nand2 I152_249(w_152_249, w_049_282, w_139_283);
  not1 I152_253(w_152_253, w_044_1405);
  or2  I152_345(w_152_345, w_076_155, w_013_098);
  or2  I152_358(w_152_358, w_113_053, w_125_733);
  not1 I152_367(w_152_367, w_123_508);
  nand2 I152_417(w_152_417, w_105_956, w_113_979);
  and2 I152_430(w_152_430, w_137_012, w_111_485);
  or2  I152_510(w_152_510, w_037_1637, w_122_399);
  nand2 I152_511(w_152_511, w_052_461, w_072_053);
  or2  I153_143(w_153_143, w_152_510, w_047_391);
  and2 I153_156(w_153_156, w_115_569, w_003_077);
  and2 I153_162(w_153_162, w_012_650, w_074_1032);
  nand2 I153_233(w_153_233, w_127_298, w_019_637);
  not1 I153_356(w_153_356, w_003_052);
  and2 I153_373(w_153_373, w_076_335, w_143_1303);
  not1 I153_475(w_153_475, w_109_175);
  nand2 I153_496(w_153_496, w_037_1349, w_128_058);
  nand2 I153_505(w_153_505, w_081_578, w_020_1040);
  and2 I153_641(w_153_641, w_114_632, w_010_140);
  not1 I153_728(w_153_728, w_071_529);
  or2  I153_745(w_153_745, w_050_1374, w_091_099);
  and2 I153_814(w_153_814, w_086_267, w_106_363);
  or2  I153_843(w_153_843, w_116_086, w_071_064);
  and2 I153_886(w_153_886, w_081_290, w_073_096);
  and2 I153_1016(w_153_1016, w_145_013, w_033_1104);
  and2 I153_1254(w_153_1254, w_036_1336, w_025_029);
  not1 I153_1324(w_153_1324, w_047_280);
  or2  I154_000(w_154_000, w_140_1554, w_071_012);
  and2 I154_008(w_154_008, w_000_1316, w_033_660);
  or2  I154_013(w_154_013, w_028_243, w_034_521);
  or2  I154_015(w_154_015, w_089_081, w_024_1059);
  and2 I154_051(w_154_051, w_075_001, w_046_105);
  not1 I154_066(w_154_066, w_066_900);
  not1 I154_071(w_154_071, w_064_266);
  or2  I154_073(w_154_073, w_118_664, w_117_474);
  or2  I154_096(w_154_096, w_133_853, w_054_366);
  nand2 I154_098(w_154_098, w_038_183, w_065_003);
  not1 I154_106(w_154_106, w_130_035);
  nand2 I154_112(w_154_112, w_103_1375, w_029_389);
  not1 I154_123(w_154_123, w_130_212);
  or2  I154_124(w_154_124, w_130_029, w_027_556);
  and2 I154_136(w_154_136, w_051_268, w_046_130);
  and2 I154_142(w_154_142, w_129_518, w_115_020);
  nand2 I154_148(w_154_148, w_009_038, w_037_923);
  and2 I154_171(w_154_171, w_041_271, w_003_282);
  and2 I154_181(w_154_181, w_048_406, w_016_010);
  not1 I154_182(w_154_182, w_059_333);
  nand2 I155_006(w_155_006, w_059_509, w_041_062);
  nand2 I155_073(w_155_073, w_128_061, w_018_138);
  and2 I155_074(w_155_074, w_134_1109, w_108_022);
  and2 I155_174(w_155_174, w_050_169, w_141_267);
  not1 I155_207(w_155_207, w_032_210);
  or2  I155_284(w_155_284, w_087_021, w_012_116);
  or2  I155_561(w_155_561, w_088_437, w_080_050);
  nand2 I155_762(w_155_762, w_068_050, w_004_983);
  or2  I155_784(w_155_784, w_050_220, w_045_005);
  nand2 I155_805(w_155_805, w_093_017, w_063_1164);
  nand2 I155_838(w_155_838, w_050_038, w_001_187);
  and2 I155_982(w_155_982, w_059_298, w_153_886);
  nand2 I155_1152(w_155_1152, w_053_007, w_094_046);
  and2 I155_1257(w_155_1257, w_038_192, w_134_321);
  and2 I155_1682(w_155_1682, w_015_021, w_146_424);
  nand2 I156_023(w_156_023, w_106_520, w_132_029);
  or2  I156_038(w_156_038, w_052_1126, w_054_170);
  nand2 I156_041(w_156_041, w_077_494, w_064_677);
  not1 I156_059(w_156_059, w_135_606);
  not1 I156_065(w_156_065, w_061_255);
  not1 I156_124(w_156_124, w_023_642);
  and2 I156_132(w_156_132, w_044_462, w_089_066);
  or2  I156_160(w_156_160, w_015_264, w_030_565);
  nand2 I156_193(w_156_193, w_005_1494, w_030_150);
  or2  I156_322(w_156_322, w_014_309, w_070_391);
  not1 I156_348(w_156_348, w_014_142);
  not1 I156_359(w_156_359, w_128_170);
  nand2 I156_368(w_156_368, w_061_216, w_135_459);
  and2 I156_447(w_156_447, w_074_039, w_038_348);
  nand2 I156_471(w_156_471, w_025_180, w_100_777);
  nand2 I156_497(w_156_497, w_112_602, w_022_045);
  and2 I156_524(w_156_524, w_051_246, w_022_332);
  and2 I156_558(w_156_558, w_005_1551, w_019_905);
  or2  I156_598(w_156_598, w_126_403, w_079_363);
  and2 I157_020(w_157_020, w_097_555, w_067_589);
  or2  I157_040(w_157_040, w_100_550, w_055_423);
  nand2 I157_065(w_157_065, w_081_572, w_039_1232);
  not1 I157_174(w_157_174, w_146_202);
  nand2 I157_188(w_157_188, w_132_011, w_033_001);
  nand2 I157_230(w_157_230, w_108_500, w_153_1324);
  nand2 I157_337(w_157_337, w_119_1092, w_082_691);
  and2 I157_357(w_157_357, w_076_058, w_024_173);
  nand2 I157_405(w_157_405, w_073_011, w_093_062);
  nand2 I157_489(w_157_489, w_025_437, w_082_527);
  or2  I157_563(w_157_563, w_121_704, w_089_377);
  not1 I157_739(w_157_739, w_066_378);
  not1 I157_762(w_157_762, w_034_430);
  not1 I157_993(w_157_993, w_082_510);
  nand2 I157_1078(w_157_1078, w_003_313, w_076_046);
  and2 I157_1082(w_157_1082, w_041_045, w_153_233);
  or2  I157_1161(w_157_1161, w_056_658, w_066_069);
  and2 I157_1237(w_157_1237, w_149_1125, w_091_097);
  or2  I158_036(w_158_036, w_005_830, w_146_220);
  and2 I158_042(w_158_042, w_156_160, w_051_190);
  not1 I158_074(w_158_074, w_114_511);
  not1 I158_092(w_158_092, w_093_005);
  not1 I158_094(w_158_094, w_016_013);
  not1 I158_099(w_158_099, w_129_010);
  and2 I158_122(w_158_122, w_036_037, w_055_090);
  and2 I158_162(w_158_162, w_096_227, w_089_080);
  and2 I158_180(w_158_180, w_095_576, w_022_308);
  and2 I158_205(w_158_205, w_106_1249, w_020_598);
  nand2 I158_257(w_158_257, w_103_523, w_076_049);
  and2 I158_277(w_158_277, w_072_049, w_035_083);
  and2 I158_336(w_158_336, w_055_856, w_041_201);
  not1 I158_355(w_158_355, w_075_097);
  not1 I158_358(w_158_358, w_154_008);
  and2 I158_371(w_158_371, w_138_017, w_026_396);
  not1 I158_375(w_158_375, w_146_366);
  not1 I159_149(w_159_149, w_011_235);
  nand2 I159_186(w_159_186, w_005_1577, w_028_698);
  nand2 I159_215(w_159_215, w_086_108, w_012_229);
  not1 I159_336(w_159_336, w_091_100);
  nand2 I159_344(w_159_344, w_039_1372, w_100_278);
  not1 I159_596(w_159_596, w_035_1502);
  not1 I159_767(w_159_767, w_122_098);
  or2  I159_802(w_159_802, w_091_128, w_020_133);
  and2 I159_806(w_159_806, w_068_197, w_023_596);
  or2  I159_842(w_159_842, w_047_579, w_065_003);
  and2 I159_858(w_159_858, w_121_417, w_092_311);
  not1 I159_974(w_159_974, w_043_043);
  not1 I159_1151(w_159_1151, w_120_165);
  nand2 I159_1268(w_159_1268, w_134_1192, w_061_643);
  not1 I159_1288(w_159_1288, w_107_055);
  nand2 I160_009(w_160_009, w_117_028, w_146_260);
  nand2 I160_016(w_160_016, w_099_214, w_133_147);
  not1 I160_041(w_160_041, w_144_1102);
  or2  I160_053(w_160_053, w_133_475, w_127_802);
  or2  I160_082(w_160_082, w_146_134, w_055_647);
  or2  I160_100(w_160_100, w_126_001, w_062_720);
  or2  I160_145(w_160_145, w_027_409, w_017_269);
  nand2 I160_154(w_160_154, w_098_254, w_095_329);
  and2 I160_196(w_160_196, w_081_415, w_066_562);
  nand2 I160_212(w_160_212, w_010_228, w_131_410);
  nand2 I160_220(w_160_220, w_025_1351, w_058_743);
  nand2 I160_228(w_160_228, w_038_150, w_158_074);
  or2  I160_237(w_160_237, w_062_998, w_009_005);
  not1 I160_337(w_160_337, w_148_806);
  nand2 I160_339(w_160_339, w_010_212, w_024_940);
  not1 I161_027(w_161_027, w_149_594);
  and2 I161_029(w_161_029, w_078_1184, w_079_539);
  or2  I161_072(w_161_072, w_112_865, w_144_609);
  or2  I161_116(w_161_116, w_147_008, w_089_1277);
  nand2 I161_120(w_161_120, w_011_093, w_148_1796);
  and2 I161_121(w_161_121, w_031_594, w_003_015);
  not1 I161_171(w_161_171, w_009_106);
  and2 I161_175(w_161_175, w_065_003, w_103_554);
  not1 I161_178(w_161_178, w_112_707);
  not1 I161_200(w_161_200, w_059_450);
  and2 I161_250(w_161_250, w_044_1330, w_139_076);
  or2  I161_272(w_161_272, w_119_1202, w_055_061);
  or2  I161_298(w_161_298, w_013_170, w_014_144);
  and2 I161_328(w_161_328, w_089_191, w_023_062);
  and2 I161_368(w_161_368, w_040_852, w_017_1595);
  not1 I161_455(w_161_455, w_049_335);
  or2  I161_515(w_161_515, w_034_145, w_157_337);
  and2 I161_520(w_161_520, w_131_071, w_086_677);
  not1 I162_019(w_162_019, w_090_414);
  and2 I162_027(w_162_027, w_144_197, w_158_042);
  nand2 I162_093(w_162_093, w_018_262, w_048_752);
  nand2 I162_105(w_162_105, w_143_370, w_121_102);
  and2 I162_117(w_162_117, w_078_778, w_142_140);
  not1 I162_130(w_162_130, w_067_017);
  nand2 I162_242(w_162_242, w_036_826, w_154_123);
  nand2 I162_278(w_162_278, w_097_556, w_019_951);
  and2 I162_340(w_162_340, w_077_209, w_013_075);
  not1 I162_591(w_162_591, w_123_1084);
  or2  I162_746(w_162_746, w_061_430, w_050_352);
  nand2 I162_795(w_162_795, w_040_757, w_021_226);
  not1 I162_808(w_162_808, w_119_078);
  or2  I162_813(w_162_813, w_127_399, w_086_402);
  nand2 I162_890(w_162_890, w_090_172, w_055_610);
  nand2 I162_894(w_162_894, w_114_1175, w_034_391);
  or2  I162_904(w_162_904, w_100_1408, w_058_828);
  nand2 I163_015(w_163_015, w_123_428, w_060_052);
  and2 I163_041(w_163_041, w_037_1659, w_161_175);
  not1 I163_147(w_163_147, w_146_115);
  not1 I163_216(w_163_216, w_091_065);
  not1 I163_272(w_163_272, w_104_800);
  nand2 I163_290(w_163_290, w_027_204, w_074_954);
  not1 I163_331(w_163_331, w_094_068);
  and2 I163_614(w_163_614, w_075_152, w_007_981);
  or2  I163_779(w_163_779, w_117_179, w_098_498);
  and2 I163_790(w_163_790, w_119_616, w_006_075);
  or2  I163_792(w_163_792, w_050_448, w_150_849);
  or2  I163_1322(w_163_1322, w_118_143, w_142_050);
  or2  I163_1548(w_163_1548, w_141_024, w_086_342);
  or2  I163_1558(w_163_1558, w_034_134, w_121_356);
  not1 I163_1572(w_163_1572, w_106_753);
  or2  I163_1585(w_163_1585, w_006_238, w_145_036);
  not1 I163_1642(w_163_1642, w_027_389);
  or2  I164_034(w_164_034, w_048_142, w_079_577);
  and2 I164_060(w_164_060, w_030_126, w_082_265);
  not1 I164_070(w_164_070, w_150_1759);
  nand2 I164_078(w_164_078, w_044_1505, w_029_628);
  not1 I164_093(w_164_093, w_041_250);
  not1 I164_134(w_164_134, w_149_218);
  or2  I164_146(w_164_146, w_038_111, w_028_300);
  nand2 I164_204(w_164_204, w_044_1268, w_062_1307);
  and2 I164_269(w_164_269, w_110_254, w_085_496);
  or2  I164_307(w_164_307, w_161_027, w_016_009);
  or2  I164_337(w_164_337, w_021_103, w_086_288);
  nand2 I164_359(w_164_359, w_106_533, w_060_080);
  not1 I164_369(w_164_369, w_078_1286);
  or2  I164_498(w_164_498, w_115_376, w_154_148);
  nand2 I164_565(w_164_565, w_048_777, w_149_028);
  not1 I164_732(w_164_732, w_101_655);
  not1 I164_761(w_164_761, w_050_1148);
  not1 I164_782(w_164_782, w_036_842);
  not1 I164_795(w_164_795, w_059_175);
  not1 I164_888(w_164_888, w_129_041);
  nand2 I165_030(w_165_030, w_036_850, w_090_1067);
  or2  I165_058(w_165_058, w_163_272, w_069_1600);
  nand2 I165_106(w_165_106, w_118_721, w_148_530);
  or2  I165_130(w_165_130, w_118_945, w_085_536);
  and2 I165_136(w_165_136, w_110_201, w_031_631);
  not1 I165_163(w_165_163, w_128_133);
  and2 I165_170(w_165_170, w_047_641, w_059_518);
  and2 I165_227(w_165_227, w_009_109, w_016_031);
  nand2 I165_253(w_165_253, w_151_350, w_143_1529);
  nand2 I165_264(w_165_264, w_100_1567, w_060_094);
  or2  I166_048(w_166_048, w_081_532, w_147_041);
  not1 I166_057(w_166_057, w_060_003);
  nand2 I166_104(w_166_104, w_065_001, w_143_1478);
  or2  I166_148(w_166_148, w_079_651, w_011_171);
  or2  I166_162(w_166_162, w_059_383, w_134_352);
  and2 I166_227(w_166_227, w_065_004, w_026_797);
  nand2 I166_233(w_166_233, w_036_914, w_055_786);
  nand2 I166_249(w_166_249, w_087_289, w_145_024);
  not1 I166_333(w_166_333, w_011_144);
  nand2 I166_335(w_166_335, w_139_244, w_111_251);
  or2  I166_509(w_166_509, w_121_240, w_013_278);
  or2  I166_531(w_166_531, w_126_243, w_125_887);
  and2 I166_597(w_166_597, w_002_293, w_127_932);
  nand2 I166_615(w_166_615, w_133_267, w_129_245);
  not1 I166_628(w_166_628, w_029_945);
  nand2 I166_656(w_166_656, w_102_294, w_073_022);
  or2  I166_699(w_166_699, w_002_020, w_014_583);
  or2  I166_812(w_166_812, w_121_103, w_130_977);
  nand2 I167_004(w_167_004, w_072_035, w_076_006);
  or2  I167_006(w_167_006, w_031_021, w_001_048);
  not1 I167_010(w_167_010, w_046_127);
  nand2 I167_012(w_167_012, w_124_740, w_029_402);
  nand2 I167_026(w_167_026, w_031_113, w_098_685);
  not1 I167_028(w_167_028, w_026_275);
  not1 I167_033(w_167_033, w_070_250);
  and2 I167_054(w_167_054, w_058_794, w_155_074);
  or2  I167_055(w_167_055, w_131_1014, w_032_066);
  nand2 I167_059(w_167_059, w_044_115, w_014_038);
  not1 I167_071(w_167_071, w_001_722);
  not1 I167_079(w_167_079, w_144_147);
  or2  I167_088(w_167_088, w_104_430, w_049_738);
  or2  I167_089(w_167_089, w_145_033, w_059_139);
  not1 I167_102(w_167_102, w_010_358);
  not1 I167_127(w_167_127, w_089_604);
  and2 I167_132(w_167_132, w_105_297, w_104_613);
  nand2 I168_005(w_168_005, w_152_367, w_049_909);
  or2  I168_035(w_168_035, w_164_070, w_037_201);
  not1 I168_077(w_168_077, w_038_331);
  and2 I168_225(w_168_225, w_044_1684, w_141_060);
  not1 I168_240(w_168_240, w_099_796);
  and2 I168_259(w_168_259, w_144_965, w_019_019);
  not1 I168_320(w_168_320, w_137_344);
  or2  I168_341(w_168_341, w_160_196, w_073_023);
  not1 I168_399(w_168_399, w_057_1445);
  not1 I168_402(w_168_402, w_089_427);
  nand2 I168_470(w_168_470, w_134_096, w_046_076);
  or2  I168_529(w_168_529, w_132_042, w_039_752);
  and2 I168_608(w_168_608, w_068_021, w_117_492);
  or2  I168_649(w_168_649, w_133_761, w_160_100);
  nand2 I169_068(w_169_068, w_103_329, w_068_189);
  not1 I169_241(w_169_241, w_054_549);
  not1 I169_308(w_169_308, w_142_350);
  or2  I169_372(w_169_372, w_075_167, w_139_1735);
  or2  I169_408(w_169_408, w_047_639, w_007_849);
  and2 I169_480(w_169_480, w_134_828, w_055_243);
  or2  I169_499(w_169_499, w_010_385, w_144_274);
  nand2 I169_507(w_169_507, w_069_1276, w_087_115);
  and2 I169_548(w_169_548, w_156_471, w_056_333);
  nand2 I169_577(w_169_577, w_154_051, w_070_080);
  and2 I169_676(w_169_676, w_080_111, w_026_175);
  nand2 I169_742(w_169_742, w_094_006, w_102_1199);
  nand2 I169_1109(w_169_1109, w_001_1068, w_074_582);
  nand2 I169_1242(w_169_1242, w_144_726, w_000_961);
  nand2 I169_1286(w_169_1286, w_117_148, w_106_764);
  not1 I169_1320(w_169_1320, w_049_429);
  or2  I170_045(w_170_045, w_026_666, w_056_112);
  not1 I170_095(w_170_095, w_000_031);
  or2  I170_167(w_170_167, w_113_771, w_117_1219);
  not1 I170_196(w_170_196, w_153_373);
  or2  I170_322(w_170_322, w_157_188, w_024_1645);
  nand2 I170_364(w_170_364, w_150_817, w_160_016);
  not1 I170_623(w_170_623, w_053_031);
  or2  I170_642(w_170_642, w_054_546, w_103_031);
  or2  I170_766(w_170_766, w_134_804, w_053_077);
  and2 I170_819(w_170_819, w_080_115, w_132_012);
  or2  I170_903(w_170_903, w_123_134, w_107_000);
  or2  I170_947(w_170_947, w_112_137, w_068_163);
  not1 I170_988(w_170_988, w_123_1098);
  or2  I170_991(w_170_991, w_134_468, w_091_033);
  or2  I170_1050(w_170_1050, w_020_685, w_092_335);
  or2  I170_1270(w_170_1270, w_019_808, w_161_120);
  and2 I170_1475(w_170_1475, w_151_922, w_140_406);
  or2  I170_1654(w_170_1654, w_100_1090, w_115_066);
  nand2 I170_1720(w_170_1720, w_055_232, w_109_184);
  or2  I170_1727(w_170_1727, w_025_629, w_050_802);
  nand2 I170_1808(w_170_1808, w_149_252, w_138_010);
  nand2 I170_1844(w_170_1844, w_031_384, w_137_507);
  nand2 I171_037(w_171_037, w_144_704, w_036_451);
  and2 I171_053(w_171_053, w_159_806, w_025_1083);
  not1 I171_085(w_171_085, w_109_039);
  not1 I171_095(w_171_095, w_153_496);
  nand2 I171_101(w_171_101, w_090_413, w_032_058);
  and2 I171_109(w_171_109, w_158_336, w_123_399);
  and2 I171_112(w_171_112, w_019_294, w_138_132);
  or2  I171_152(w_171_152, w_151_370, w_079_564);
  nand2 I171_237(w_171_237, w_169_308, w_050_614);
  nand2 I171_267(w_171_267, w_145_027, w_118_004);
  or2  I171_290(w_171_290, w_114_1212, w_094_036);
  nand2 I171_471(w_171_471, w_037_1462, w_035_574);
  not1 I171_493(w_171_493, w_045_1264);
  not1 I171_505(w_171_505, w_161_272);
  or2  I171_539(w_171_539, w_062_887, w_114_1015);
  not1 I171_593(w_171_593, w_112_296);
  and2 I171_654(w_171_654, w_079_126, w_051_425);
  nand2 I171_704(w_171_704, w_158_180, w_082_734);
  nand2 I171_731(w_171_731, w_169_480, w_128_197);
  nand2 I171_750(w_171_750, w_057_832, w_121_231);
  nand2 I171_794(w_171_794, w_167_132, w_064_193);
  and2 I171_858(w_171_858, w_041_002, w_055_181);
  nand2 I171_971(w_171_971, w_126_363, w_017_774);
  and2 I171_1112(w_171_1112, w_154_000, w_034_590);
  not1 I172_003(w_172_003, w_122_605);
  nand2 I172_004(w_172_004, w_147_074, w_129_607);
  and2 I172_015(w_172_015, w_107_332, w_057_1360);
  and2 I172_046(w_172_046, w_027_277, w_128_109);
  nand2 I172_059(w_172_059, w_121_422, w_064_884);
  nand2 I172_071(w_172_071, w_090_314, w_136_321);
  and2 I172_081(w_172_081, w_045_1052, w_154_015);
  and2 I172_087(w_172_087, w_141_369, w_119_815);
  or2  I172_088(w_172_088, w_156_059, w_100_155);
  not1 I172_095(w_172_095, w_095_900);
  not1 I172_119(w_172_119, w_089_962);
  nand2 I172_120(w_172_120, w_152_176, w_092_129);
  and2 I172_131(w_172_131, w_010_378, w_078_969);
  nand2 I172_145(w_172_145, w_087_1062, w_142_544);
  and2 I172_150(w_172_150, w_016_024, w_088_594);
  not1 I173_079(w_173_079, w_167_033);
  or2  I173_112(w_173_112, w_030_339, w_103_462);
  nand2 I173_258(w_173_258, w_067_376, w_030_742);
  and2 I173_425(w_173_425, w_155_561, w_004_989);
  nand2 I173_447(w_173_447, w_172_088, w_120_152);
  not1 I173_470(w_173_470, w_033_248);
  not1 I173_537(w_173_537, w_123_334);
  nand2 I173_558(w_173_558, w_060_035, w_036_786);
  and2 I173_569(w_173_569, w_068_097, w_017_476);
  and2 I173_612(w_173_612, w_092_158, w_089_438);
  not1 I173_762(w_173_762, w_054_060);
  not1 I173_948(w_173_948, w_040_759);
  and2 I173_991(w_173_991, w_082_120, w_070_379);
  not1 I173_1074(w_173_1074, w_123_088);
  or2  I173_1159(w_173_1159, w_145_038, w_016_011);
  or2  I174_048(w_174_048, w_164_134, w_132_021);
  nand2 I174_073(w_174_073, w_028_066, w_137_039);
  and2 I174_078(w_174_078, w_088_030, w_039_1605);
  or2  I174_324(w_174_324, w_038_353, w_107_432);
  not1 I174_370(w_174_370, w_166_162);
  or2  I174_380(w_174_380, w_010_332, w_099_553);
  not1 I174_392(w_174_392, w_158_358);
  not1 I174_401(w_174_401, w_097_717);
  and2 I174_581(w_174_581, w_172_046, w_019_439);
  and2 I174_624(w_174_624, w_142_649, w_055_494);
  or2  I174_675(w_174_675, w_092_151, w_120_168);
  and2 I174_742(w_174_742, w_028_706, w_077_201);
  or2  I174_780(w_174_780, w_081_578, w_092_129);
  and2 I175_047(w_175_047, w_002_452, w_106_524);
  or2  I175_050(w_175_050, w_058_1019, w_092_648);
  or2  I175_062(w_175_062, w_140_267, w_137_514);
  nand2 I175_064(w_175_064, w_141_148, w_117_099);
  or2  I175_066(w_175_066, w_174_073, w_076_354);
  not1 I175_076(w_175_076, w_132_089);
  nand2 I175_080(w_175_080, w_036_594, w_014_692);
  nand2 I175_084(w_175_084, w_085_059, w_122_202);
  nand2 I175_088(w_175_088, w_169_1286, w_140_1319);
  nand2 I175_090(w_175_090, w_062_418, w_172_004);
  and2 I175_091(w_175_091, w_119_455, w_043_043);
  not1 I175_094(w_175_094, w_074_298);
  or2  I175_102(w_175_102, w_058_1006, w_111_069);
  and2 I175_110(w_175_110, w_132_079, w_131_803);
  nand2 I175_111(w_175_111, w_150_1570, w_013_024);
  and2 I176_041(w_176_041, w_145_023, w_012_639);
  nand2 I176_168(w_176_168, w_172_081, w_100_323);
  not1 I176_212(w_176_212, w_063_1500);
  or2  I176_355(w_176_355, w_078_455, w_162_340);
  not1 I176_366(w_176_366, w_157_489);
  not1 I176_396(w_176_396, w_024_1522);
  or2  I176_449(w_176_449, w_127_482, w_118_360);
  or2  I176_513(w_176_513, w_036_837, w_059_082);
  not1 I176_700(w_176_700, w_144_874);
  or2  I176_763(w_176_763, w_144_058, w_148_1730);
  nand2 I176_823(w_176_823, w_083_001, w_023_775);
  not1 I176_863(w_176_863, w_153_143);
  not1 I176_1151(w_176_1151, w_103_196);
  and2 I176_1327(w_176_1327, w_115_603, w_072_059);
  or2  I176_1462(w_176_1462, w_093_049, w_060_034);
  or2  I177_208(w_177_208, w_006_009, w_000_1242);
  nand2 I177_222(w_177_222, w_027_019, w_032_086);
  nand2 I177_782(w_177_782, w_092_926, w_004_1122);
  not1 I177_900(w_177_900, w_094_013);
  not1 I177_917(w_177_917, w_063_093);
  nand2 I177_1001(w_177_1001, w_104_938, w_016_018);
  and2 I177_1126(w_177_1126, w_018_101, w_113_925);
  not1 I177_1191(w_177_1191, w_006_128);
  nand2 I177_1314(w_177_1314, w_147_036, w_133_907);
  and2 I177_1547(w_177_1547, w_167_012, w_108_734);
  and2 I177_1601(w_177_1601, w_017_1823, w_049_275);
  nand2 I177_1639(w_177_1639, w_022_395, w_173_569);
  or2  I177_1895(w_177_1895, w_119_276, w_116_805);
  and2 I178_031(w_178_031, w_058_521, w_004_182);
  or2  I178_032(w_178_032, w_150_421, w_099_412);
  not1 I178_123(w_178_123, w_087_146);
  or2  I178_285(w_178_285, w_149_381, w_148_274);
  nand2 I178_361(w_178_361, w_156_322, w_016_005);
  and2 I178_365(w_178_365, w_109_162, w_022_382);
  nand2 I178_455(w_178_455, w_097_370, w_035_1146);
  or2  I178_479(w_178_479, w_052_1133, w_020_1222);
  not1 I178_552(w_178_552, w_007_652);
  and2 I178_586(w_178_586, w_105_1809, w_060_060);
  and2 I178_635(w_178_635, w_005_625, w_150_1409);
  or2  I178_658(w_178_658, w_005_844, w_111_666);
  or2  I179_029(w_179_029, w_050_395, w_158_205);
  and2 I179_031(w_179_031, w_056_298, w_056_936);
  not1 I179_116(w_179_116, w_046_083);
  not1 I179_122(w_179_122, w_016_002);
  nand2 I179_222(w_179_222, w_088_139, w_044_1342);
  nand2 I179_226(w_179_226, w_120_104, w_152_169);
  and2 I179_260(w_179_260, w_025_1338, w_112_301);
  not1 I179_351(w_179_351, w_075_065);
  or2  I179_361(w_179_361, w_026_717, w_159_767);
  nand2 I179_397(w_179_397, w_083_003, w_109_208);
  and2 I179_717(w_179_717, w_053_109, w_123_400);
  or2  I179_748(w_179_748, w_157_405, w_103_1313);
  or2  I179_807(w_179_807, w_127_889, w_139_942);
  nand2 I179_974(w_179_974, w_107_286, w_147_153);
  and2 I179_1212(w_179_1212, w_177_782, w_153_745);
  not1 I179_1221(w_179_1221, w_071_303);
  or2  I179_1418(w_179_1418, w_110_529, w_023_811);
  or2  I179_1432(w_179_1432, w_039_610, w_076_311);
  nand2 I179_1625(w_179_1625, w_045_1161, w_111_125);
  and2 I180_015(w_180_015, w_093_023, w_085_576);
  or2  I180_040(w_180_040, w_043_102, w_165_030);
  nand2 I180_056(w_180_056, w_024_918, w_076_149);
  not1 I180_132(w_180_132, w_109_046);
  and2 I180_179(w_180_179, w_024_1404, w_038_378);
  not1 I180_239(w_180_239, w_013_245);
  not1 I180_291(w_180_291, w_143_116);
  not1 I180_313(w_180_313, w_114_252);
  not1 I180_322(w_180_322, w_170_947);
  not1 I180_336(w_180_336, w_157_1078);
  or2  I180_352(w_180_352, w_169_676, w_010_210);
  not1 I180_356(w_180_356, w_010_416);
  or2  I180_418(w_180_418, w_069_1356, w_132_065);
  nand2 I180_422(w_180_422, w_109_335, w_047_007);
  or2  I180_443(w_180_443, w_179_748, w_066_223);
  nand2 I180_447(w_180_447, w_046_266, w_080_061);
  not1 I180_482(w_180_482, w_068_163);
  nand2 I180_529(w_180_529, w_123_984, w_141_077);
  or2  I180_551(w_180_551, w_092_240, w_026_844);
  or2  I180_572(w_180_572, w_152_065, w_156_598);
  not1 I180_575(w_180_575, w_132_017);
  and2 I181_001(w_181_001, w_052_309, w_063_695);
  not1 I181_095(w_181_095, w_160_009);
  nand2 I181_202(w_181_202, w_017_1750, w_157_563);
  nand2 I181_306(w_181_306, w_149_093, w_118_268);
  nand2 I181_478(w_181_478, w_150_1761, w_175_062);
  or2  I181_622(w_181_622, w_085_513, w_066_731);
  or2  I181_782(w_181_782, w_151_553, w_061_426);
  not1 I181_839(w_181_839, w_073_012);
  or2  I181_849(w_181_849, w_040_134, w_096_039);
  nand2 I181_1114(w_181_1114, w_131_311, w_133_719);
  nand2 I182_019(w_182_019, w_146_395, w_145_034);
  and2 I182_066(w_182_066, w_163_790, w_111_331);
  and2 I182_109(w_182_109, w_089_1169, w_097_386);
  nand2 I182_157(w_182_157, w_088_067, w_142_1185);
  not1 I182_194(w_182_194, w_132_046);
  not1 I182_234(w_182_234, w_123_616);
  or2  I182_241(w_182_241, w_096_183, w_073_072);
  and2 I182_243(w_182_243, w_000_1190, w_068_224);
  and2 I182_285(w_182_285, w_053_004, w_034_566);
  and2 I182_309(w_182_309, w_102_519, w_147_176);
  and2 I182_361(w_182_361, w_058_1478, w_056_679);
  and2 I182_398(w_182_398, w_024_211, w_064_891);
  not1 I182_401(w_182_401, w_117_827);
  and2 I182_439(w_182_439, w_070_013, w_006_022);
  nand2 I183_035(w_183_035, w_010_320, w_024_245);
  nand2 I183_051(w_183_051, w_150_1648, w_094_014);
  not1 I183_054(w_183_054, w_029_849);
  and2 I183_130(w_183_130, w_126_270, w_101_166);
  or2  I183_147(w_183_147, w_031_384, w_088_210);
  not1 I183_273(w_183_273, w_177_1895);
  or2  I183_299(w_183_299, w_019_031, w_051_455);
  or2  I183_362(w_183_362, w_102_520, w_050_353);
  or2  I183_438(w_183_438, w_066_909, w_005_1358);
  nand2 I183_455(w_183_455, w_059_561, w_133_214);
  and2 I183_481(w_183_481, w_055_325, w_072_055);
  nand2 I183_686(w_183_686, w_171_750, w_015_091);
  and2 I183_740(w_183_740, w_022_144, w_104_723);
  nand2 I183_998(w_183_998, w_051_582, w_048_792);
  not1 I183_1020(w_183_1020, w_038_028);
  nand2 I183_1069(w_183_1069, w_095_503, w_096_173);
  and2 I183_1281(w_183_1281, w_093_040, w_017_864);
  and2 I183_1551(w_183_1551, w_007_294, w_040_189);
  nand2 I183_1567(w_183_1567, w_140_212, w_059_346);
  nand2 I183_1770(w_183_1770, w_159_149, w_171_731);
  or2  I183_1773(w_183_1773, w_056_650, w_018_244);
  nand2 I183_1795(w_183_1795, w_060_082, w_020_301);
  nand2 I184_001(w_184_001, w_015_056, w_147_053);
  not1 I184_002(w_184_002, w_058_780);
  and2 I184_003(w_184_003, w_145_017, w_118_540);
  and2 I184_004(w_184_004, w_089_222, w_065_000);
  nand2 I184_006(w_184_006, w_042_119, w_118_1079);
  or2  I184_007(w_184_007, w_041_043, w_076_078);
  and2 I184_008(w_184_008, w_039_501, w_074_1265);
  or2  I184_009(w_184_009, w_058_938, w_182_194);
  or2  I184_010(w_184_010, w_046_066, w_168_470);
  or2  I185_077(w_185_077, w_064_728, w_029_679);
  nand2 I185_333(w_185_333, w_063_1247, w_047_174);
  and2 I185_506(w_185_506, w_096_003, w_083_026);
  not1 I185_943(w_185_943, w_039_1151);
  nand2 I185_1010(w_185_1010, w_064_305, w_164_060);
  nand2 I185_1161(w_185_1161, w_063_407, w_133_293);
  not1 I185_1466(w_185_1466, w_151_454);
  and2 I185_1801(w_185_1801, w_082_527, w_108_007);
  not1 I185_1853(w_185_1853, w_147_093);
  and2 I186_000(w_186_000, w_016_021, w_001_006);
  and2 I186_011(w_186_011, w_029_603, w_106_720);
  not1 I186_015(w_186_015, w_013_026);
  and2 I186_025(w_186_025, w_106_848, w_073_004);
  nand2 I186_064(w_186_064, w_071_488, w_165_106);
  and2 I186_119(w_186_119, w_007_136, w_071_437);
  nand2 I186_151(w_186_151, w_044_390, w_142_945);
  nand2 I186_162(w_186_162, w_135_601, w_042_125);
  or2  I186_165(w_186_165, w_015_057, w_143_103);
  nand2 I186_180(w_186_180, w_021_003, w_015_120);
  nand2 I186_191(w_186_191, w_055_370, w_123_455);
  nand2 I186_203(w_186_203, w_131_070, w_018_032);
  nand2 I186_295(w_186_295, w_009_051, w_149_580);
  or2  I186_307(w_186_307, w_155_805, w_015_128);
  or2  I186_315(w_186_315, w_073_016, w_003_132);
  or2  I186_332(w_186_332, w_179_1432, w_059_457);
  not1 I186_344(w_186_344, w_059_008);
  and2 I186_379(w_186_379, w_148_1020, w_072_006);
  or2  I186_385(w_186_385, w_002_193, w_112_804);
  nand2 I187_067(w_187_067, w_164_204, w_181_001);
  nand2 I187_075(w_187_075, w_093_005, w_112_831);
  and2 I187_078(w_187_078, w_098_274, w_186_315);
  or2  I187_081(w_187_081, w_130_707, w_011_459);
  nand2 I187_222(w_187_222, w_008_627, w_176_763);
  nand2 I187_243(w_187_243, w_053_109, w_132_031);
  and2 I187_263(w_187_263, w_133_170, w_004_1649);
  not1 I187_264(w_187_264, w_118_1036);
  nand2 I187_270(w_187_270, w_091_133, w_047_019);
  and2 I187_330(w_187_330, w_164_732, w_091_089);
  not1 I187_346(w_187_346, w_151_097);
  nand2 I187_394(w_187_394, w_062_1296, w_016_001);
  or2  I187_411(w_187_411, w_083_030, w_105_117);
  or2  I187_436(w_187_436, w_085_030, w_036_895);
  nand2 I188_057(w_188_057, w_142_752, w_042_137);
  or2  I188_082(w_188_082, w_022_217, w_024_1261);
  or2  I188_159(w_188_159, w_079_721, w_045_483);
  nand2 I188_178(w_188_178, w_126_165, w_039_1753);
  or2  I188_238(w_188_238, w_071_227, w_076_039);
  not1 I188_247(w_188_247, w_123_865);
  not1 I188_313(w_188_313, w_091_088);
  nand2 I188_329(w_188_329, w_043_063, w_086_1316);
  and2 I188_384(w_188_384, w_028_191, w_124_142);
  not1 I188_417(w_188_417, w_066_558);
  or2  I188_436(w_188_436, w_081_437, w_105_635);
  not1 I188_553(w_188_553, w_078_801);
  or2  I189_010(w_189_010, w_021_010, w_128_002);
  not1 I189_011(w_189_011, w_106_215);
  or2  I189_015(w_189_015, w_144_1387, w_155_838);
  and2 I189_019(w_189_019, w_057_1047, w_043_101);
  not1 I189_024(w_189_024, w_188_247);
  or2  I189_026(w_189_026, w_140_691, w_055_226);
  nand2 I189_043(w_189_043, w_162_019, w_087_1097);
  nand2 I189_052(w_189_052, w_126_138, w_063_1149);
  nand2 I190_004(w_190_004, w_176_212, w_181_782);
  or2  I190_036(w_190_036, w_106_347, w_116_1268);
  and2 I190_121(w_190_121, w_101_033, w_152_253);
  nand2 I190_135(w_190_135, w_050_1369, w_070_459);
  nand2 I190_391(w_190_391, w_058_1346, w_120_141);
  not1 I190_479(w_190_479, w_066_412);
  nand2 I190_664(w_190_664, w_082_422, w_124_393);
  or2  I190_1082(w_190_1082, w_092_396, w_152_081);
  not1 I190_1290(w_190_1290, w_180_056);
  and2 I190_1332(w_190_1332, w_079_202, w_106_1269);
  and2 I190_1392(w_190_1392, w_085_181, w_032_001);
  nand2 I190_1437(w_190_1437, w_070_371, w_100_467);
  nand2 I190_1779(w_190_1779, w_181_622, w_171_109);
  or2  I190_1780(w_190_1780, w_151_1090, w_119_797);
  not1 I191_076(w_191_076, w_114_1047);
  and2 I191_098(w_191_098, w_109_182, w_043_075);
  not1 I191_138(w_191_138, w_138_005);
  nand2 I191_221(w_191_221, w_007_066, w_014_599);
  or2  I191_270(w_191_270, w_043_096, w_124_046);
  or2  I191_375(w_191_375, w_083_005, w_117_394);
  and2 I191_445(w_191_445, w_009_083, w_161_250);
  or2  I191_626(w_191_626, w_051_480, w_151_434);
  not1 I191_793(w_191_793, w_064_364);
  and2 I191_816(w_191_816, w_047_175, w_061_182);
  and2 I191_841(w_191_841, w_028_051, w_011_877);
  and2 I191_1010(w_191_1010, w_109_180, w_140_067);
  not1 I191_1058(w_191_1058, w_155_073);
  and2 I191_1112(w_191_1112, w_169_577, w_171_493);
  or2  I191_1190(w_191_1190, w_115_079, w_019_675);
  or2  I191_1216(w_191_1216, w_166_148, w_160_082);
  nand2 I191_1390(w_191_1390, w_136_629, w_138_040);
  or2  I191_1487(w_191_1487, w_171_237, w_103_994);
  and2 I191_1753(w_191_1753, w_066_430, w_151_1043);
  and2 I192_087(w_192_087, w_037_1532, w_062_497);
  nand2 I192_089(w_192_089, w_047_496, w_057_1817);
  nand2 I192_108(w_192_108, w_132_055, w_045_1590);
  nand2 I192_118(w_192_118, w_104_385, w_174_780);
  nand2 I192_190(w_192_190, w_074_1578, w_093_034);
  and2 I192_318(w_192_318, w_151_179, w_128_222);
  or2  I192_328(w_192_328, w_116_878, w_101_324);
  not1 I192_338(w_192_338, w_016_005);
  and2 I192_346(w_192_346, w_089_1258, w_053_064);
  or2  I192_359(w_192_359, w_095_167, w_071_044);
  or2  I192_382(w_192_382, w_060_016, w_024_1276);
  not1 I192_428(w_192_428, w_084_458);
  not1 I192_461(w_192_461, w_051_1001);
  not1 I192_473(w_192_473, w_107_544);
  or2  I192_486(w_192_486, w_044_784, w_147_190);
  or2  I193_008(w_193_008, w_021_053, w_084_260);
  nand2 I193_032(w_193_032, w_016_003, w_044_1117);
  nand2 I193_095(w_193_095, w_147_189, w_137_339);
  not1 I193_139(w_193_139, w_062_032);
  or2  I193_173(w_193_173, w_016_027, w_050_1537);
  nand2 I193_179(w_193_179, w_143_515, w_158_277);
  or2  I193_189(w_193_189, w_053_045, w_111_029);
  nand2 I193_336(w_193_336, w_112_596, w_009_091);
  and2 I193_422(w_193_422, w_024_028, w_046_274);
  or2  I194_074(w_194_074, w_072_047, w_049_601);
  nand2 I194_103(w_194_103, w_177_1639, w_110_610);
  and2 I194_234(w_194_234, w_123_063, w_143_1469);
  or2  I194_257(w_194_257, w_125_221, w_143_363);
  or2  I194_467(w_194_467, w_056_114, w_182_241);
  not1 I194_552(w_194_552, w_102_130);
  nand2 I194_580(w_194_580, w_004_1281, w_091_141);
  or2  I194_643(w_194_643, w_072_032, w_191_1753);
  or2  I194_705(w_194_705, w_171_704, w_045_335);
  nand2 I194_797(w_194_797, w_119_410, w_110_297);
  not1 I194_853(w_194_853, w_031_762);
  and2 I194_862(w_194_862, w_088_900, w_139_1263);
  or2  I195_041(w_195_041, w_136_511, w_143_404);
  or2  I195_079(w_195_079, w_040_461, w_072_051);
  or2  I195_086(w_195_086, w_040_212, w_026_060);
  not1 I195_194(w_195_194, w_105_1042);
  not1 I195_202(w_195_202, w_012_324);
  nand2 I195_311(w_195_311, w_188_238, w_184_003);
  and2 I195_410(w_195_410, w_089_629, w_053_031);
  not1 I195_498(w_195_498, w_193_008);
  or2  I195_1310(w_195_1310, w_058_1160, w_052_925);
  and2 I195_1332(w_195_1332, w_011_628, w_193_139);
  nand2 I195_1391(w_195_1391, w_175_050, w_122_570);
  not1 I195_1485(w_195_1485, w_001_1276);
  nand2 I196_050(w_196_050, w_152_216, w_026_011);
  or2  I196_160(w_196_160, w_077_642, w_106_334);
  not1 I196_282(w_196_282, w_139_156);
  or2  I196_289(w_196_289, w_061_009, w_161_178);
  not1 I196_349(w_196_349, w_007_725);
  and2 I196_432(w_196_432, w_018_007, w_079_578);
  or2  I196_440(w_196_440, w_180_529, w_130_259);
  and2 I196_463(w_196_463, w_012_353, w_052_952);
  nand2 I196_555(w_196_555, w_145_016, w_149_095);
  not1 I196_697(w_196_697, w_044_087);
  and2 I197_073(w_197_073, w_155_284, w_173_948);
  not1 I197_082(w_197_082, w_149_805);
  or2  I197_288(w_197_288, w_048_202, w_153_728);
  or2  I197_296(w_197_296, w_177_208, w_016_004);
  or2  I197_493(w_197_493, w_030_016, w_079_847);
  and2 I197_707(w_197_707, w_129_332, w_171_290);
  nand2 I197_777(w_197_777, w_156_124, w_160_237);
  and2 I197_860(w_197_860, w_084_317, w_127_783);
  and2 I197_1015(w_197_1015, w_017_967, w_054_220);
  not1 I197_1036(w_197_1036, w_046_251);
  not1 I197_1099(w_197_1099, w_093_040);
  nand2 I197_1182(w_197_1182, w_133_374, w_172_071);
  nand2 I198_122(w_198_122, w_035_640, w_065_001);
  and2 I198_198(w_198_198, w_151_380, w_094_046);
  and2 I198_224(w_198_224, w_027_380, w_081_385);
  nand2 I198_290(w_198_290, w_116_1036, w_004_1831);
  nand2 I198_398(w_198_398, w_005_163, w_172_120);
  or2  I198_481(w_198_481, w_087_1307, w_131_345);
  nand2 I198_625(w_198_625, w_190_121, w_031_828);
  not1 I198_923(w_198_923, w_014_272);
  nand2 I198_926(w_198_926, w_164_337, w_152_220);
  not1 I198_1118(w_198_1118, w_190_135);
  and2 I198_1152(w_198_1152, w_125_362, w_037_1357);
  nand2 I198_1352(w_198_1352, w_171_095, w_001_378);
  not1 I198_1377(w_198_1377, w_066_767);
  nand2 I198_1645(w_198_1645, w_007_194, w_142_457);
  not1 I198_1667(w_198_1667, w_075_049);
  not1 I198_1676(w_198_1676, w_189_026);
  nand2 I198_1725(w_198_1725, w_035_116, w_106_096);
  not1 I199_005(w_199_005, w_048_162);
  nand2 I199_041(w_199_041, w_110_293, w_168_259);
  and2 I199_095(w_199_095, w_113_438, w_030_042);
  or2  I199_127(w_199_127, w_188_057, w_190_036);
  nand2 I199_480(w_199_480, w_174_392, w_087_063);
  and2 I199_620(w_199_620, w_060_055, w_001_1529);
  and2 I199_771(w_199_771, w_029_921, w_052_1621);
  not1 I199_865(w_199_865, w_131_038);
  not1 I199_989(w_199_989, w_136_898);
  or2  I199_1086(w_199_1086, w_061_517, w_157_739);
  not1 I199_1092(w_199_1092, w_043_077);
  not1 I199_1351(w_199_1351, w_094_044);
  or2  I199_1604(w_199_1604, w_172_071, w_084_207);
  and2 I199_1644(w_199_1644, w_033_1210, w_077_664);
  nand2 I200_051(w_200_051, w_139_580, w_144_352);
  nand2 I200_056(w_200_056, w_056_441, w_120_085);
  and2 I200_067(w_200_067, w_068_216, w_173_447);
  or2  I200_137(w_200_137, w_046_270, w_188_313);
  and2 I200_143(w_200_143, w_043_071, w_158_094);
  and2 I200_145(w_200_145, w_007_354, w_007_518);
  nand2 I200_163(w_200_163, w_116_115, w_003_023);
  nand2 I200_197(w_200_197, w_108_266, w_197_707);
  not1 I200_278(w_200_278, w_198_1645);
  nand2 I200_293(w_200_293, w_088_597, w_149_1158);
  not1 I200_312(w_200_312, w_015_136);
  not1 I200_317(w_200_317, w_044_1783);
  nand2 I200_341(w_200_341, w_144_1226, w_106_1235);
  nand2 I200_386(w_200_386, w_060_084, w_120_010);
  and2 I200_395(w_200_395, w_086_748, w_012_460);
  or2  I200_406(w_200_406, w_083_017, w_088_258);
  not1 I200_422(w_200_422, w_078_261);
  not1 I200_432(w_200_432, w_072_013);
  not1 I201_006(w_201_006, w_127_807);
  or2  I201_021(w_201_021, w_104_1694, w_118_651);
  or2  I201_025(w_201_025, w_119_1318, w_123_478);
  or2  I201_029(w_201_029, w_192_108, w_170_1475);
  nand2 I201_031(w_201_031, w_075_184, w_032_206);
  nand2 I201_033(w_201_033, w_138_041, w_181_849);
  nand2 I201_058(w_201_058, w_161_116, w_010_180);
  not1 I201_059(w_201_059, w_200_067);
  or2  I201_117(w_201_117, w_180_443, w_005_786);
  or2  I201_130(w_201_130, w_068_114, w_032_135);
  not1 I201_166(w_201_166, w_021_001);
  not1 I201_184(w_201_184, w_033_1239);
  or2  I201_230(w_201_230, w_125_047, w_191_841);
  or2  I201_265(w_201_265, w_067_763, w_195_498);
  and2 I201_314(w_201_314, w_125_560, w_154_171);
  nand2 I202_090(w_202_090, w_170_1050, w_141_267);
  not1 I202_095(w_202_095, w_061_392);
  not1 I202_356(w_202_356, w_024_1098);
  not1 I202_372(w_202_372, w_164_078);
  or2  I202_431(w_202_431, w_200_056, w_140_100);
  not1 I202_662(w_202_662, w_003_184);
  not1 I202_727(w_202_727, w_111_153);
  and2 I202_782(w_202_782, w_034_559, w_054_540);
  or2  I202_924(w_202_924, w_116_359, w_075_091);
  nand2 I202_1120(w_202_1120, w_088_239, w_201_031);
  or2  I202_1580(w_202_1580, w_051_143, w_011_044);
  and2 I202_1780(w_202_1780, w_039_178, w_163_1322);
  nand2 I203_305(w_203_305, w_140_570, w_176_396);
  not1 I203_384(w_203_384, w_045_752);
  and2 I203_566(w_203_566, w_159_336, w_127_476);
  or2  I203_599(w_203_599, w_076_355, w_027_210);
  or2  I203_650(w_203_650, w_030_630, w_018_142);
  or2  I203_766(w_203_766, w_093_070, w_171_505);
  or2  I204_064(w_204_064, w_126_181, w_049_047);
  not1 I204_196(w_204_196, w_019_165);
  not1 I204_245(w_204_245, w_037_849);
  and2 I204_353(w_204_353, w_143_098, w_009_086);
  and2 I204_438(w_204_438, w_155_174, w_180_015);
  nand2 I204_674(w_204_674, w_197_288, w_191_816);
  nand2 I204_725(w_204_725, w_138_007, w_091_069);
  or2  I204_1002(w_204_1002, w_151_165, w_049_457);
  or2  I204_1159(w_204_1159, w_081_582, w_125_981);
  and2 I204_1212(w_204_1212, w_027_591, w_025_243);
  nand2 I205_298(w_205_298, w_079_536, w_137_389);
  nand2 I205_483(w_205_483, w_041_207, w_069_039);
  and2 I205_554(w_205_554, w_145_005, w_063_1422);
  nand2 I205_699(w_205_699, w_196_349, w_200_312);
  and2 I205_721(w_205_721, w_197_1036, w_146_057);
  nand2 I205_933(w_205_933, w_152_358, w_141_004);
  or2  I205_1143(w_205_1143, w_180_313, w_058_242);
  and2 I206_165(w_206_165, w_193_032, w_056_124);
  and2 I206_484(w_206_484, w_044_794, w_097_743);
  and2 I206_621(w_206_621, w_122_177, w_020_305);
  not1 I206_712(w_206_712, w_025_198);
  nand2 I206_741(w_206_741, w_156_359, w_137_449);
  and2 I206_775(w_206_775, w_018_240, w_177_1314);
  not1 I206_918(w_206_918, w_159_344);
  or2  I206_964(w_206_964, w_133_303, w_120_133);
  nand2 I207_160(w_207_160, w_089_1077, w_176_700);
  and2 I207_233(w_207_233, w_157_040, w_037_649);
  and2 I207_479(w_207_479, w_023_010, w_129_795);
  or2  I207_585(w_207_585, w_164_093, w_034_476);
  and2 I207_587(w_207_587, w_064_1433, w_179_717);
  nand2 I207_668(w_207_668, w_138_058, w_137_146);
  not1 I207_727(w_207_727, w_112_022);
  and2 I207_1006(w_207_1006, w_059_229, w_124_064);
  nand2 I207_1070(w_207_1070, w_022_335, w_038_081);
  and2 I207_1116(w_207_1116, w_079_797, w_151_595);
  nand2 I207_1312(w_207_1312, w_037_1531, w_197_860);
  nand2 I207_1454(w_207_1454, w_183_051, w_088_447);
  not1 I207_1687(w_207_1687, w_171_112);
  and2 I208_175(w_208_175, w_175_110, w_131_847);
  not1 I208_304(w_208_304, w_008_017);
  nand2 I208_305(w_208_305, w_150_1721, w_150_894);
  or2  I208_324(w_208_324, w_189_019, w_109_206);
  not1 I208_518(w_208_518, w_166_048);
  nand2 I208_573(w_208_573, w_052_166, w_095_054);
  or2  I208_663(w_208_663, w_053_050, w_058_1023);
  or2  I208_702(w_208_702, w_182_285, w_104_176);
  or2  I208_813(w_208_813, w_063_270, w_166_335);
  and2 I208_912(w_208_912, w_168_005, w_019_437);
  or2  I208_1069(w_208_1069, w_064_159, w_044_1523);
  not1 I208_1436(w_208_1436, w_110_835);
  and2 I209_000(w_209_000, w_058_649, w_103_1337);
  and2 I209_084(w_209_084, w_057_551, w_141_591);
  and2 I209_174(w_209_174, w_136_458, w_115_111);
  and2 I209_313(w_209_313, w_144_511, w_168_608);
  or2  I209_517(w_209_517, w_034_463, w_060_095);
  or2  I209_638(w_209_638, w_081_223, w_059_065);
  not1 I209_764(w_209_764, w_150_144);
  or2  I209_1088(w_209_1088, w_057_1525, w_008_760);
  or2  I209_1546(w_209_1548, w_015_155, w_209_1547);
  or2  I209_1547(w_209_1549, w_096_042, w_209_1548);
  nand2 I209_1548(w_209_1550, w_189_015, w_209_1549);
  and2 I209_1549(w_209_1551, w_006_088, w_209_1550);
  or2  I209_1550(w_209_1552, w_146_191, w_209_1551);
  nand2 I209_1551(w_209_1553, w_209_1552, w_108_245);
  not1 I209_1552(w_209_1554, w_209_1553);
  nand2 I209_1553(w_209_1555, w_209_1554, w_007_1020);
  and2 I209_1554(w_209_1547, w_209_1555, w_105_074);
  and2 I210_033(w_210_033, w_017_1214, w_124_377);
  nand2 I210_113(w_210_113, w_064_380, w_111_256);
  or2  I210_344(w_210_344, w_081_055, w_167_004);
  not1 I210_367(w_210_367, w_059_065);
  not1 I210_372(w_210_372, w_116_228);
  or2  I210_375(w_210_375, w_043_098, w_006_054);
  nand2 I210_412(w_210_412, w_134_487, w_095_734);
  nand2 I210_428(w_210_428, w_087_1426, w_082_813);
  nand2 I210_430(w_210_430, w_153_843, w_050_1383);
  nand2 I210_614(w_210_614, w_208_1436, w_175_064);
  not1 I210_1039(w_210_1039, w_087_1279);
  or2  I210_1199(w_210_1199, w_199_480, w_198_926);
  not1 I210_1329(w_210_1329, w_141_148);
  nand2 I211_021(w_211_021, w_050_276, w_090_266);
  or2  I211_042(w_211_042, w_191_221, w_027_437);
  and2 I211_043(w_211_043, w_190_1392, w_201_059);
  or2  I211_104(w_211_104, w_184_009, w_176_1151);
  not1 I211_155(w_211_155, w_029_367);
  not1 I211_212(w_211_212, w_111_239);
  and2 I211_294(w_211_294, w_113_432, w_163_779);
  and2 I211_336(w_211_336, w_115_598, w_075_082);
  not1 I211_365(w_211_365, w_186_191);
  and2 I212_009(w_212_009, w_023_158, w_128_012);
  and2 I212_066(w_212_066, w_112_850, w_170_1727);
  or2  I212_134(w_212_134, w_193_179, w_010_108);
  or2  I212_332(w_212_332, w_043_067, w_099_818);
  not1 I212_762(w_212_762, w_037_807);
  and2 I212_1185(w_212_1185, w_142_022, w_183_481);
  and2 I212_1705(w_212_1705, w_052_547, w_113_148);
  or2  I213_020(w_213_020, w_045_1599, w_039_075);
  nand2 I213_021(w_213_021, w_151_765, w_021_218);
  and2 I213_035(w_213_035, w_141_070, w_114_000);
  nand2 I213_041(w_213_041, w_191_1010, w_200_278);
  and2 I213_152(w_213_152, w_099_495, w_180_575);
  nand2 I213_172(w_213_172, w_091_030, w_001_566);
  and2 I213_342(w_213_342, w_118_921, w_185_1010);
  nand2 I213_379(w_213_379, w_116_730, w_095_528);
  not1 I213_423(w_213_423, w_058_1040);
  or2  I213_469(w_213_469, w_089_1140, w_192_461);
  nand2 I213_512(w_213_512, w_043_041, w_068_095);
  and2 I213_562(w_213_562, w_086_742, w_154_015);
  or2  I213_743(w_213_743, w_019_763, w_025_208);
  nand2 I214_015(w_214_015, w_129_066, w_014_132);
  and2 I214_075(w_214_075, w_048_072, w_026_993);
  nand2 I214_078(w_214_078, w_144_014, w_145_012);
  nand2 I214_082(w_214_082, w_147_126, w_173_470);
  nand2 I214_230(w_214_230, w_148_1416, w_020_445);
  and2 I214_277(w_214_277, w_047_329, w_147_080);
  or2  I214_282(w_214_282, w_129_783, w_162_890);
  and2 I214_392(w_214_392, w_139_715, w_190_1779);
  or2  I214_394(w_214_394, w_146_028, w_001_199);
  nand2 I214_401(w_214_401, w_037_502, w_027_122);
  nand2 I214_469(w_214_469, w_086_326, w_188_384);
  nand2 I214_542(w_214_542, w_015_171, w_200_395);
  not1 I214_558(w_214_558, w_213_152);
  or2  I214_568(w_214_568, w_116_364, w_033_1448);
  and2 I214_620(w_214_620, w_030_146, w_169_742);
  and2 I214_697(w_214_697, w_002_144, w_130_195);
  not1 I214_704(w_214_704, w_027_120);
  or2  I214_754(w_214_754, w_146_403, w_103_692);
  or2  I215_125(w_215_125, w_019_002, w_170_642);
  and2 I215_143(w_215_143, w_032_068, w_156_497);
  nand2 I215_199(w_215_199, w_214_401, w_190_1437);
  or2  I215_746(w_215_746, w_163_792, w_128_033);
  and2 I215_1078(w_215_1078, w_070_244, w_212_1705);
  nand2 I216_232(w_216_232, w_139_129, w_019_010);
  nand2 I216_236(w_216_236, w_051_804, w_019_192);
  not1 I216_266(w_216_266, w_080_095);
  nand2 I216_299(w_216_299, w_007_022, w_119_536);
  and2 I216_306(w_216_306, w_178_658, w_039_1768);
  nand2 I216_318(w_216_318, w_119_989, w_214_277);
  and2 I216_467(w_216_467, w_074_246, w_189_052);
  and2 I216_540(w_216_540, w_029_524, w_143_753);
  and2 I216_642(w_216_642, w_120_094, w_040_754);
  and2 I216_644(w_216_644, w_138_101, w_096_225);
  nand2 I216_649(w_216_649, w_208_304, w_155_762);
  or2  I216_667(w_216_667, w_075_179, w_128_038);
  or2  I216_731(w_216_731, w_151_1014, w_113_013);
  and2 I216_743(w_216_743, w_180_447, w_173_112);
  and2 I216_759(w_216_759, w_098_031, w_039_1097);
  or2  I216_873(w_216_873, w_118_342, w_099_1080);
  not1 I216_1118(w_216_1118, w_204_196);
  and2 I216_1133(w_216_1133, w_150_768, w_079_162);
  and2 I217_005(w_217_005, w_056_1391, w_208_305);
  and2 I217_007(w_217_007, w_097_579, w_007_1068);
  nand2 I217_023(w_217_023, w_118_228, w_004_025);
  nand2 I217_031(w_217_031, w_170_623, w_101_244);
  nand2 I217_072(w_217_072, w_105_819, w_211_042);
  or2  I217_073(w_217_073, w_055_363, w_109_340);
  not1 I217_076(w_217_076, w_001_560);
  or2  I217_186(w_217_186, w_207_585, w_084_144);
  and2 I217_197(w_217_197, w_145_032, w_096_162);
  and2 I217_203(w_217_203, w_140_529, w_084_036);
  not1 I218_058(w_218_058, w_122_063);
  not1 I218_066(w_218_066, w_048_546);
  or2  I218_302(w_218_302, w_001_302, w_135_336);
  nand2 I218_338(w_218_338, w_042_065, w_168_402);
  and2 I218_385(w_218_385, w_094_008, w_008_415);
  nand2 I218_388(w_218_388, w_199_989, w_105_1171);
  not1 I218_404(w_218_404, w_049_1165);
  nand2 I218_555(w_218_555, w_170_766, w_211_294);
  not1 I218_637(w_218_637, w_086_909);
  or2  I218_640(w_218_640, w_181_202, w_126_256);
  not1 I218_721(w_218_721, w_206_741);
  or2  I218_739(w_218_739, w_067_160, w_052_574);
  or2  I218_783(w_218_783, w_128_242, w_129_090);
  not1 I218_833(w_218_833, w_108_134);
  not1 I218_1074(w_218_1074, w_180_572);
  or2  I218_1258(w_218_1258, w_073_100, w_184_007);
  or2  I219_020(w_219_020, w_061_548, w_027_512);
  nand2 I219_036(w_219_036, w_035_160, w_050_1433);
  and2 I219_172(w_219_172, w_074_713, w_000_853);
  nand2 I219_184(w_219_184, w_206_775, w_045_1002);
  and2 I220_1285(w_220_1285, w_112_166, w_057_883);
  and2 I221_482(w_221_482, w_144_1570, w_001_1240);
  not1 I221_531(w_221_531, w_063_966);
  or2  I221_1056(w_221_1056, w_184_008, w_016_014);
  and2 I221_1147(w_221_1147, w_217_186, w_146_407);
  and2 I222_066(w_222_066, w_102_594, w_045_574);
  nand2 I222_116(w_222_116, w_072_005, w_021_072);
  not1 I222_411(w_222_411, w_054_469);
  and2 I222_545(w_222_545, w_011_631, w_186_203);
  or2  I222_633(w_222_633, w_173_558, w_030_305);
  nand2 I222_642(w_222_642, w_056_114, w_146_297);
  or2  I222_818(w_222_818, w_180_551, w_159_1288);
  not1 I222_957(w_222_957, w_098_734);
  not1 I222_1038(w_222_1038, w_098_370);
  nand2 I222_1290(w_222_1290, w_067_727, w_098_1010);
  or2  I223_022(w_223_022, w_093_055, w_006_178);
  nand2 I223_179(w_223_179, w_105_1249, w_218_739);
  nand2 I223_221(w_223_221, w_164_359, w_042_118);
  or2  I223_272(w_223_272, w_040_356, w_135_553);
  not1 I223_338(w_223_338, w_150_229);
  or2  I223_536(w_223_536, w_111_482, w_072_053);
  and2 I223_721(w_223_721, w_179_029, w_016_019);
  nand2 I223_990(w_223_990, w_194_862, w_014_156);
  nand2 I223_1010(w_223_1010, w_162_746, w_018_234);
  nand2 I223_1210(w_223_1210, w_209_313, w_174_324);
  or2  I223_1368(w_223_1368, w_118_129, w_089_408);
  not1 I224_049(w_224_049, w_087_462);
  not1 I224_145(w_224_145, w_075_132);
  not1 I224_249(w_224_249, w_125_448);
  nand2 I224_413(w_224_413, w_132_015, w_108_428);
  nand2 I224_605(w_224_605, w_046_248, w_056_1176);
  nand2 I224_834(w_224_834, w_087_607, w_198_1152);
  and2 I225_186(w_225_186, w_200_386, w_216_266);
  not1 I225_276(w_225_276, w_103_146);
  or2  I225_418(w_225_418, w_158_355, w_089_127);
  and2 I225_547(w_225_547, w_091_054, w_151_1378);
  or2  I225_642(w_225_642, w_198_398, w_216_644);
  nand2 I225_802(w_225_802, w_047_562, w_177_917);
  not1 I225_915(w_225_915, w_001_188);
  not1 I225_962(w_225_962, w_064_1643);
  or2  I226_005(w_226_005, w_136_168, w_145_016);
  and2 I226_239(w_226_239, w_095_130, w_013_206);
  and2 I226_257(w_226_257, w_114_294, w_060_100);
  or2  I226_276(w_226_276, w_214_542, w_127_624);
  not1 I226_350(w_226_350, w_204_725);
  or2  I226_439(w_226_439, w_058_616, w_063_1171);
  not1 I226_477(w_226_477, w_160_145);
  and2 I226_631(w_226_631, w_138_049, w_095_834);
  not1 I226_639(w_226_639, w_105_740);
  not1 I226_655(w_226_655, w_214_568);
  or2  I226_665(w_226_665, w_214_620, w_139_348);
  nand2 I227_002(w_227_002, w_145_006, w_122_410);
  and2 I227_009(w_227_009, w_023_339, w_043_063);
  and2 I227_085(w_227_085, w_201_314, w_088_293);
  or2  I227_104(w_227_104, w_171_085, w_062_408);
  nand2 I227_172(w_227_172, w_210_372, w_064_330);
  nand2 I228_032(w_228_032, w_011_809, w_176_366);
  not1 I228_090(w_228_090, w_221_1056);
  or2  I228_137(w_228_137, w_005_542, w_079_145);
  and2 I228_153(w_228_153, w_157_1161, w_020_500);
  and2 I228_179(w_228_179, w_195_079, w_223_1010);
  not1 I228_186(w_228_186, w_083_021);
  or2  I228_194(w_228_194, w_063_1157, w_044_908);
  and2 I229_071(w_229_071, w_117_762, w_043_063);
  nand2 I229_075(w_229_075, w_095_836, w_007_090);
  nand2 I229_192(w_229_192, w_180_322, w_043_042);
  not1 I229_279(w_229_279, w_022_155);
  nand2 I229_1171(w_229_1171, w_027_374, w_056_164);
  and2 I229_1253(w_229_1253, w_161_328, w_030_214);
  not1 I229_1356(w_229_1356, w_076_046);
  or2  I229_1460(w_229_1460, w_144_688, w_093_020);
  or2  I229_1499(w_229_1499, w_003_269, w_112_554);
  or2  I229_1590(w_229_1590, w_132_034, w_157_230);
  nand2 I229_1608(w_229_1608, w_213_342, w_082_358);
  and2 I230_121(w_230_121, w_180_356, w_201_058);
  and2 I230_132(w_230_132, w_211_043, w_082_155);
  or2  I230_237(w_230_237, w_186_385, w_028_313);
  not1 I230_275(w_230_275, w_070_056);
  and2 I230_282(w_230_282, w_008_546, w_067_871);
  nand2 I230_560(w_230_560, w_073_005, w_122_601);
  nand2 I230_594(w_230_594, w_020_696, w_015_127);
  nand2 I230_606(w_230_606, w_020_1265, w_105_476);
  not1 I230_630(w_230_630, w_090_226);
  not1 I231_023(w_231_023, w_155_982);
  nand2 I231_482(w_231_482, w_098_197, w_184_008);
  and2 I231_484(w_231_484, w_222_116, w_124_387);
  nand2 I231_978(w_231_978, w_124_457, w_226_350);
  nand2 I231_1101(w_231_1101, w_117_997, w_150_1283);
  nand2 I231_1104(w_231_1104, w_073_010, w_159_842);
  not1 I231_1239(w_231_1239, w_022_302);
  and2 I231_1269(w_231_1269, w_097_390, w_173_612);
  not1 I231_1286(w_231_1286, w_037_387);
  not1 I231_1321(w_231_1321, w_123_1173);
  nand2 I231_1386(w_231_1386, w_165_264, w_217_007);
  nand2 I231_1618(w_231_1618, w_187_436, w_009_029);
  not1 I231_1772(w_231_1772, w_100_000);
  or2  I232_002(w_232_002, w_154_096, w_201_021);
  not1 I232_153(w_232_153, w_062_447);
  and2 I232_183(w_232_183, w_157_1082, w_007_1388);
  or2  I232_385(w_232_385, w_077_997, w_050_154);
  and2 I232_388(w_232_388, w_058_814, w_205_554);
  nand2 I232_480(w_232_480, w_200_432, w_039_1770);
  not1 I232_507(w_232_507, w_222_957);
  not1 I232_608(w_232_608, w_020_581);
  or2  I232_641(w_232_641, w_083_000, w_128_243);
  and2 I232_667(w_232_667, w_171_794, w_216_667);
  not1 I233_056(w_233_056, w_197_1099);
  not1 I233_083(w_233_083, w_052_1783);
  and2 I233_120(w_233_120, w_172_095, w_066_063);
  not1 I233_152(w_233_152, w_182_109);
  not1 I233_161(w_233_161, w_095_755);
  or2  I233_219(w_233_219, w_188_159, w_203_766);
  nand2 I233_228(w_233_228, w_132_051, w_023_826);
  and2 I233_242(w_233_242, w_075_159, w_195_1310);
  or2  I233_251(w_233_251, w_073_071, w_145_020);
  or2  I233_279(w_233_279, w_036_543, w_186_332);
  or2  I234_011(w_234_011, w_131_031, w_164_269);
  and2 I234_048(w_234_048, w_124_274, w_192_190);
  and2 I234_255(w_234_255, w_176_355, w_229_1608);
  nand2 I234_284(w_234_284, w_006_032, w_115_405);
  nand2 I234_445(w_234_445, w_147_105, w_071_481);
  not1 I234_462(w_234_462, w_133_345);
  and2 I234_587(w_234_587, w_210_033, w_218_721);
  or2  I234_664(w_234_664, w_137_355, w_063_060);
  not1 I234_819(w_234_819, w_024_1079);
  and2 I234_1004(w_234_1004, w_183_1773, w_022_296);
  or2  I234_1075(w_234_1075, w_177_222, w_155_207);
  not1 I234_1138(w_234_1138, w_116_901);
  and2 I235_106(w_235_106, w_216_649, w_088_455);
  nand2 I235_291(w_235_291, w_118_264, w_128_116);
  not1 I235_327(w_235_327, w_210_1329);
  or2  I235_350(w_235_350, w_186_151, w_096_058);
  nand2 I235_371(w_235_371, w_096_012, w_223_272);
  nand2 I235_498(w_235_498, w_125_811, w_221_531);
  nand2 I235_551(w_235_551, w_100_770, w_056_504);
  not1 I235_573(w_235_573, w_064_1658);
  nand2 I235_640(w_235_640, w_070_031, w_187_067);
  not1 I235_669(w_235_669, w_208_813);
  not1 I235_733(w_235_733, w_021_083);
  not1 I235_757(w_235_757, w_119_483);
  or2  I235_791(w_235_791, w_095_020, w_011_372);
  or2  I235_892(w_235_892, w_198_122, w_032_187);
  nand2 I235_947(w_235_947, w_172_131, w_131_127);
  or2  I235_1041(w_235_1043, w_229_1171, w_235_1042);
  nand2 I235_1042(w_235_1044, w_092_881, w_235_1043);
  not1 I235_1043(w_235_1045, w_235_1044);
  and2 I235_1044(w_235_1046, w_028_805, w_235_1045);
  or2  I235_1045(w_235_1047, w_235_1046, w_235_1062);
  or2  I235_1046(w_235_1048, w_235_1047, w_214_282);
  or2  I235_1047(w_235_1042, w_235_1048, w_148_932);
  or2  I235_1048(w_235_1053, w_062_783, w_235_1052);
  and2 I235_1049(w_235_1054, w_192_089, w_235_1053);
  not1 I235_1050(w_235_1055, w_235_1054);
  or2  I235_1051(w_235_1056, w_235_1055, w_017_1706);
  and2 I235_1052(w_235_1057, w_002_177, w_235_1056);
  and2 I235_1053(w_235_1058, w_062_876, w_235_1057);
  or2  I235_1054(w_235_1059, w_235_1058, w_064_1337);
  or2  I235_1055(w_235_1060, w_235_1059, w_124_135);
  not1 I235_1056(w_235_1052, w_235_1047);
  and2 I235_1057(w_235_1062, w_113_814, w_235_1060);
  not1 I236_005(w_236_005, w_105_000);
  or2  I236_099(w_236_099, w_191_1112, w_004_1229);
  and2 I236_182(w_236_182, w_231_1321, w_045_583);
  or2  I236_391(w_236_391, w_073_083, w_107_430);
  not1 I236_403(w_236_403, w_081_619);
  or2  I237_042(w_237_042, w_152_511, w_135_506);
  nand2 I237_138(w_237_138, w_094_085, w_141_009);
  not1 I237_475(w_237_475, w_090_210);
  not1 I237_519(w_237_519, w_228_186);
  not1 I237_569(w_237_569, w_179_116);
  not1 I237_638(w_237_638, w_125_956);
  or2  I237_705(w_237_705, w_130_562, w_111_417);
  and2 I237_819(w_237_819, w_041_035, w_164_034);
  not1 I238_062(w_238_062, w_143_056);
  or2  I238_073(w_238_073, w_191_1487, w_140_442);
  nand2 I238_085(w_238_085, w_215_125, w_225_418);
  nand2 I238_139(w_238_139, w_148_1819, w_134_097);
  not1 I238_143(w_238_143, w_057_1003);
  nand2 I238_272(w_238_272, w_198_1118, w_179_222);
  and2 I238_332(w_238_332, w_129_429, w_218_555);
  not1 I238_366(w_238_366, w_056_023);
  or2  I238_425(w_238_425, w_192_473, w_058_108);
  not1 I238_509(w_238_509, w_218_783);
  nand2 I239_061(w_239_061, w_166_333, w_042_081);
  not1 I239_196(w_239_196, w_087_566);
  and2 I239_367(w_239_367, w_044_201, w_018_129);
  or2  I239_566(w_239_566, w_031_256, w_038_385);
  or2  I239_601(w_239_601, w_001_335, w_063_566);
  or2  I239_726(w_239_726, w_160_339, w_184_002);
  not1 I240_270(w_240_270, w_043_032);
  and2 I240_317(w_240_317, w_175_076, w_165_130);
  or2  I240_427(w_240_427, w_108_054, w_208_324);
  or2  I240_531(w_240_531, w_059_125, w_007_1423);
  and2 I240_576(w_240_576, w_012_497, w_213_035);
  nand2 I240_590(w_240_590, w_166_615, w_043_071);
  and2 I240_888(w_240_888, w_026_318, w_101_203);
  and2 I240_1305(w_240_1305, w_132_043, w_216_759);
  nand2 I241_010(w_241_010, w_023_1273, w_038_459);
  nand2 I241_064(w_241_064, w_197_296, w_187_264);
  not1 I241_096(w_241_096, w_159_1268);
  not1 I241_299(w_241_299, w_104_1546);
  or2  I241_502(w_241_502, w_089_1209, w_093_005);
  not1 I241_1084(w_241_1084, w_003_176);
  or2  I241_1472(w_241_1472, w_180_179, w_015_141);
  not1 I242_001(w_242_001, w_090_615);
  and2 I242_012(w_242_012, w_204_1159, w_051_291);
  not1 I242_014(w_242_014, w_217_197);
  nand2 I242_017(w_242_017, w_200_143, w_125_683);
  or2  I242_030(w_242_030, w_008_670, w_096_108);
  nand2 I242_046(w_242_046, w_005_1519, w_085_363);
  or2  I242_064(w_242_064, w_123_374, w_100_401);
  not1 I242_075(w_242_075, w_019_596);
  or2  I242_084(w_242_084, w_180_132, w_054_057);
  and2 I243_096(w_243_096, w_135_482, w_108_261);
  and2 I243_197(w_243_197, w_216_1133, w_139_404);
  and2 I243_657(w_243_657, w_056_1623, w_112_254);
  or2  I243_851(w_243_851, w_220_1285, w_019_556);
  or2  I243_975(w_243_975, w_166_057, w_010_328);
  not1 I243_1061(w_243_1061, w_172_015);
  and2 I243_1147(w_243_1147, w_044_1629, w_166_104);
  nand2 I243_1362(w_243_1362, w_103_445, w_239_196);
  nand2 I243_1460(w_243_1460, w_112_597, w_054_103);
  or2  I244_026(w_244_026, w_074_128, w_114_490);
  and2 I244_200(w_244_200, w_045_344, w_177_1191);
  not1 I244_317(w_244_317, w_060_040);
  not1 I244_535(w_244_535, w_092_004);
  nand2 I244_543(w_244_543, w_167_088, w_043_070);
  or2  I244_796(w_244_796, w_162_027, w_084_362);
  nand2 I244_892(w_244_892, w_108_207, w_127_697);
  not1 I245_076(w_245_076, w_028_346);
  not1 I245_306(w_245_306, w_176_366);
  or2  I245_1128(w_245_1128, w_170_1720, w_228_179);
  not1 I245_1762(w_245_1762, w_068_239);
  and2 I246_016(w_246_016, w_141_140, w_055_111);
  or2  I246_112(w_246_112, w_033_210, w_167_127);
  nand2 I246_168(w_246_168, w_207_668, w_109_373);
  not1 I246_881(w_246_881, w_054_320);
  nand2 I246_986(w_246_986, w_175_111, w_083_008);
  not1 I246_1367(w_246_1367, w_073_053);
  nand2 I246_1436(w_246_1436, w_089_1266, w_022_362);
  or2  I246_1548(w_246_1548, w_031_153, w_046_145);
  not1 I246_1608(w_246_1608, w_183_130);
  nand2 I247_514(w_247_514, w_152_031, w_083_022);
  not1 I247_604(w_247_604, w_000_1704);
  and2 I247_657(w_247_657, w_213_469, w_238_425);
  or2  I247_759(w_247_759, w_178_635, w_026_1443);
  not1 I247_786(w_247_786, w_136_769);
  not1 I247_877(w_247_877, w_041_254);
  not1 I247_1352(w_247_1352, w_106_172);
  not1 I247_1659(w_247_1659, w_099_037);
  or2  I248_024(w_248_024, w_199_1604, w_135_226);
  and2 I248_028(w_248_028, w_231_1386, w_141_328);
  or2  I248_051(w_248_051, w_218_066, w_088_291);
  or2  I248_059(w_248_059, w_214_015, w_234_284);
  and2 I248_124(w_248_124, w_015_285, w_089_155);
  not1 I248_127(w_248_127, w_231_978);
  not1 I248_147(w_248_147, w_247_514);
  nand2 I248_161(w_248_161, w_211_155, w_213_379);
  and2 I248_291(w_248_291, w_105_012, w_229_192);
  nand2 I248_327(w_248_327, w_088_528, w_040_320);
  and2 I248_354(w_248_354, w_013_142, w_127_251);
  and2 I248_445(w_248_445, w_167_055, w_187_411);
  not1 I248_450(w_248_450, w_078_500);
  nand2 I249_066(w_249_066, w_193_189, w_207_1070);
  nand2 I249_123(w_249_123, w_200_341, w_210_344);
  nand2 I249_423(w_249_423, w_012_535, w_157_174);
  and2 I249_488(w_249_488, w_197_1182, w_104_1049);
  nand2 I249_765(w_249_765, w_101_496, w_197_777);
  or2  I249_943(w_249_943, w_153_505, w_178_123);
  nand2 I250_051(w_250_051, w_121_744, w_246_1548);
  or2  I250_116(w_250_116, w_216_873, w_126_039);
  or2  I250_183(w_250_183, w_011_706, w_167_055);
  not1 I250_207(w_250_207, w_092_517);
  not1 I250_208(w_250_208, w_210_113);
  nand2 I250_222(w_250_222, w_173_537, w_005_022);
  nand2 I250_245(w_250_245, w_106_854, w_224_145);
  and2 I251_010(w_251_010, w_030_727, w_228_137);
  or2  I251_109(w_251_109, w_119_1278, w_112_215);
  or2  I251_123(w_251_123, w_050_368, w_192_328);
  and2 I251_157(w_251_157, w_070_314, w_241_010);
  and2 I251_169(w_251_169, w_250_051, w_040_1003);
  nand2 I251_204(w_251_204, w_036_310, w_040_075);
  and2 I251_245(w_251_245, w_122_436, w_101_566);
  nand2 I251_281(w_251_281, w_018_018, w_152_430);
  and2 I251_282(w_251_282, w_005_610, w_079_848);
  not1 I252_005(w_252_005, w_097_712);
  not1 I252_160(w_252_160, w_037_547);
  or2  I252_191(w_252_191, w_187_222, w_076_057);
  or2  I252_284(w_252_284, w_108_251, w_042_068);
  not1 I252_349(w_252_349, w_080_067);
  and2 I252_382(w_252_382, w_115_212, w_060_034);
  not1 I252_500(w_252_500, w_183_273);
  and2 I252_591(w_252_591, w_115_321, w_044_569);
  nand2 I252_597(w_252_597, w_094_049, w_008_177);
  nand2 I252_617(w_252_617, w_107_651, w_036_815);
  not1 I252_658(w_252_658, w_198_198);
  not1 I253_001(w_253_001, w_159_1151);
  and2 I253_003(w_253_003, w_014_579, w_070_183);
  not1 I253_005(w_253_005, w_222_066);
  or2  I254_015(w_254_015, w_213_562, w_182_234);
  not1 I254_039(w_254_039, w_170_045);
  or2  I254_114(w_254_114, w_146_055, w_229_279);
  nand2 I254_167(w_254_167, w_085_109, w_186_015);
  and2 I254_340(w_254_340, w_234_819, w_235_291);
  not1 I255_042(w_255_042, w_092_970);
  and2 I255_132(w_255_132, w_241_1084, w_010_380);
  nand2 I255_136(w_255_136, w_048_021, w_075_238);
  not1 I255_140(w_255_140, w_180_291);
  not1 I255_196(w_255_196, w_011_470);
  or2  I255_206(w_255_206, w_083_029, w_070_015);
  or2  I255_230(w_255_230, w_138_109, w_057_1060);
  nand2 I255_238(w_255_238, w_179_1418, w_176_041);
  or2  I256_060(w_256_060, w_101_154, w_182_401);
  or2  I256_122(w_256_122, w_046_090, w_030_502);
  not1 I256_321(w_256_321, w_218_833);
  nand2 I256_362(w_256_362, w_112_635, w_235_350);
  or2  I256_421(w_256_421, w_159_186, w_007_961);
  nand2 I256_436(w_256_436, w_007_046, w_184_004);
  not1 I256_496(w_256_496, w_230_275);
  nand2 I256_516(w_256_516, w_108_309, w_153_1016);
  not1 I256_553(w_256_553, w_214_075);
  not1 I256_557(w_256_557, w_034_016);
  or2  I256_622(w_256_622, w_255_238, w_210_614);
  not1 I256_894(w_256_894, w_048_770);
  or2  I256_915(w_256_915, w_143_323, w_140_1423);
  and2 I256_943(w_256_943, w_162_117, w_233_228);
  nand2 I256_957(w_256_957, w_111_383, w_183_147);
  nand2 I257_146(w_257_146, w_166_628, w_024_061);
  and2 I257_235(w_257_235, w_183_1567, w_229_1460);
  and2 I257_360(w_257_360, w_070_005, w_088_189);
  or2  I257_796(w_257_796, w_097_817, w_033_138);
  not1 I257_1198(w_257_1198, w_122_102);
  and2 I257_1239(w_257_1239, w_112_677, w_087_524);
  not1 I257_1369(w_257_1369, w_209_084);
  or2  I257_1467(w_257_1467, w_025_172, w_238_366);
  and2 I258_154(w_258_154, w_084_016, w_240_531);
  and2 I258_178(w_258_178, w_131_011, w_240_270);
  or2  I258_378(w_258_378, w_079_261, w_055_001);
  or2  I258_413(w_258_413, w_046_195, w_136_402);
  nand2 I259_070(w_259_070, w_186_064, w_079_425);
  or2  I259_081(w_259_081, w_030_186, w_088_663);
  nand2 I259_220(w_259_220, w_198_625, w_041_199);
  not1 I259_272(w_259_272, w_106_677);
  and2 I259_392(w_259_392, w_098_263, w_062_240);
  or2  I260_008(w_260_008, w_227_172, w_169_548);
  or2  I260_029(w_260_029, w_112_274, w_117_1471);
  not1 I260_033(w_260_033, w_128_191);
  not1 I260_043(w_260_043, w_028_046);
  or2  I260_048(w_260_048, w_161_029, w_031_284);
  nand2 I261_075(w_261_075, w_199_041, w_202_924);
  not1 I261_128(w_261_128, w_175_110);
  nand2 I261_168(w_261_168, w_260_008, w_147_159);
  nand2 I261_278(w_261_278, w_007_1338, w_216_299);
  or2  I262_119(w_262_119, w_134_430, w_116_421);
  not1 I262_131(w_262_131, w_099_429);
  nand2 I262_144(w_262_144, w_083_022, w_165_163);
  nand2 I262_184(w_262_184, w_218_338, w_108_055);
  nand2 I262_238(w_262_238, w_217_073, w_186_000);
  nand2 I262_290(w_262_290, w_155_1682, w_080_103);
  nand2 I263_000(w_263_000, w_089_328, w_229_075);
  and2 I263_053(w_263_053, w_176_168, w_086_991);
  not1 I263_115(w_263_115, w_167_059);
  nand2 I263_216(w_263_216, w_039_910, w_173_991);
  nand2 I263_293(w_263_293, w_000_1448, w_030_038);
  and2 I263_422(w_263_422, w_127_476, w_228_153);
  or2  I263_426(w_263_426, w_225_642, w_044_778);
  nand2 I263_558(w_263_558, w_167_089, w_218_404);
  not1 I264_021(w_264_021, w_183_455);
  nand2 I264_181(w_264_181, w_105_146, w_182_309);
  or2  I264_257(w_264_257, w_216_467, w_139_001);
  nand2 I264_337(w_264_337, w_075_239, w_012_355);
  and2 I264_425(w_264_425, w_087_1547, w_184_009);
  nand2 I264_430(w_264_430, w_110_625, w_047_141);
  nand2 I264_435(w_264_435, w_211_104, w_183_1281);
  nand2 I264_438(w_264_438, w_059_509, w_033_643);
  or2  I264_518(w_264_518, w_153_156, w_130_000);
  or2  I264_556(w_264_556, w_074_357, w_122_259);
  not1 I265_098(w_265_098, w_176_513);
  not1 I265_127(w_265_127, w_152_249);
  not1 I265_223(w_265_223, w_146_335);
  not1 I265_335(w_265_335, w_153_475);
  not1 I265_375(w_265_375, w_185_1801);
  or2  I265_456(w_265_456, w_132_055, w_042_027);
  nand2 I265_476(w_265_476, w_168_341, w_214_394);
  and2 I265_699(w_265_699, w_111_418, w_162_105);
  and2 I265_1117(w_265_1117, w_104_813, w_002_493);
  nand2 I265_1327(w_265_1327, w_100_472, w_121_524);
  nand2 I265_1382(w_265_1382, w_200_422, w_041_248);
  not1 I265_1397(w_265_1397, w_235_371);
  not1 I266_035(w_266_035, w_154_142);
  nand2 I266_061(w_266_061, w_209_764, w_257_1239);
  or2  I266_233(w_266_233, w_102_507, w_148_715);
  not1 I266_295(w_266_295, w_027_247);
  not1 I266_332(w_266_332, w_122_018);
  nand2 I266_478(w_266_478, w_092_540, w_091_097);
  not1 I266_497(w_266_497, w_105_048);
  not1 I266_543(w_266_543, w_189_015);
  or2  I267_180(w_267_180, w_109_057, w_095_506);
  and2 I267_201(w_267_201, w_123_182, w_091_177);
  nand2 I267_254(w_267_254, w_047_073, w_057_816);
  nand2 I267_329(w_267_329, w_032_224, w_124_061);
  and2 I267_397(w_267_397, w_151_103, w_066_075);
  and2 I267_399(w_267_399, w_049_1157, w_004_1689);
  not1 I267_432(w_267_432, w_181_478);
  and2 I267_476(w_267_476, w_266_061, w_097_887);
  not1 I267_705(w_267_705, w_003_277);
  not1 I267_861(w_267_861, w_145_020);
  or2  I267_865(w_267_865, w_141_495, w_113_1021);
  or2  I268_033(w_268_033, w_138_044, w_152_345);
  or2  I268_357(w_268_357, w_091_145, w_182_398);
  and2 I268_361(w_268_361, w_033_1044, w_190_664);
  or2  I268_1259(w_268_1259, w_111_289, w_119_1282);
  not1 I269_453(w_269_453, w_186_344);
  nand2 I269_1665(w_269_1665, w_107_211, w_000_773);
  and2 I269_1751(w_269_1751, w_135_145, w_137_276);
  or2  I269_1792(w_269_1792, w_208_663, w_098_977);
  nand2 I269_1961(w_269_1961, w_082_265, w_080_110);
  nand2 I269_1979(w_269_1979, w_126_106, w_040_1005);
  nand2 I270_079(w_270_079, w_258_178, w_097_887);
  or2  I270_226(w_270_226, w_107_581, w_267_399);
  nand2 I270_265(w_270_265, w_054_553, w_212_134);
  and2 I270_271(w_270_271, w_066_222, w_095_476);
  and2 I270_345(w_270_345, w_050_185, w_106_585);
  not1 I270_392(w_270_392, w_138_049);
  and2 I270_531(w_270_531, w_234_445, w_264_518);
  or2  I270_663(w_270_663, w_222_545, w_265_1382);
  and2 I271_056(w_271_056, w_252_191, w_081_490);
  nand2 I271_175(w_271_175, w_147_156, w_071_323);
  nand2 I271_200(w_271_200, w_004_719, w_037_1730);
  and2 I271_323(w_271_323, w_150_1118, w_089_693);
  nand2 I271_982(w_271_982, w_188_417, w_058_196);
  or2  I272_054(w_272_054, w_167_079, w_015_170);
  and2 I272_095(w_272_095, w_236_099, w_226_257);
  and2 I272_366(w_272_366, w_083_013, w_183_299);
  or2  I272_662(w_272_662, w_160_053, w_024_1583);
  and2 I272_679(w_272_679, w_111_204, w_267_705);
  or2  I272_972(w_272_972, w_051_422, w_024_299);
  nand2 I272_974(w_272_974, w_242_084, w_026_230);
  nand2 I273_071(w_273_071, w_000_720, w_255_042);
  and2 I273_075(w_273_075, w_199_771, w_009_076);
  nand2 I273_156(w_273_156, w_263_422, w_226_439);
  and2 I273_350(w_273_350, w_171_471, w_263_426);
  not1 I273_376(w_273_376, w_124_662);
  or2  I273_595(w_273_595, w_101_672, w_242_014);
  or2  I273_610(w_273_610, w_018_066, w_063_1561);
  and2 I273_623(w_273_623, w_246_1367, w_111_604);
  or2  I273_751(w_273_751, w_021_261, w_179_1625);
  not1 I273_869(w_273_869, w_192_118);
  nand2 I273_880(w_273_880, w_080_109, w_126_122);
  or2  I274_015(w_274_015, w_035_1475, w_098_389);
  nand2 I274_028(w_274_028, w_019_389, w_054_537);
  nand2 I274_034(w_274_034, w_248_127, w_174_675);
  and2 I274_039(w_274_039, w_001_206, w_192_087);
  or2  I274_044(w_274_044, w_201_006, w_230_630);
  or2  I274_045(w_274_045, w_078_092, w_147_189);
  and2 I274_052(w_274_052, w_060_066, w_075_065);
  or2  I274_054(w_274_054, w_083_031, w_229_1590);
  and2 I274_070(w_274_070, w_208_573, w_022_210);
  or2  I274_071(w_274_071, w_047_537, w_205_483);
  and2 I274_077(w_274_077, w_096_143, w_234_462);
  nand2 I275_027(w_275_027, w_104_663, w_172_059);
  not1 I275_365(w_275_365, w_119_026);
  or2  I275_392(w_275_392, w_072_079, w_109_277);
  not1 I275_420(w_275_420, w_243_1061);
  or2  I275_427(w_275_427, w_272_366, w_189_043);
  or2  I275_486(w_275_486, w_207_1312, w_055_661);
  not1 I275_490(w_275_490, w_140_799);
  and2 I276_024(w_276_024, w_205_298, w_091_022);
  not1 I276_078(w_276_078, w_231_1101);
  nand2 I276_091(w_276_091, w_243_197, w_110_1508);
  and2 I276_119(w_276_119, w_060_033, w_091_003);
  not1 I276_134(w_276_134, w_143_110);
  nand2 I276_145(w_276_145, w_145_032, w_262_144);
  nand2 I276_176(w_276_176, w_158_162, w_070_022);
  not1 I276_188(w_276_188, w_002_191);
  not1 I277_056(w_277_056, w_249_943);
  nand2 I277_085(w_277_085, w_221_1147, w_225_547);
  and2 I277_292(w_277_292, w_030_626, w_109_313);
  not1 I278_052(w_278_052, w_049_253);
  or2  I278_414(w_278_414, w_034_067, w_096_147);
  and2 I278_502(w_278_502, w_058_186, w_267_865);
  nand2 I278_723(w_278_723, w_013_296, w_010_173);
  and2 I278_772(w_278_772, w_218_385, w_151_190);
  not1 I278_946(w_278_946, w_092_1194);
  and2 I278_1207(w_278_1207, w_086_1430, w_153_162);
  nand2 I278_1377(w_278_1377, w_260_033, w_152_142);
  nand2 I279_118(w_279_118, w_166_509, w_092_201);
  and2 I279_187(w_279_187, w_052_731, w_115_410);
  nand2 I279_205(w_279_205, w_085_511, w_040_791);
  and2 I279_250(w_279_250, w_156_065, w_164_795);
  and2 I279_362(w_279_362, w_178_552, w_128_008);
  not1 I279_544(w_279_544, w_267_201);
  not1 I279_570(w_279_570, w_022_039);
  nand2 I279_589(w_279_589, w_012_273, w_050_749);
  nand2 I280_045(w_280_045, w_184_007, w_214_469);
  nand2 I280_266(w_280_266, w_240_317, w_124_488);
  nand2 I280_365(w_280_365, w_150_106, w_076_333);
  not1 I280_389(w_280_389, w_165_170);
  not1 I281_044(w_281_044, w_120_111);
  not1 I281_131(w_281_131, w_216_1118);
  nand2 I281_393(w_281_393, w_008_013, w_029_444);
  or2  I281_595(w_281_595, w_145_015, w_240_576);
  nand2 I281_879(w_281_879, w_062_1222, w_186_011);
  not1 I281_975(w_281_975, w_090_672);
  not1 I282_305(w_282_305, w_267_180);
  nand2 I282_474(w_282_474, w_055_170, w_047_103);
  nand2 I282_537(w_282_537, w_166_249, w_237_705);
  nand2 I282_707(w_282_707, w_098_1076, w_229_071);
  or2  I282_1923(w_282_1923, w_162_904, w_179_260);
  or2  I283_034(w_283_034, w_036_1339, w_070_150);
  or2  I283_086(w_283_086, w_051_046, w_099_714);
  or2  I283_135(w_283_135, w_058_553, w_166_699);
  and2 I283_224(w_283_224, w_191_138, w_155_1152);
  nand2 I283_357(w_283_357, w_207_1687, w_140_483);
  or2  I283_663(w_283_663, w_103_1422, w_047_149);
  or2  I283_992(w_283_992, w_245_076, w_162_808);
  not1 I283_1042(w_283_1042, w_149_090);
  or2  I283_1149(w_283_1149, w_168_529, w_048_797);
  nand2 I283_1219(w_283_1219, w_028_159, w_168_240);
  nand2 I283_1343(w_283_1343, w_046_173, w_006_038);
  or2  I283_1410(w_283_1410, w_274_028, w_127_866);
  nand2 I283_1461(w_283_1461, w_037_674, w_230_282);
  nand2 I283_1561(w_283_1561, w_243_975, w_068_157);
  not1 I283_1724(w_283_1724, w_254_340);
  nand2 I284_047(w_284_047, w_196_050, w_039_289);
  not1 I284_140(w_284_140, w_203_599);
  or2  I284_147(w_284_147, w_179_031, w_211_365);
  or2  I284_819(w_284_819, w_196_463, w_187_346);
  nand2 I284_987(w_284_987, w_190_391, w_282_707);
  or2  I284_1406(w_284_1406, w_266_497, w_283_135);
  not1 I284_1530(w_284_1530, w_112_359);
  and2 I285_021(w_285_021, w_226_005, w_154_182);
  or2  I285_142(w_285_142, w_005_789, w_142_644);
  or2  I285_152(w_285_152, w_003_159, w_154_000);
  not1 I285_264(w_285_264, w_001_210);
  not1 I285_314(w_285_314, w_093_034);
  not1 I285_457(w_285_457, w_184_001);
  or2  I285_470(w_285_470, w_138_004, w_128_197);
  and2 I285_507(w_285_507, w_003_273, w_025_779);
  and2 I285_671(w_285_671, w_167_071, w_217_076);
  and2 I286_076(w_286_076, w_060_057, w_163_216);
  not1 I286_086(w_286_086, w_215_199);
  nand2 I286_163(w_286_163, w_215_143, w_232_667);
  nand2 I286_239(w_286_239, w_204_353, w_095_148);
  not1 I286_530(w_286_530, w_172_150);
  and2 I286_531(w_286_531, w_191_793, w_155_006);
  and2 I286_538(w_286_538, w_176_449, w_225_276);
  or2  I286_539(w_286_539, w_176_863, w_003_259);
  or2  I287_020(w_287_020, w_016_017, w_270_392);
  not1 I287_022(w_287_022, w_007_005);
  nand2 I287_027(w_287_027, w_261_168, w_242_075);
  not1 I287_129(w_287_129, w_052_338);
  not1 I287_148(w_287_148, w_246_1436);
  or2  I287_194(w_287_194, w_103_590, w_076_244);
  and2 I287_271(w_287_271, w_126_139, w_118_481);
  nand2 I287_287(w_287_287, w_202_095, w_249_488);
  or2  I287_352(w_287_352, w_205_721, w_146_120);
  not1 I288_036(w_288_036, w_052_205);
  not1 I288_172(w_288_172, w_131_169);
  and2 I288_272(w_288_272, w_192_318, w_217_023);
  not1 I288_321(w_288_321, w_090_384);
  nand2 I288_700(w_288_700, w_167_102, w_063_966);
  and2 I288_709(w_288_709, w_105_1029, w_248_291);
  and2 I288_823(w_288_823, w_173_425, w_195_202);
  and2 I289_199(w_289_199, w_099_080, w_003_036);
  not1 I289_281(w_289_281, w_265_335);
  or2  I289_377(w_289_377, w_143_347, w_048_672);
  not1 I289_398(w_289_398, w_115_524);
  or2  I289_817(w_289_817, w_105_1812, w_201_130);
  nand2 I289_856(w_289_856, w_113_176, w_272_679);
  and2 I289_921(w_289_921, w_146_375, w_263_115);
  and2 I289_1017(w_289_1017, w_168_077, w_148_903);
  not1 I289_1199(w_289_1199, w_006_099);
  not1 I290_007(w_290_007, w_039_024);
  and2 I290_095(w_290_095, w_057_606, w_198_224);
  not1 I290_110(w_290_110, w_147_040);
  or2  I290_217(w_290_217, w_183_1770, w_029_105);
  not1 I290_254(w_290_254, w_014_136);
  or2  I290_399(w_290_399, w_014_500, w_065_004);
  nand2 I291_126(w_291_126, w_223_990, w_173_258);
  nand2 I291_244(w_291_244, w_004_1674, w_256_516);
  or2  I291_638(w_291_638, w_288_709, w_035_101);
  and2 I291_793(w_291_793, w_166_812, w_137_952);
  or2  I292_019(w_292_019, w_251_245, w_065_003);
  or2  I292_033(w_292_033, w_286_531, w_214_704);
  and2 I292_145(w_292_145, w_027_108, w_128_084);
  or2  I292_461(w_292_461, w_026_161, w_078_1342);
  nand2 I292_557(w_292_557, w_162_813, w_230_594);
  nand2 I292_708(w_292_708, w_190_1290, w_027_029);
  nand2 I292_732(w_292_732, w_109_145, w_041_204);
  not1 I292_765(w_292_765, w_285_264);
  nand2 I292_804(w_292_804, w_281_879, w_089_688);
  or2  I292_892(w_292_892, w_172_003, w_269_1665);
  not1 I293_147(w_293_147, w_256_496);
  not1 I293_212(w_293_212, w_057_1158);
  not1 I293_441(w_293_441, w_272_054);
  and2 I293_464(w_293_464, w_146_007, w_039_260);
  or2  I293_484(w_293_484, w_001_940, w_041_217);
  nand2 I293_535(w_293_535, w_146_234, w_148_1863);
  not1 I293_608(w_293_608, w_278_502);
  or2  I293_660(w_293_660, w_276_024, w_232_507);
  not1 I293_759(w_293_759, w_233_242);
  not1 I293_875(w_293_875, w_152_045);
  not1 I293_989(w_293_989, w_092_526);
  or2  I293_1017(w_293_1017, w_184_010, w_087_590);
  and2 I293_1517(w_293_1517, w_051_294, w_199_095);
  not1 I294_087(w_294_087, w_177_900);
  and2 I294_252(w_294_252, w_233_279, w_026_1407);
  not1 I294_314(w_294_314, w_054_052);
  not1 I294_499(w_294_499, w_246_016);
  not1 I294_564(w_294_564, w_082_240);
  not1 I294_630(w_294_630, w_276_188);
  nand2 I294_813(w_294_813, w_076_240, w_031_395);
  not1 I295_332(w_295_332, w_165_253);
  nand2 I295_369(w_295_369, w_283_086, w_057_915);
  and2 I295_422(w_295_422, w_078_1349, w_153_814);
  not1 I295_546(w_295_546, w_226_276);
  nand2 I295_616(w_295_616, w_109_222, w_010_408);
  and2 I295_718(w_295_718, w_117_651, w_255_140);
  nand2 I295_949(w_295_949, w_075_097, w_294_630);
  nand2 I295_1351(w_295_1351, w_089_524, w_078_055);
  nand2 I295_1365(w_295_1365, w_286_163, w_049_157);
  not1 I296_305(w_296_305, w_100_298);
  nand2 I296_333(w_296_333, w_235_551, w_269_1792);
  not1 I296_491(w_296_491, w_253_001);
  nand2 I296_801(w_296_801, w_066_077, w_072_002);
  or2  I297_041(w_297_041, w_136_806, w_126_105);
  or2  I297_083(w_297_083, w_218_1074, w_047_015);
  or2  I297_111(w_297_111, w_254_167, w_286_086);
  or2  I298_387(w_298_387, w_033_752, w_149_1027);
  and2 I298_578(w_298_578, w_010_202, w_145_005);
  or2  I298_675(w_298_675, w_177_1126, w_165_136);
  or2  I298_828(w_298_828, w_090_457, w_148_490);
  nand2 I298_1289(w_298_1289, w_158_092, w_110_1010);
  or2  I298_1342(w_298_1342, w_218_1258, w_205_1143);
  nand2 I298_1674(w_298_1674, w_233_152, w_248_327);
  not1 I299_086(w_299_086, w_171_267);
  nand2 I299_100(w_299_100, w_126_344, w_131_634);
  not1 I299_113(w_299_113, w_266_295);
  not1 I299_308(w_299_308, w_084_073);
  nand2 I299_340(w_299_340, w_187_078, w_156_348);
  nand2 I299_691(w_299_691, w_028_231, w_107_995);
  not1 I299_740(w_299_740, w_034_185);
  and2 I299_1020(w_299_1020, w_175_084, w_252_284);
  and2 I299_1159(w_299_1159, w_044_1614, w_096_161);
  or2  I299_1179(w_299_1179, w_118_923, w_296_491);
  or2  I299_1221(w_299_1221, w_037_1421, w_033_086);
  and2 I299_1489(w_299_1489, w_207_233, w_209_517);
  nand2 I299_1560(w_299_1560, w_100_1550, w_221_482);
  not1 I299_1758(w_299_1760, w_299_1759);
  nand2 I299_1759(w_299_1761, w_235_733, w_299_1760);
  not1 I299_1760(w_299_1759, w_299_1761);
  not1 I300_014(w_300_014, w_247_786);
  nand2 I300_714(w_300_714, w_275_420, w_088_114);
  not1 I300_853(w_300_853, w_241_1472);
  or2  I300_1378(w_300_1378, w_082_083, w_049_110);
  and2 I300_1448(w_300_1448, w_027_107, w_155_784);
  nand2 I301_1084(w_301_1084, w_035_516, w_240_888);
  not1 I301_1225(w_301_1225, w_262_290);
  or2  I301_1280(w_301_1280, w_269_1961, w_142_557);
  not1 I301_1829(w_301_1829, w_256_122);
  not1 I302_121(w_302_121, w_266_035);
  or2  I302_122(w_302_122, w_061_279, w_131_981);
  nand2 I302_195(w_302_195, w_230_560, w_096_109);
  and2 I302_321(w_302_321, w_090_984, w_283_992);
  not1 I302_402(w_302_402, w_000_1267);
  or2  I302_624(w_302_624, w_049_515, w_290_095);
  nand2 I302_660(w_302_660, w_161_520, w_171_794);
  nand2 I302_1277(w_302_1277, w_219_184, w_206_712);
  not1 I302_1591(w_302_1591, w_070_005);
  not1 I303_008(w_303_008, w_163_1572);
  and2 I303_045(w_303_045, w_186_025, w_078_347);
  and2 I303_690(w_303_690, w_073_090, w_011_079);
  nand2 I304_846(w_304_846, w_060_047, w_008_818);
  and2 I304_1341(w_304_1341, w_008_259, w_169_241);
  nand2 I304_1575(w_304_1575, w_028_381, w_225_915);
  nand2 I304_1593(w_304_1593, w_288_823, w_235_327);
  nand2 I305_000(w_305_000, w_242_012, w_170_095);
  or2  I305_006(w_305_006, w_032_061, w_178_365);
  or2  I305_008(w_305_008, w_293_147, w_034_494);
  and2 I305_011(w_305_011, w_106_089, w_236_403);
  not1 I305_012(w_305_012, w_126_389);
  or2  I305_017(w_305_019, w_003_006, w_305_018);
  not1 I305_018(w_305_020, w_305_019);
  or2  I305_019(w_305_021, w_209_638, w_305_020);
  not1 I305_020(w_305_022, w_305_021);
  not1 I305_021(w_305_023, w_305_022);
  or2  I305_022(w_305_024, w_071_312, w_305_023);
  and2 I305_023(w_305_018, w_185_1853, w_305_024);
  or2  I306_005(w_306_005, w_175_094, w_051_020);
  not1 I306_282(w_306_282, w_146_401);
  not1 I306_427(w_306_427, w_053_032);
  and2 I306_1195(w_306_1195, w_007_793, w_074_278);
  and2 I306_1228(w_306_1228, w_265_223, w_087_1383);
  or2  I306_1282(w_306_1282, w_170_988, w_137_178);
  not1 I307_008(w_307_008, w_112_465);
  or2  I307_013(w_307_013, w_036_1373, w_052_1771);
  nand2 I307_048(w_307_048, w_036_1005, w_122_331);
  and2 I307_119(w_307_119, w_063_613, w_208_518);
  not1 I307_203(w_307_203, w_167_026);
  nand2 I307_230(w_307_230, w_152_417, w_195_410);
  and2 I307_243(w_307_243, w_050_197, w_292_765);
  nand2 I307_271(w_307_271, w_082_414, w_196_697);
  or2  I307_274(w_307_274, w_199_865, w_181_839);
  not1 I308_235(w_308_235, w_242_017);
  and2 I308_256(w_308_256, w_126_420, w_273_071);
  nand2 I308_281(w_308_281, w_018_212, w_090_467);
  nand2 I308_457(w_308_457, w_307_119, w_185_077);
  nand2 I308_778(w_308_778, w_106_380, w_005_1081);
  or2  I308_1117(w_308_1117, w_154_112, w_209_174);
  nand2 I308_1148(w_308_1148, w_100_1177, w_117_142);
  and2 I309_001(w_309_001, w_273_156, w_302_1277);
  or2  I309_086(w_309_086, w_202_356, w_247_1352);
  or2  I309_136(w_309_136, w_231_1618, w_057_250);
  or2  I309_174(w_309_174, w_122_327, w_157_357);
  nand2 I310_019(w_310_019, w_063_1059, w_162_278);
  or2  I310_043(w_310_043, w_226_477, w_070_080);
  or2  I310_065(w_310_065, w_184_009, w_053_014);
  nand2 I310_136(w_310_136, w_069_474, w_273_610);
  nand2 I310_189(w_310_189, w_101_356, w_028_071);
  and2 I310_223(w_310_223, w_198_290, w_171_053);
  not1 I310_274(w_310_274, w_138_106);
  not1 I310_332(w_310_332, w_250_245);
  and2 I310_477(w_310_477, w_170_1844, w_163_1585);
  or2  I310_505(w_310_505, w_231_1239, w_190_1332);
  nand2 I311_135(w_311_135, w_302_624, w_272_972);
  nand2 I311_230(w_311_230, w_006_058, w_302_121);
  and2 I311_245(w_311_245, w_216_731, w_129_744);
  nand2 I311_254(w_311_254, w_179_226, w_195_1332);
  or2  I311_386(w_311_386, w_228_194, w_022_234);
  nand2 I311_453(w_311_453, w_084_343, w_253_001);
  and2 I311_514(w_311_514, w_124_112, w_310_136);
  nand2 I311_641(w_311_641, w_132_057, w_138_100);
  nand2 I312_054(w_312_054, w_197_1015, w_274_045);
  and2 I312_133(w_312_133, w_232_183, w_110_1502);
  nand2 I312_146(w_312_146, w_111_080, w_052_1458);
  nand2 I312_162(w_312_162, w_295_949, w_170_364);
  or2  I312_218(w_312_218, w_158_371, w_104_1704);
  not1 I312_425(w_312_425, w_201_184);
  nand2 I312_514(w_312_514, w_003_007, w_285_457);
  and2 I313_000(w_313_000, w_182_019, w_119_1341);
  and2 I313_001(w_313_001, w_185_506, w_017_174);
  or2  I313_005(w_313_005, w_192_338, w_222_818);
  and2 I313_017(w_313_017, w_125_394, w_056_876);
  nand2 I313_025(w_313_025, w_090_747, w_184_009);
  nand2 I313_028(w_313_028, w_128_176, w_051_571);
  not1 I313_033(w_313_033, w_091_182);
  and2 I314_151(w_314_151, w_144_993, w_051_576);
  nand2 I314_499(w_314_499, w_092_126, w_164_369);
  nand2 I315_093(w_315_093, w_177_1001, w_285_470);
  and2 I315_232(w_315_232, w_049_404, w_069_1285);
  nand2 I315_234(w_315_234, w_089_360, w_227_085);
  or2  I315_444(w_315_444, w_040_981, w_041_156);
  nand2 I315_445(w_315_445, w_061_552, w_161_515);
  and2 I315_556(w_315_556, w_020_648, w_293_989);
  not1 I315_720(w_315_720, w_044_189);
  and2 I316_082(w_316_082, w_244_026, w_073_093);
  nand2 I316_101(w_316_101, w_263_293, w_180_418);
  nand2 I316_288(w_316_288, w_057_1615, w_248_124);
  nand2 I316_510(w_316_510, w_203_305, w_206_484);
  and2 I316_915(w_316_915, w_017_1369, w_240_1305);
  and2 I317_092(w_317_092, w_243_096, w_213_020);
  nand2 I317_649(w_317_649, w_068_085, w_115_333);
  or2  I317_1030(w_317_1030, w_043_016, w_111_151);
  nand2 I317_1544(w_317_1544, w_131_539, w_235_498);
  nand2 I317_1547(w_317_1547, w_266_332, w_032_179);
  not1 I317_1606(w_317_1606, w_054_599);
  not1 I318_012(w_318_012, w_313_017);
  and2 I318_097(w_318_097, w_117_052, w_057_1337);
  or2  I318_192(w_318_192, w_021_195, w_147_198);
  not1 I318_277(w_318_277, w_089_067);
  nand2 I318_336(w_318_336, w_135_182, w_084_391);
  and2 I318_360(w_318_360, w_178_031, w_084_333);
  nand2 I318_507(w_318_507, w_041_178, w_202_782);
  not1 I319_307(w_319_307, w_040_203);
  and2 I319_1589(w_319_1589, w_310_043, w_142_776);
  not1 I320_201(w_320_201, w_145_035);
  or2  I320_214(w_320_214, w_024_289, w_254_039);
  or2  I320_484(w_320_484, w_105_671, w_042_018);
  nand2 I320_632(w_320_632, w_237_569, w_072_077);
  not1 I321_082(w_321_082, w_096_073);
  not1 I321_092(w_321_092, w_261_128);
  not1 I321_097(w_321_097, w_134_375);
  not1 I321_120(w_321_120, w_251_109);
  and2 I321_129(w_321_129, w_037_567, w_194_234);
  not1 I321_196(w_321_196, w_270_226);
  nand2 I322_112(w_322_112, w_296_333, w_111_447);
  or2  I322_143(w_322_143, w_263_216, w_275_365);
  nand2 I322_296(w_322_296, w_139_069, w_165_058);
  nand2 I322_1155(w_322_1155, w_064_1204, w_223_536);
  nand2 I323_111(w_323_111, w_279_362, w_115_540);
  nand2 I323_288(w_323_288, w_267_397, w_118_1139);
  nand2 I323_305(w_323_305, w_307_230, w_071_056);
  and2 I323_309(w_323_309, w_115_460, w_243_1460);
  not1 I323_312(w_323_312, w_178_479);
  or2  I323_386(w_323_386, w_071_341, w_245_306);
  not1 I323_403(w_323_403, w_216_236);
  nand2 I323_446(w_323_446, w_169_499, w_059_020);
  nand2 I323_461(w_323_461, w_186_379, w_038_320);
  nand2 I324_008(w_324_008, w_253_001, w_158_036);
  or2  I324_092(w_324_092, w_131_766, w_063_1411);
  not1 I324_105(w_324_105, w_037_226);
  nand2 I324_145(w_324_145, w_028_479, w_055_044);
  not1 I324_183(w_324_183, w_253_003);
  nand2 I324_469(w_324_469, w_272_095, w_103_718);
  and2 I324_530(w_324_530, w_298_1674, w_011_103);
  and2 I324_742(w_324_742, w_079_588, w_117_017);
  and2 I325_661(w_325_661, w_297_111, w_125_397);
  nand2 I325_1102(w_325_1102, w_265_375, w_170_322);
  or2  I325_1215(w_325_1215, w_145_036, w_047_253);
  nand2 I325_1228(w_325_1228, w_172_145, w_279_589);
  not1 I325_1468(w_325_1468, w_154_106);
  and2 I325_1534(w_325_1534, w_064_926, w_120_152);
  not1 I326_363(w_326_363, w_315_445);
  or2  I326_383(w_326_383, w_257_1198, w_101_615);
  or2  I326_737(w_326_737, w_031_684, w_321_120);
  not1 I326_1155(w_326_1155, w_201_265);
  not1 I327_290(w_327_290, w_047_442);
  or2  I327_428(w_327_428, w_142_697, w_125_1361);
  not1 I327_516(w_327_516, w_270_345);
  and2 I327_519(w_327_519, w_199_1351, w_139_120);
  nand2 I327_1023(w_327_1023, w_024_081, w_105_063);
  nand2 I327_1107(w_327_1107, w_010_163, w_212_1185);
  not1 I328_005(w_328_005, w_175_090);
  nand2 I328_006(w_328_006, w_161_368, w_080_119);
  nand2 I328_008(w_328_008, w_084_080, w_310_274);
  and2 I328_010(w_328_010, w_064_036, w_324_183);
  or2  I328_013(w_328_013, w_267_861, w_293_464);
  or2  I329_059(w_329_059, w_013_069, w_178_361);
  and2 I329_203(w_329_203, w_106_043, w_259_220);
  not1 I329_228(w_329_228, w_092_1039);
  nand2 I329_249(w_329_249, w_103_375, w_020_139);
  not1 I329_262(w_329_262, w_118_692);
  not1 I329_460(w_329_460, w_137_463);
  and2 I330_248(w_330_248, w_213_172, w_112_552);
  and2 I330_693(w_330_693, w_238_085, w_013_253);
  or2  I330_731(w_330_731, w_308_1117, w_032_208);
  or2  I330_753(w_330_753, w_100_576, w_195_194);
  not1 I330_814(w_330_814, w_256_943);
  not1 I330_958(w_330_958, w_289_199);
  and2 I330_1024(w_330_1024, w_293_484, w_112_279);
  not1 I331_107(w_331_107, w_156_023);
  nand2 I331_550(w_331_550, w_026_379, w_004_1613);
  and2 I331_838(w_331_838, w_055_435, w_091_090);
  not1 I331_899(w_331_899, w_149_581);
  or2  I332_063(w_332_063, w_120_041, w_001_861);
  and2 I332_177(w_332_177, w_231_1269, w_005_1467);
  and2 I332_319(w_332_319, w_324_530, w_274_077);
  not1 I332_572(w_332_572, w_226_631);
  and2 I332_617(w_332_617, w_206_964, w_101_367);
  or2  I332_1090(w_332_1090, w_295_1351, w_313_001);
  or2  I333_070(w_333_070, w_038_308, w_295_718);
  and2 I334_223(w_334_223, w_091_124, w_009_009);
  and2 I334_261(w_334_261, w_071_339, w_328_010);
  nand2 I334_343(w_334_343, w_040_011, w_121_486);
  not1 I334_566(w_334_566, w_234_255);
  or2  I334_567(w_334_567, w_215_746, w_201_029);
  nand2 I334_597(w_334_597, w_201_033, w_060_069);
  not1 I334_650(w_334_650, w_224_834);
  and2 I335_006(w_335_006, w_063_041, w_272_974);
  nand2 I335_072(w_335_072, w_193_422, w_291_638);
  or2  I335_362(w_335_362, w_065_003, w_156_368);
  not1 I336_141(w_336_141, w_112_034);
  and2 I336_181(w_336_181, w_052_1284, w_207_160);
  nand2 I336_577(w_336_577, w_263_000, w_083_030);
  or2  I336_663(w_336_663, w_013_145, w_303_690);
  or2  I336_1049(w_336_1049, w_078_872, w_095_099);
  and2 I336_1116(w_336_1116, w_048_963, w_103_062);
  nand2 I336_1225(w_336_1225, w_314_151, w_241_502);
  not1 I336_1630(w_336_1630, w_300_714);
  or2  I337_027(w_337_027, w_132_015, w_006_153);
  not1 I337_038(w_337_038, w_200_145);
  and2 I337_094(w_337_094, w_200_163, w_265_127);
  nand2 I337_158(w_337_158, w_327_1023, w_257_796);
  and2 I337_234(w_337_234, w_183_740, w_034_405);
  not1 I337_266(w_337_266, w_140_045);
  or2  I337_369(w_337_369, w_161_298, w_334_223);
  nand2 I338_073(w_338_073, w_231_023, w_320_201);
  nand2 I338_1435(w_338_1435, w_064_085, w_005_024);
  nand2 I338_1654(w_338_1654, w_251_281, w_231_1286);
  nand2 I338_1705(w_338_1705, w_214_082, w_125_1050);
  or2  I339_121(w_339_121, w_143_466, w_293_1517);
  and2 I339_235(w_339_235, w_262_238, w_140_745);
  nand2 I339_405(w_339_405, w_066_823, w_244_543);
  or2  I339_439(w_339_439, w_191_270, w_048_671);
  nand2 I339_524(w_339_524, w_014_008, w_080_007);
  or2  I340_114(w_340_114, w_027_430, w_179_974);
  or2  I341_141(w_341_141, w_035_117, w_191_1216);
  and2 I341_249(w_341_249, w_318_360, w_267_254);
  nand2 I341_302(w_341_302, w_100_186, w_299_1489);
  or2  I342_013(w_342_013, w_061_212, w_020_1155);
  not1 I342_1028(w_342_1028, w_101_437);
  and2 I342_1576(w_342_1576, w_252_591, w_011_680);
  or2  I342_1767(w_342_1769, w_309_174, w_342_1768);
  and2 I342_1768(w_342_1770, w_323_305, w_342_1769);
  not1 I342_1769(w_342_1771, w_342_1770);
  not1 I342_1770(w_342_1772, w_342_1771);
  or2  I342_1771(w_342_1773, w_264_438, w_342_1772);
  or2  I342_1772(w_342_1774, w_129_681, w_342_1773);
  or2  I342_1773(w_342_1775, w_342_1774, w_342_1788);
  and2 I342_1774(w_342_1776, w_156_524, w_342_1775);
  and2 I342_1775(w_342_1777, w_166_233, w_342_1776);
  and2 I342_1776(w_342_1768, w_342_1777, w_149_329);
  and2 I342_1777(w_342_1782, w_216_743, w_342_1781);
  or2  I342_1778(w_342_1783, w_342_1782, w_305_000);
  not1 I342_1779(w_342_1784, w_342_1783);
  and2 I342_1780(w_342_1785, w_083_008, w_342_1784);
  and2 I342_1781(w_342_1786, w_311_514, w_342_1785);
  not1 I342_1782(w_342_1781, w_342_1775);
  and2 I342_1783(w_342_1788, w_089_647, w_342_1786);
  and2 I343_016(w_343_016, w_295_332, w_014_659);
  nand2 I343_227(w_343_227, w_039_1891, w_053_098);
  nand2 I343_894(w_343_894, w_161_072, w_197_082);
  nand2 I343_1177(w_343_1177, w_138_008, w_044_718);
  or2  I344_052(w_344_052, w_301_1084, w_002_035);
  and2 I344_117(w_344_117, w_084_168, w_184_007);
  or2  I344_139(w_344_139, w_280_266, w_015_127);
  and2 I344_141(w_344_141, w_086_1168, w_082_529);
  or2  I344_150(w_344_150, w_174_401, w_293_759);
  nand2 I344_207(w_344_207, w_322_296, w_337_094);
  not1 I345_1056(w_345_1056, w_202_431);
  not1 I345_1240(w_345_1240, w_158_122);
  and2 I345_1481(w_345_1481, w_324_092, w_047_100);
  and2 I346_341(w_346_341, w_043_064, w_098_004);
  not1 I346_528(w_346_528, w_040_353);
  nand2 I346_640(w_346_640, w_288_700, w_082_745);
  nand2 I346_679(w_346_679, w_117_365, w_327_519);
  nand2 I347_053(w_347_053, w_294_252, w_153_641);
  nand2 I347_705(w_347_705, w_256_915, w_232_641);
  or2  I347_950(w_347_950, w_082_303, w_115_501);
  and2 I347_1219(w_347_1219, w_282_474, w_160_154);
  and2 I347_1311(w_347_1311, w_243_851, w_046_168);
  not1 I347_1576(w_347_1576, w_274_052);
  not1 I347_1601(w_347_1601, w_186_295);
  and2 I348_167(w_348_167, w_039_033, w_188_436);
  nand2 I349_052(w_349_052, w_198_1725, w_086_235);
  or2  I349_104(w_349_104, w_334_343, w_260_043);
  or2  I350_207(w_350_207, w_167_132, w_199_1086);
  not1 I350_314(w_350_314, w_183_1020);
  not1 I350_377(w_350_377, w_287_287);
  and2 I350_444(w_350_444, w_186_162, w_275_486);
  nand2 I350_527(w_350_527, w_087_304, w_157_065);
  or2  I350_529(w_350_529, w_111_264, w_019_865);
  not1 I351_000(w_351_000, w_069_1818);
  or2  I351_021(w_351_021, w_022_003, w_085_505);
  not1 I351_028(w_351_028, w_263_053);
  and2 I351_035(w_351_035, w_216_232, w_081_093);
  or2  I352_320(w_352_320, w_074_869, w_238_139);
  and2 I352_406(w_352_406, w_014_487, w_133_042);
  not1 I352_422(w_352_422, w_132_043);
  and2 I352_672(w_352_672, w_332_572, w_237_475);
  and2 I353_138(w_353_138, w_148_120, w_072_005);
  and2 I353_181(w_353_181, w_056_929, w_191_1058);
  nand2 I353_240(w_353_240, w_022_061, w_256_553);
  nand2 I353_380(w_353_380, w_134_006, w_087_840);
  not1 I353_448(w_353_448, w_145_037);
  and2 I353_531(w_353_531, w_076_208, w_108_067);
  nand2 I353_691(w_353_691, w_108_652, w_137_871);
  nand2 I353_720(w_353_720, w_283_663, w_224_605);
  and2 I353_985(w_353_985, w_020_015, w_307_048);
  not1 I353_1174(w_353_1174, w_223_338);
  and2 I354_064(w_354_064, w_135_378, w_300_1378);
  or2  I354_278(w_354_278, w_211_021, w_306_005);
  and2 I354_391(w_354_391, w_025_298, w_311_254);
  not1 I354_412(w_354_412, w_353_138);
  or2  I354_460(w_354_460, w_148_1903, w_258_154);
  and2 I354_1250(w_354_1250, w_120_047, w_342_013);
  nand2 I354_1261(w_354_1261, w_093_062, w_163_614);
  and2 I355_018(w_355_018, w_235_640, w_286_539);
  or2  I355_076(w_355_076, w_352_320, w_179_1212);
  not1 I355_089(w_355_089, w_342_1576);
  or2  I355_155(w_355_155, w_298_387, w_191_375);
  and2 I355_213(w_355_213, w_216_318, w_066_602);
  or2  I355_226(w_355_226, w_162_591, w_309_136);
  and2 I355_291(w_355_291, w_136_823, w_053_014);
  not1 I355_525(w_355_525, w_208_1069);
  nand2 I356_068(w_356_068, w_157_1237, w_083_001);
  and2 I356_335(w_356_335, w_272_662, w_009_026);
  or2  I356_714(w_356_714, w_299_1179, w_136_665);
  not1 I357_026(w_357_026, w_207_727);
  not1 I357_083(w_357_083, w_007_043);
  not1 I357_141(w_357_141, w_059_014);
  or2  I357_293(w_357_293, w_204_245, w_302_1591);
  not1 I357_401(w_357_401, w_105_1183);
  nand2 I358_471(w_358_471, w_347_950, w_123_237);
  nand2 I358_675(w_358_675, w_351_035, w_172_087);
  not1 I358_692(w_358_692, w_330_814);
  nand2 I358_1178(w_358_1178, w_073_034, w_347_705);
  or2  I358_1499(w_358_1499, w_170_1808, w_028_038);
  or2  I359_131(w_359_131, w_182_361, w_319_1589);
  nand2 I359_526(w_359_526, w_029_1059, w_248_445);
  not1 I359_650(w_359_650, w_224_049);
  not1 I359_1125(w_359_1125, w_140_1596);
  or2  I360_496(w_360_496, w_103_064, w_128_264);
  and2 I360_542(w_360_542, w_135_570, w_209_000);
  nand2 I360_762(w_360_762, w_279_118, w_057_284);
  not1 I361_090(w_361_090, w_144_1115);
  or2  I361_238(w_361_238, w_325_1215, w_143_1344);
  and2 I361_317(w_361_317, w_022_234, w_184_003);
  or2  I362_105(w_362_105, w_332_319, w_122_572);
  or2  I362_212(w_362_212, w_137_007, w_352_406);
  or2  I362_293(w_362_293, w_329_249, w_291_126);
  and2 I362_337(w_362_337, w_323_309, w_028_636);
  not1 I362_481(w_362_481, w_217_072);
  nand2 I362_483(w_362_483, w_026_570, w_194_467);
  not1 I362_1655(w_362_1655, w_161_121);
  not1 I363_075(w_363_075, w_285_152);
  and2 I363_507(w_363_507, w_318_507, w_061_633);
  and2 I363_598(w_363_598, w_350_377, w_139_1379);
  nand2 I363_803(w_363_803, w_110_1241, w_171_593);
  or2  I364_185(w_364_185, w_154_071, w_057_653);
  or2  I364_233(w_364_233, w_320_214, w_354_412);
  not1 I364_722(w_364_722, w_026_480);
  or2  I364_1423(w_364_1423, w_292_557, w_041_064);
  nand2 I365_064(w_365_064, w_298_675, w_217_005);
  or2  I365_198(w_365_198, w_151_1182, w_352_422);
  and2 I365_216(w_365_216, w_104_684, w_121_501);
  or2  I365_534(w_365_534, w_317_1606, w_350_444);
  or2  I365_536(w_365_536, w_256_321, w_335_362);
  and2 I365_620(w_365_620, w_231_484, w_054_444);
  nand2 I365_832(w_365_832, w_012_271, w_164_307);
  not1 I365_858(w_365_858, w_239_726);
  and2 I366_011(w_366_011, w_236_005, w_216_642);
  not1 I367_489(w_367_489, w_185_943);
  nand2 I368_156(w_368_156, w_062_689, w_287_129);
  and2 I368_455(w_368_455, w_143_941, w_012_522);
  not1 I368_653(w_368_653, w_203_566);
  nand2 I368_783(w_368_783, w_098_801, w_110_914);
  nand2 I368_986(w_368_986, w_091_140, w_289_817);
  or2  I368_1314(w_368_1314, w_303_008, w_257_146);
  nand2 I368_1526(w_368_1526, w_116_599, w_317_092);
  and2 I368_1696(w_368_1696, w_300_853, w_072_054);
  and2 I369_228(w_369_228, w_161_200, w_354_391);
  and2 I369_346(w_369_346, w_163_331, w_083_010);
  nand2 I369_649(w_369_649, w_154_013, w_183_686);
  not1 I369_1046(w_369_1046, w_316_082);
  nand2 I369_1193(w_369_1193, w_146_418, w_182_157);
  not1 I369_1531(w_369_1531, w_287_194);
  or2  I370_066(w_370_066, w_160_337, w_005_357);
  not1 I370_067(w_370_067, w_230_606);
  and2 I370_077(w_370_077, w_071_523, w_141_255);
  and2 I370_616(w_370_616, w_318_097, w_063_194);
  not1 I370_890(w_370_890, w_311_230);
  or2  I370_1007(w_370_1007, w_201_025, w_019_525);
  not1 I370_1459(w_370_1459, w_121_092);
  not1 I371_092(w_371_092, w_055_525);
  not1 I371_098(w_371_098, w_189_010);
  or2  I371_343(w_371_343, w_233_161, w_251_123);
  and2 I371_387(w_371_387, w_015_232, w_044_791);
  or2  I371_548(w_371_548, w_102_931, w_064_1456);
  and2 I371_710(w_371_710, w_190_004, w_103_1398);
  or2  I372_215(w_372_215, w_082_337, w_125_175);
  nand2 I372_317(w_372_317, w_184_003, w_276_119);
  and2 I372_366(w_372_366, w_369_649, w_148_1503);
  or2  I372_404(w_372_404, w_070_427, w_292_033);
  not1 I372_428(w_372_428, w_241_096);
  or2  I373_465(w_373_465, w_186_307, w_016_011);
  nand2 I373_471(w_373_471, w_122_556, w_213_021);
  or2  I373_1442(w_373_1442, w_072_079, w_172_119);
  and2 I373_1800(w_373_1800, w_160_228, w_069_1807);
  and2 I374_012(w_374_012, w_219_036, w_174_380);
  nand2 I374_145(w_374_145, w_246_881, w_158_277);
  or2  I374_304(w_374_304, w_355_076, w_001_717);
  and2 I374_798(w_374_798, w_131_376, w_082_589);
  nand2 I374_1192(w_374_1192, w_329_228, w_053_105);
  nand2 I374_1496(w_374_1496, w_187_330, w_109_032);
  and2 I375_1233(w_375_1233, w_374_012, w_233_251);
  or2  I376_209(w_376_209, w_035_004, w_048_253);
  and2 I376_513(w_376_513, w_337_038, w_092_091);
  not1 I376_677(w_376_677, w_035_397);
  or2  I376_750(w_376_750, w_026_1260, w_127_734);
  nand2 I377_072(w_377_072, w_111_292, w_077_658);
  not1 I377_193(w_377_193, w_271_323);
  not1 I377_256(w_377_256, w_028_748);
  nand2 I378_048(w_378_048, w_377_256, w_232_608);
  nand2 I378_278(w_378_278, w_168_035, w_213_423);
  nand2 I378_565(w_378_565, w_244_317, w_210_430);
  or2  I378_597(w_378_597, w_026_777, w_130_221);
  or2  I379_043(w_379_043, w_245_1762, w_060_020);
  or2  I379_194(w_379_194, w_347_1576, w_102_010);
  not1 I379_781(w_379_781, w_284_819);
  and2 I379_829(w_379_829, w_046_255, w_175_047);
  nand2 I380_321(w_380_321, w_196_160, w_141_336);
  nand2 I380_434(w_380_434, w_087_110, w_237_569);
  nand2 I381_179(w_381_179, w_252_597, w_104_1580);
  and2 I381_531(w_381_531, w_315_093, w_241_064);
  and2 I381_634(w_381_634, w_378_278, w_077_151);
  nand2 I381_839(w_381_839, w_042_107, w_265_098);
  and2 I382_163(w_382_163, w_336_1225, w_338_1705);
  nand2 I382_185(w_382_185, w_218_640, w_356_714);
  not1 I382_653(w_382_653, w_279_544);
  and2 I382_672(w_382_672, w_335_006, w_158_257);
  not1 I382_678(w_382_678, w_305_006);
  and2 I383_097(w_383_097, w_076_103, w_003_193);
  or2  I383_133(w_383_133, w_009_055, w_022_186);
  not1 I383_187(w_383_187, w_078_434);
  or2  I383_219(w_383_219, w_014_225, w_205_699);
  and2 I383_235(w_383_235, w_133_138, w_248_161);
  not1 I383_377(w_383_377, w_014_822);
  not1 I384_1443(w_384_1443, w_345_1481);
  and2 I385_227(w_385_227, w_287_027, w_368_653);
  not1 I385_326(w_385_326, w_264_337);
  nand2 I386_011(w_386_011, w_299_1221, w_319_307);
  and2 I386_236(w_386_236, w_012_252, w_006_262);
  and2 I387_317(w_387_317, w_156_132, w_308_457);
  or2  I387_619(w_387_619, w_325_1102, w_305_012);
  nand2 I387_691(w_387_691, w_163_1558, w_031_724);
  nand2 I387_720(w_387_720, w_171_858, w_311_641);
  not1 I387_967(w_387_967, w_153_1254);
  nand2 I388_219(w_388_219, w_173_1074, w_147_049);
  or2  I388_339(w_388_339, w_364_722, w_274_034);
  and2 I388_630(w_388_630, w_090_919, w_010_325);
  nand2 I388_751(w_388_751, w_281_595, w_362_337);
  nand2 I388_936(w_388_936, w_166_227, w_370_077);
  or2  I389_671(w_389_671, w_244_200, w_132_046);
  or2  I389_787(w_389_787, w_256_362, w_386_236);
  not1 I389_1252(w_389_1252, w_035_1053);
  and2 I389_1431(w_389_1431, w_292_708, w_125_545);
  not1 I389_1549(w_389_1549, w_129_877);
  and2 I389_1637(w_389_1637, w_233_219, w_022_223);
  nand2 I390_195(w_390_195, w_264_556, w_109_032);
  nand2 I390_434(w_390_434, w_365_216, w_120_000);
  or2  I390_717(w_390_717, w_062_064, w_044_314);
  not1 I391_015(w_391_015, w_151_1109);
  nand2 I391_048(w_391_048, w_202_727, w_159_974);
  or2  I392_480(w_392_480, w_240_427, w_194_257);
  nand2 I392_598(w_392_598, w_149_590, w_310_189);
  nand2 I392_982(w_392_982, w_388_630, w_368_156);
  and2 I392_1327(w_392_1327, w_183_1551, w_005_1252);
  not1 I392_1798(w_392_1798, w_207_1006);
  or2  I393_523(w_393_523, w_152_430, w_138_064);
  or2  I394_008(w_394_008, w_075_001, w_094_005);
  and2 I394_013(w_394_013, w_307_013, w_266_233);
  and2 I394_030(w_394_030, w_310_505, w_054_313);
  and2 I394_037(w_394_037, w_094_055, w_296_305);
  nand2 I395_657(w_395_657, w_131_405, w_299_1159);
  nand2 I395_966(w_395_966, w_322_112, w_369_228);
  not1 I396_001(w_396_001, w_213_743);
  and2 I396_254(w_396_254, w_283_1561, w_067_292);
  or2  I396_282(w_396_282, w_214_078, w_186_180);
  and2 I396_560(w_396_560, w_238_062, w_353_448);
  not1 I397_455(w_397_455, w_380_434);
  not1 I397_673(w_397_673, w_129_608);
  or2  I397_1350(w_397_1350, w_273_376, w_373_1442);
  nand2 I397_1463(w_397_1463, w_341_141, w_152_120);
  or2  I398_086(w_398_086, w_139_070, w_318_012);
  not1 I398_235(w_398_235, w_179_807);
  nand2 I398_258(w_398_258, w_317_1030, w_196_282);
  not1 I398_887(w_398_887, w_329_059);
  nand2 I398_1205(w_398_1205, w_179_122, w_100_1813);
  or2  I398_1585(w_398_1585, w_256_894, w_080_030);
  or2  I399_076(w_399_076, w_024_212, w_110_026);
  nand2 I399_191(w_399_191, w_021_143, w_317_1547);
  nand2 I399_563(w_399_563, w_327_1107, w_312_514);
  and2 I399_1417(w_399_1417, w_192_428, w_384_1443);
  not1 I399_1787(w_399_1789, w_399_1788);
  not1 I399_1788(w_399_1790, w_399_1789);
  and2 I399_1789(w_399_1791, w_399_1806, w_399_1790);
  not1 I399_1790(w_399_1792, w_399_1791);
  or2  I399_1791(w_399_1793, w_399_1792, w_079_747);
  not1 I399_1792(w_399_1794, w_399_1793);
  or2  I399_1793(w_399_1795, w_399_1794, w_368_455);
  not1 I399_1794(w_399_1796, w_399_1795);
  not1 I399_1795(w_399_1797, w_399_1796);
  not1 I399_1796(w_399_1798, w_399_1797);
  and2 I399_1797(w_399_1788, w_399_1798, w_141_123);
  not1 I399_1798(w_399_1803, w_399_1802);
  not1 I399_1799(w_399_1804, w_399_1803);
  not1 I399_1800(w_399_1802, w_399_1791);
  and2 I399_1801(w_399_1806, w_250_208, w_399_1804);
  or2  I400_067(w_400_067, w_139_697, w_059_214);
  nand2 I400_224(w_400_224, w_145_040, w_086_780);
  and2 I401_063(w_401_063, w_382_678, w_087_242);
  nand2 I401_383(w_401_383, w_029_719, w_087_1123);
  not1 I401_517(w_401_517, w_275_427);
  not1 I401_544(w_401_544, w_170_1654);
  and2 I402_176(w_402_176, w_265_1117, w_292_732);
  nand2 I402_569(w_402_569, w_383_187, w_094_100);
  not1 I402_632(w_402_632, w_011_111);
  and2 I402_872(w_402_872, w_368_783, w_173_1159);
  or2  I402_998(w_402_998, w_339_439, w_034_276);
  nand2 I403_004(w_403_004, w_345_1240, w_101_221);
  and2 I403_097(w_403_097, w_196_440, w_368_1314);
  and2 I403_146(w_403_146, w_009_063, w_021_086);
  not1 I403_215(w_403_215, w_293_212);
  and2 I403_223(w_403_223, w_383_235, w_311_245);
  and2 I404_052(w_404_052, w_101_670, w_189_011);
  or2  I404_266(w_404_266, w_025_1442, w_370_616);
  not1 I404_800(w_404_800, w_271_982);
  nand2 I405_122(w_405_122, w_214_697, w_146_075);
  not1 I405_171(w_405_171, w_173_079);
  nand2 I405_284(w_405_284, w_397_455, w_065_003);
  nand2 I406_175(w_406_175, w_104_1248, w_097_469);
  and2 I406_471(w_406_471, w_143_109, w_151_834);
  or2  I406_554(w_406_554, w_072_007, w_061_367);
  and2 I406_677(w_406_677, w_331_107, w_142_170);
  nand2 I406_835(w_406_835, w_108_467, w_195_1485);
  nand2 I406_870(w_406_870, w_364_233, w_161_171);
  and2 I406_964(w_406_964, w_134_1230, w_170_167);
  nand2 I407_014(w_407_014, w_330_753, w_056_1388);
  and2 I407_182(w_407_182, w_068_086, w_355_291);
  or2  I408_005(w_408_005, w_028_638, w_398_235);
  or2  I408_011(w_408_011, w_119_1518, w_023_1163);
  not1 I408_015(w_408_015, w_369_1046);
  not1 I408_017(w_408_017, w_214_558);
  nand2 I409_138(w_409_138, w_283_224, w_394_008);
  and2 I409_623(w_409_623, w_367_489, w_057_1156);
  and2 I409_732(w_409_732, w_289_921, w_183_054);
  nand2 I409_773(w_409_773, w_279_187, w_212_066);
  nand2 I410_008(w_410_008, w_359_1125, w_106_370);
  not1 I410_069(w_410_069, w_295_546);
  nand2 I410_103(w_410_103, w_291_244, w_132_068);
  not1 I410_111(w_410_111, w_304_1575);
  not1 I410_164(w_410_164, w_118_152);
  or2  I411_668(w_411_668, w_312_425, w_408_015);
  not1 I411_987(w_411_987, w_183_035);
  and2 I411_1244(w_411_1244, w_156_558, w_093_052);
  or2  I411_1382(w_411_1382, w_116_1531, w_391_015);
  and2 I411_1447(w_411_1447, w_194_643, w_296_801);
  not1 I412_000(w_412_000, w_117_499);
  or2  I412_028(w_412_028, w_123_1252, w_409_623);
  or2  I412_161(w_412_161, w_252_500, w_325_1468);
  not1 I412_437(w_412_437, w_178_032);
  not1 I413_194(w_413_194, w_069_980);
  or2  I414_110(w_414_110, w_245_1128, w_191_098);
  or2  I415_024(w_415_024, w_091_081, w_016_020);
  nand2 I415_058(w_415_058, w_159_215, w_283_1042);
  or2  I415_207(w_415_207, w_357_141, w_201_166);
  not1 I416_198(w_416_198, w_305_008);
  or2  I416_298(w_416_298, w_200_406, w_167_028);
  and2 I416_307(w_416_307, w_111_712, w_249_765);
  and2 I416_364(w_416_364, w_164_761, w_104_1647);
  not1 I416_432(w_416_432, w_354_1261);
  and2 I416_600(w_416_600, w_108_374, w_306_427);
  nand2 I416_1113(w_416_1113, w_003_139, w_100_579);
  and2 I417_017(w_417_017, w_381_839, w_268_361);
  nand2 I417_456(w_417_456, w_032_077, w_273_075);
  or2  I418_170(w_418_170, w_273_623, w_299_340);
  not1 I418_475(w_418_475, w_112_631);
  nand2 I418_479(w_418_479, w_163_1548, w_344_150);
  not1 I418_673(w_418_673, w_017_1131);
  not1 I418_1325(w_418_1325, w_234_664);
  or2  I418_1382(w_418_1382, w_357_026, w_240_590);
  not1 I419_069(w_419_069, w_169_372);
  not1 I419_087(w_419_087, w_235_573);
  or2  I419_178(w_419_178, w_208_175, w_154_098);
  or2  I420_832(w_420_832, w_360_762, w_410_111);
  and2 I420_1439(w_420_1439, w_113_575, w_264_430);
  nand2 I421_031(w_421_031, w_186_119, w_013_274);
  or2  I421_096(w_421_096, w_360_496, w_180_529);
  nand2 I421_143(w_421_143, w_027_351, w_232_002);
  not1 I421_154(w_421_154, w_398_887);
  not1 I421_269(w_421_269, w_060_095);
  or2  I421_275(w_421_275, w_289_377, w_412_161);
  nand2 I421_311(w_421_311, w_238_332, w_051_960);
  not1 I422_251(w_422_251, w_050_875);
  nand2 I422_306(w_422_306, w_389_671, w_234_1004);
  or2  I422_351(w_422_351, w_238_143, w_084_197);
  not1 I422_384(w_422_384, w_289_398);
  not1 I422_579(w_422_579, w_332_617);
  or2  I423_080(w_423_080, w_207_587, w_190_1780);
  not1 I423_206(w_423_206, w_323_111);
  not1 I424_002(w_424_002, w_113_007);
  or2  I424_010(w_424_010, w_135_078, w_265_1327);
  not1 I424_016(w_424_016, w_299_086);
  or2  I424_021(w_424_021, w_019_773, w_212_009);
  and2 I424_022(w_424_022, w_405_171, w_030_318);
  and2 I424_025(w_424_025, w_106_1199, w_062_878);
  nand2 I425_174(w_425_174, w_145_009, w_075_105);
  and2 I425_247(w_425_247, w_389_1431, w_195_086);
  and2 I426_621(w_426_621, w_085_676, w_144_1212);
  not1 I427_021(w_427_021, w_064_096);
  and2 I427_055(w_427_055, w_159_596, w_182_066);
  and2 I427_082(w_427_082, w_084_139, w_122_127);
  not1 I427_169(w_427_169, w_048_627);
  and2 I427_172(w_427_172, w_378_048, w_318_277);
  not1 I427_245(w_427_245, w_242_030);
  not1 I427_257(w_427_257, w_046_062);
  and2 I428_864(w_428_864, w_305_011, w_130_648);
  nand2 I429_200(w_429_200, w_278_772, w_104_128);
  or2  I429_1594(w_429_1594, w_338_073, w_322_143);
  or2  I430_014(w_430_014, w_353_691, w_168_649);
  not1 I430_067(w_430_067, w_378_597);
  not1 I430_069(w_430_069, w_351_021);
  or2  I430_088(w_430_088, w_086_755, w_325_661);
  nand2 I430_130(w_430_130, w_288_272, w_128_246);
  or2  I431_218(w_431_218, w_197_493, w_084_058);
  and2 I431_239(w_431_239, w_285_021, w_092_204);
  and2 I431_1031(w_431_1031, w_223_721, w_111_352);
  and2 I431_1266(w_431_1266, w_283_357, w_230_132);
  or2  I432_171(w_432_171, w_108_705, w_355_155);
  not1 I432_725(w_432_727, w_432_726);
  or2  I432_726(w_432_728, w_170_196, w_432_727);
  not1 I432_727(w_432_729, w_432_728);
  not1 I432_728(w_432_730, w_432_729);
  and2 I432_729(w_432_731, w_336_663, w_432_730);
  nand2 I432_730(w_432_726, w_432_731, w_432_741);
  or2  I432_731(w_432_736, w_059_353, w_432_735);
  and2 I432_732(w_432_737, w_144_1040, w_432_736);
  and2 I432_733(w_432_738, w_068_126, w_432_737);
  not1 I432_734(w_432_739, w_432_738);
  not1 I432_735(w_432_735, w_432_726);
  and2 I432_736(w_432_741, w_394_013, w_432_739);
  and2 I433_070(w_433_070, w_087_1021, w_392_1798);
  not1 I433_394(w_433_394, w_081_311);
  and2 I433_430(w_433_430, w_248_450, w_354_278);
  nand2 I433_560(w_433_560, w_269_1979, w_294_087);
  nand2 I433_592(w_433_592, w_409_732, w_252_160);
  or2  I433_631(w_433_631, w_430_069, w_123_590);
  and2 I433_824(w_433_824, w_115_508, w_004_134);
  not1 I434_621(w_434_621, w_363_598);
  not1 I434_633(w_434_633, w_426_621);
  nand2 I435_916(w_435_916, w_107_398, w_276_176);
  nand2 I436_667(w_436_667, w_343_894, w_371_548);
  not1 I436_1391(w_436_1391, w_433_430);
  and2 I436_1601(w_436_1601, w_278_1377, w_111_122);
  and2 I437_1451(w_437_1451, w_355_018, w_255_206);
  or2  I437_1574(w_437_1574, w_086_178, w_217_031);
  and2 I438_1586(w_438_1586, w_163_015, w_234_048);
  nand2 I439_508(w_439_508, w_239_061, w_120_057);
  not1 I439_531(w_439_531, w_141_297);
  not1 I440_591(w_440_591, w_418_170);
  and2 I440_709(w_440_709, w_064_636, w_350_527);
  not1 I440_814(w_440_814, w_083_019);
  nand2 I440_896(w_440_896, w_074_115, w_371_343);
  or2  I441_128(w_441_128, w_059_246, w_423_080);
  nand2 I441_750(w_441_750, w_059_179, w_406_175);
  not1 I441_948(w_441_948, w_124_260);
  not1 I442_118(w_442_118, w_202_1120);
  not1 I442_759(w_442_759, w_237_519);
  nand2 I442_803(w_442_803, w_233_120, w_207_1116);
  not1 I442_1693(w_442_1693, w_143_988);
  and2 I443_305(w_443_305, w_238_509, w_389_1549);
  nand2 I443_369(w_443_369, w_431_1266, w_100_021);
  and2 I443_718(w_443_718, w_054_065, w_141_073);
  or2  I444_085(w_444_085, w_075_109, w_183_1795);
  not1 I444_113(w_444_113, w_265_1397);
  or2  I445_301(w_445_301, w_174_624, w_372_317);
  not1 I445_361(w_445_361, w_387_619);
  nand2 I445_394(w_445_394, w_299_1560, w_334_566);
  and2 I446_046(w_446_046, w_154_136, w_408_017);
  and2 I446_247(w_446_247, w_069_1270, w_031_248);
  nand2 I446_536(w_446_536, w_130_700, w_113_372);
  and2 I446_605(w_446_605, w_175_088, w_208_702);
  and2 I446_698(w_446_698, w_192_346, w_358_675);
  not1 I446_722(w_446_722, w_157_993);
  and2 I446_752(w_446_752, w_399_076, w_163_1642);
  or2  I447_169(w_447_169, w_442_803, w_410_069);
  and2 I448_252(w_448_252, w_306_1282, w_191_445);
  or2  I448_423(w_448_423, w_283_1724, w_235_757);
  not1 I449_347(w_449_347, w_141_180);
  or2  I449_402(w_449_402, w_082_431, w_159_802);
  nand2 I449_1041(w_449_1041, w_195_1391, w_175_102);
  nand2 I451_401(w_451_401, w_268_1259, w_284_147);
  or2  I451_616(w_451_616, w_362_1655, w_121_216);
  and2 I451_632(w_451_632, w_062_105, w_020_154);
  or2  I452_108(w_452_108, w_210_367, w_031_733);
  not1 I452_176(w_452_176, w_007_1379);
  not1 I452_289(w_452_289, w_282_537);
  or2  I452_775(w_452_775, w_075_116, w_264_021);
  nand2 I453_073(w_453_073, w_226_239, w_084_304);
  and2 I453_109(w_453_109, w_047_434, w_346_679);
  not1 I453_115(w_453_115, w_008_254);
  nand2 I453_196(w_453_196, w_339_235, w_421_096);
  nand2 I454_021(w_454_021, w_370_890, w_138_013);
  nand2 I454_025(w_454_025, w_406_677, w_201_230);
  or2  I454_043(w_454_043, w_250_207, w_007_752);
  or2  I454_142(w_454_142, w_324_469, w_237_819);
  nand2 I454_260(w_454_260, w_196_289, w_194_705);
  not1 I456_283(w_456_283, w_415_024);
  not1 I456_442(w_456_442, w_278_946);
  or2  I456_731(w_456_731, w_363_803, w_062_544);
  nand2 I456_769(w_456_769, w_328_008, w_392_982);
  not1 I456_979(w_456_979, w_452_176);
  nand2 I457_975(w_457_975, w_380_321, w_416_432);
  nand2 I457_1220(w_457_1222, w_034_121, w_457_1221);
  not1 I457_1221(w_457_1223, w_457_1222);
  not1 I457_1222(w_457_1224, w_457_1223);
  nand2 I457_1223(w_457_1225, w_013_110, w_457_1224);
  not1 I457_1224(w_457_1226, w_457_1225);
  nand2 I457_1225(w_457_1221, w_457_1226, w_254_114);
  nand2 I458_073(w_458_073, w_353_1174, w_170_991);
  and2 I458_412(w_458_412, w_229_1356, w_390_717);
  nand2 I458_1066(w_458_1066, w_187_394, w_454_260);
  or2  I459_383(w_459_383, w_255_196, w_032_037);
  not1 I459_833(w_459_833, w_194_103);
  and2 I460_906(w_460_906, w_440_896, w_331_899);
  and2 I460_1204(w_460_1204, w_404_800, w_279_250);
  and2 I461_047(w_461_047, w_069_350, w_071_028);
  or2  I461_171(w_461_171, w_444_085, w_218_058);
  and2 I461_280(w_461_280, w_177_1547, w_019_1031);
  and2 I461_310(w_461_310, w_178_285, w_412_000);
  or2  I461_319(w_461_319, w_200_293, w_446_046);
  not1 I461_651(w_461_651, w_116_912);
  or2  I461_696(w_461_696, w_038_260, w_256_557);
  nand2 I462_021(w_462_021, w_274_044, w_187_270);
  or2  I462_025(w_462_025, w_020_1191, w_223_1210);
  not1 I462_134(w_462_134, w_276_078);
  and2 I463_044(w_463_044, w_402_632, w_353_531);
  or2  I463_144(w_463_144, w_324_105, w_006_084);
  and2 I463_172(w_463_172, w_194_580, w_338_1654);
  or2  I463_340(w_463_340, w_403_215, w_193_336);
  nand2 I463_433(w_463_433, w_150_493, w_067_961);
  or2  I463_473(w_463_473, w_256_957, w_065_005);
  not1 I464_379(w_464_379, w_081_447);
  and2 I465_050(w_465_050, w_318_192, w_454_142);
  or2  I465_943(w_465_943, w_026_1371, w_007_264);
  and2 I466_005(w_466_005, w_042_127, w_354_064);
  not1 I466_103(w_466_103, w_134_012);
  not1 I466_234(w_466_234, w_015_066);
  or2  I466_271(w_466_271, w_046_147, w_106_158);
  and2 I467_390(w_467_390, w_247_759, w_197_073);
  nand2 I467_689(w_467_689, w_199_005, w_068_169);
  and2 I467_1137(w_467_1137, w_174_078, w_437_1451);
  or2  I468_214(w_468_214, w_026_1107, w_441_948);
  nand2 I468_249(w_468_249, w_199_1092, w_099_224);
  and2 I468_253(w_468_253, w_059_489, w_325_1228);
  or2  I469_046(w_469_046, w_057_487, w_381_634);
  nand2 I469_351(w_469_351, w_176_823, w_303_045);
  nand2 I469_529(w_469_529, w_162_894, w_323_288);
  and2 I470_456(w_470_456, w_231_482, w_184_004);
  not1 I470_1212(w_470_1212, w_153_356);
  not1 I471_265(w_471_265, w_202_090);
  and2 I471_359(w_471_359, w_224_249, w_306_282);
  not1 I471_553(w_471_553, w_120_032);
  and2 I473_022(w_473_022, w_313_028, w_268_033);
  or2  I473_245(w_473_245, w_070_051, w_214_392);
  not1 I473_1043(w_473_1043, w_416_298);
  or2  I474_300(w_474_300, w_313_005, w_322_1155);
  nand2 I474_412(w_474_412, w_049_515, w_066_863);
  and2 I475_095(w_475_095, w_213_041, w_132_033);
  not1 I475_175(w_475_175, w_286_239);
  not1 I475_219(w_475_219, w_243_1147);
  nand2 I476_073(w_476_073, w_433_824, w_336_181);
  and2 I476_096(w_476_096, w_166_104, w_418_1382);
  or2  I476_191(w_476_191, w_141_261, w_416_307);
  not1 I476_312(w_476_312, w_152_039);
  not1 I476_313(w_476_313, w_124_165);
  and2 I476_379(w_476_379, w_329_203, w_307_243);
  or2  I476_389(w_476_389, w_237_042, w_411_1447);
  nand2 I477_023(w_477_023, w_327_428, w_359_131);
  not1 I477_098(w_477_098, w_234_1138);
  and2 I477_104(w_477_104, w_072_058, w_451_616);
  not1 I478_293(w_478_293, w_058_212);
  not1 I478_367(w_478_367, w_125_1126);
  or2  I478_665(w_478_665, w_269_1751, w_045_1704);
  and2 I478_815(w_478_815, w_420_832, w_251_157);
  and2 I478_1092(w_478_1092, w_016_018, w_292_019);
  not1 I478_1191(w_478_1191, w_475_219);
  and2 I478_1446(w_478_1446, w_421_031, w_422_579);
  not1 I479_615(w_479_615, w_169_408);
  or2  I479_638(w_479_638, w_120_117, w_347_1311);
  not1 I479_643(w_479_643, w_298_578);
  nand2 I479_694(w_479_694, w_275_392, w_072_055);
  not1 I479_1024(w_479_1024, w_284_047);
  not1 I479_1741(w_479_1741, w_118_710);
  nand2 I480_021(w_480_021, w_041_073, w_335_072);
  and2 I480_062(w_480_062, w_473_245, w_339_524);
  or2  I481_093(w_481_093, w_419_178, w_300_014);
  not1 I481_1485(w_481_1485, w_187_263);
  or2  I482_410(w_482_410, w_449_402, w_222_1038);
  and2 I482_839(w_482_839, w_453_109, w_088_815);
  or2  I483_094(w_483_094, w_226_639, w_189_010);
  not1 I483_314(w_483_314, w_364_1423);
  and2 I483_425(w_483_425, w_204_1212, w_020_304);
  nand2 I484_010(w_484_010, w_140_948, w_101_523);
  nand2 I484_362(w_484_362, w_227_104, w_203_650);
  not1 I484_491(w_484_493, w_484_492);
  not1 I484_492(w_484_494, w_484_493);
  or2  I484_493(w_484_492, w_484_494, w_484_509);
  not1 I484_494(w_484_499, w_484_498);
  or2  I484_495(w_484_500, w_484_499, w_327_290);
  and2 I484_496(w_484_501, w_194_552, w_484_500);
  not1 I484_497(w_484_502, w_484_501);
  nand2 I484_498(w_484_503, w_484_502, w_033_801);
  or2  I484_499(w_484_504, w_484_503, w_166_531);
  nand2 I484_500(w_484_505, w_211_336, w_484_504);
  and2 I484_501(w_484_506, w_484_505, w_053_029);
  not1 I484_502(w_484_507, w_484_506);
  not1 I484_503(w_484_498, w_484_492);
  and2 I484_504(w_484_509, w_183_998, w_484_507);
  nand2 I485_176(w_485_176, w_271_200, w_111_376);
  not1 I487_032(w_487_032, w_093_001);
  or2  I487_525(w_487_525, w_454_021, w_418_479);
  nand2 I487_617(w_487_617, w_132_032, w_115_627);
  and2 I487_790(w_487_790, w_412_437, w_403_146);
  or2  I487_1069(w_487_1069, w_398_258, w_035_643);
  not1 I487_1147(w_487_1147, w_168_320);
  not1 I488_278(w_488_278, w_321_196);
  not1 I488_641(w_488_641, w_418_475);
  and2 I488_908(w_488_908, w_194_074, w_339_121);
  not1 I488_978(w_488_978, w_279_570);
  not1 I489_036(w_489_036, w_180_040);
  or2  I489_1324(w_489_1324, w_475_175, w_176_1462);
  or2  I489_1344(w_489_1344, w_022_418, w_150_006);
  nand2 I490_288(w_490_288, w_080_067, w_285_142);
  or2  I490_1421(w_490_1421, w_294_314, w_081_242);
  not1 I491_048(w_491_048, w_463_340);
  and2 I491_164(w_491_164, w_206_165, w_016_027);
  nand2 I492_043(w_492_043, w_049_489, w_232_388);
  nand2 I492_085(w_492_085, w_350_207, w_210_428);
  nand2 I492_086(w_492_086, w_005_255, w_092_616);
  not1 I492_128(w_492_128, w_251_169);
  or2  I493_062(w_493_062, w_164_565, w_171_539);
  or2  I493_157(w_493_157, w_299_308, w_060_077);
  nand2 I493_225(w_493_225, w_479_638, w_208_912);
  or2  I493_430(w_493_430, w_376_750, w_116_390);
  and2 I493_441(w_493_441, w_250_183, w_225_186);
  nand2 I493_571(w_493_573, w_493_589, w_493_572);
  nand2 I493_572(w_493_574, w_493_573, w_262_184);
  not1 I493_573(w_493_575, w_493_574);
  nand2 I493_574(w_493_576, w_349_104, w_493_575);
  not1 I493_575(w_493_577, w_493_576);
  not1 I493_576(w_493_578, w_493_577);
  nand2 I493_577(w_493_572, w_493_578, w_476_312);
  and2 I493_578(w_493_583, w_493_582, w_310_332);
  not1 I493_579(w_493_584, w_493_583);
  not1 I493_580(w_493_585, w_493_584);
  and2 I493_581(w_493_586, w_138_041, w_493_585);
  and2 I493_582(w_493_587, w_493_586, w_180_422);
  not1 I493_583(w_493_582, w_493_573);
  and2 I493_584(w_493_589, w_287_352, w_493_587);
  nand2 I494_945(w_494_945, w_311_135, w_404_052);
  nand2 I494_1233(w_494_1233, w_150_016, w_223_1368);
  and2 I494_1930(w_494_1932, w_494_1931, w_344_117);
  nand2 I494_1931(w_494_1933, w_461_319, w_494_1932);
  and2 I494_1932(w_494_1934, w_465_943, w_494_1933);
  and2 I494_1933(w_494_1935, w_171_152, w_494_1934);
  and2 I494_1934(w_494_1936, w_016_025, w_494_1935);
  not1 I494_1935(w_494_1931, w_494_1936);
  nand2 I495_1004(w_495_1004, w_427_257, w_339_405);
  or2  I495_1084(w_495_1084, w_133_737, w_353_985);
  not1 I496_101(w_496_101, w_061_260);
  and2 I496_495(w_496_495, w_487_617, w_350_529);
  and2 I496_628(w_496_628, w_202_1580, w_222_1290);
  nand2 I496_797(w_496_797, w_493_062, w_494_1233);
  and2 I496_959(w_496_959, w_016_016, w_174_370);
  not1 I496_1215(w_496_1215, w_402_872);
  and2 I497_331(w_497_331, w_372_366, w_184_006);
  and2 I497_364(w_497_364, w_308_281, w_278_723);
  nand2 I497_391(w_497_391, w_105_126, w_425_174);
  not1 I498_402(w_498_402, w_202_372);
  nand2 I498_507(w_498_507, w_321_129, w_019_436);
  or2  I498_636(w_498_636, w_156_038, w_312_146);
  or2  I499_181(w_499_181, w_370_066, w_019_343);
  nand2 I499_371(w_499_371, w_233_056, w_223_022);
  and2 I499_436(w_499_436, w_275_027, w_103_237);
  not1 I499_1419(w_499_1419, w_453_115);
  nand2 I499_1719(w_499_1719, w_200_051, w_062_140);
  nand2 I500_004(w_500_004, w_210_375, w_037_777);
  nand2 I500_891(w_500_891, w_008_070, w_106_336);
  and2 I500_1299(w_500_1299, w_491_164, w_139_1525);
  nand2 I501_352(w_501_352, w_294_564, w_405_122);
  not1 I502_002(w_502_002, w_453_073);
  not1 I502_250(w_502_250, w_106_252);
  not1 I502_289(w_502_289, w_371_710);
  not1 I503_023(w_503_023, w_036_696);
  nand2 I503_261(w_503_261, w_133_392, w_402_176);
  not1 I503_299(w_503_299, w_282_1923);
  or2  I503_404(w_503_404, w_454_025, w_421_275);
  or2  I503_694(w_503_694, w_383_097, w_260_048);
  and2 I504_065(w_504_065, w_422_384, w_262_119);
  or2  I504_152(w_504_152, w_034_104, w_001_1030);
  not1 I504_314(w_504_314, w_334_597);
  and2 I504_564(w_504_564, w_136_661, w_305_012);
  not1 I505_342(w_505_342, w_098_432);
  nand2 I505_916(w_505_916, w_117_559, w_500_004);
  and2 I505_1503(w_505_1503, w_145_017, w_456_979);
  and2 I505_1562(w_505_1562, w_293_608, w_047_577);
  not1 I506_135(w_506_135, w_312_218);
  nand2 I506_138(w_506_138, w_344_207, w_105_1716);
  nand2 I506_472(w_506_472, w_353_380, w_479_694);
  and2 I507_047(w_507_047, w_191_1390, w_289_856);
  not1 I507_110(w_507_110, w_019_784);
  or2  I508_018(w_508_018, w_346_341, w_332_1090);
  or2  I509_068(w_509_068, w_029_474, w_222_642);
  or2  I509_110(w_509_110, w_191_626, w_023_622);
  and2 I509_148(w_509_148, w_126_004, w_440_591);
  or2  I509_294(w_509_294, w_084_050, w_320_632);
  and2 I509_322(w_509_322, w_505_916, w_505_1562);
  and2 I509_386(w_509_386, w_281_044, w_244_535);
  and2 I510_051(w_510_051, w_490_288, w_020_1263);
  or2  I510_177(w_510_177, w_085_081, w_461_651);
  and2 I510_180(w_510_180, w_499_371, w_298_1342);
  not1 I510_260(w_510_260, w_169_1109);
  and2 I510_261(w_510_261, w_003_062, w_284_1406);
  not1 I512_268(w_512_268, w_283_1343);
  or2  I512_374(w_512_374, w_254_015, w_445_394);
  not1 I512_679(w_512_679, w_363_075);
  not1 I512_823(w_512_823, w_480_021);
  or2  I512_1078(w_512_1078, w_206_918, w_158_099);
  or2  I513_409(w_513_409, w_049_336, w_107_488);
  and2 I513_1030(w_513_1030, w_504_065, w_385_326);
  nand2 I514_053(w_514_053, w_070_231, w_134_150);
  nand2 I514_848(w_514_848, w_093_004, w_477_023);
  nand2 I514_955(w_514_955, w_344_052, w_230_121);
  or2  I514_1099(w_514_1099, w_302_321, w_307_203);
  nand2 I514_1390(w_514_1390, w_387_691, w_165_227);
  or2  I515_094(w_515_094, w_270_663, w_427_245);
  or2  I515_186(w_515_186, w_092_164, w_470_1212);
  or2  I515_456(w_515_456, w_509_294, w_487_525);
  not1 I515_657(w_515_657, w_393_523);
  and2 I515_679(w_515_679, w_191_076, w_223_179);
  or2  I516_317(w_516_317, w_052_1038, w_115_579);
  not1 I516_699(w_516_699, w_166_656);
  nand2 I517_039(w_517_039, w_118_233, w_274_015);
  nand2 I518_204(w_518_204, w_346_640, w_424_010);
  or2  I519_189(w_519_189, w_308_778, w_314_499);
  not1 I520_598(w_520_598, w_264_435);
  or2  I520_667(w_520_667, w_006_195, w_249_066);
  and2 I520_1416(w_520_1416, w_451_401, w_456_442);
  or2  I521_852(w_521_852, w_116_1491, w_265_456);
  or2  I522_090(w_522_090, w_119_924, w_372_428);
  and2 I523_021(w_523_021, w_452_289, w_372_404);
  or2  I523_688(w_523_688, w_088_1192, w_016_022);
  or2  I524_121(w_524_121, w_462_021, w_119_642);
  or2  I524_464(w_524_464, w_479_615, w_425_247);
  or2  I524_1502(w_524_1502, w_171_101, w_355_089);
  or2  I524_1505(w_524_1505, w_222_633, w_293_660);
  and2 I525_175(w_525_175, w_304_1593, w_302_660);
  or2  I525_366(w_525_366, w_394_037, w_033_093);
  or2  I525_1141(w_525_1141, w_086_1118, w_301_1829);
  nand2 I525_1399(w_525_1399, w_202_1780, w_308_1148);
  nand2 I528_041(w_528_041, w_096_176, w_006_178);
  or2  I528_110(w_528_110, w_192_486, w_491_048);
  not1 I528_145(w_528_145, w_002_378);
  nand2 I529_180(w_529_180, w_337_158, w_410_164);
  nand2 I530_1263(w_530_1263, w_154_073, w_132_039);
  not1 I530_1605(w_530_1605, w_466_234);
  nand2 I531_121(w_531_121, w_473_022, w_446_698);
  and2 I531_628(w_531_628, w_069_001, w_002_428);
  or2  I531_1377(w_531_1379, w_531_1378, w_398_1585);
  nand2 I531_1378(w_531_1380, w_531_1379, w_468_253);
  not1 I531_1379(w_531_1381, w_531_1380);
  not1 I531_1380(w_531_1382, w_531_1381);
  not1 I531_1381(w_531_1383, w_531_1382);
  nand2 I531_1382(w_531_1384, w_531_1383, w_503_404);
  or2  I531_1383(w_531_1385, w_531_1384, w_350_314);
  not1 I531_1384(w_531_1386, w_531_1385);
  not1 I531_1385(w_531_1387, w_531_1386);
  nand2 I531_1386(w_531_1388, w_531_1397, w_531_1387);
  and2 I531_1387(w_531_1378, w_531_1388, w_108_717);
  not1 I531_1388(w_531_1393, w_531_1392);
  nand2 I531_1389(w_531_1394, w_386_011, w_531_1393);
  not1 I531_1390(w_531_1395, w_531_1394);
  not1 I531_1391(w_531_1392, w_531_1388);
  and2 I531_1392(w_531_1397, w_207_479, w_531_1395);
  not1 I532_271(w_532_271, w_157_762);
  and2 I532_410(w_532_410, w_323_386, w_137_239);
  and2 I534_014(w_534_014, w_113_097, w_323_446);
  and2 I534_1008(w_534_1008, w_242_046, w_421_154);
  or2  I534_1231(w_534_1231, w_053_048, w_207_1454);
  not1 I536_150(w_536_150, w_411_1382);
  nand2 I537_388(w_537_388, w_030_561, w_117_589);
  nand2 I537_615(w_537_615, w_084_334, w_086_1493);
  nand2 I538_357(w_538_357, w_313_000, w_358_471);
  nand2 I538_363(w_538_363, w_234_587, w_351_000);
  and2 I538_713(w_538_713, w_276_091, w_107_296);
  nand2 I538_864(w_538_864, w_229_1499, w_042_105);
  not1 I539_231(w_539_231, w_062_1111);
  nand2 I540_182(w_540_182, w_015_007, w_180_482);
  or2  I540_326(w_540_326, w_330_731, w_141_636);
  not1 I540_341(w_540_341, w_331_838);
  nand2 I541_073(w_541_073, w_406_835, w_285_671);
  not1 I542_089(w_542_089, w_085_153);
  and2 I542_308(w_542_308, w_288_036, w_169_1242);
  or2  I543_374(w_543_374, w_108_731, w_043_093);
  and2 I543_594(w_543_594, w_108_398, w_457_975);
  not1 I543_740(w_543_740, w_293_875);
  or2  I544_028(w_544_028, w_138_151, w_383_133);
  and2 I544_040(w_544_040, w_539_231, w_392_598);
  and2 I544_081(w_544_081, w_265_476, w_263_558);
  and2 I544_100(w_544_100, w_063_1100, w_191_1190);
  or2  I545_1135(w_545_1135, w_315_234, w_125_252);
  not1 I545_1157(w_545_1157, w_107_971);
  and2 I546_065(w_546_065, w_072_001, w_316_510);
  or2  I546_078(w_546_078, w_273_751, w_496_628);
  or2  I546_258(w_546_258, w_382_653, w_168_225);
  not1 I546_1098(w_546_1098, w_389_787);
  and2 I547_082(w_547_082, w_385_227, w_438_1586);
  or2  I547_437(w_547_437, w_088_552, w_370_067);
  nand2 I548_325(w_548_325, w_053_031, w_292_145);
  and2 I548_356(w_548_356, w_403_004, w_329_262);
  or2  I548_509(w_548_509, w_257_1369, w_484_010);
  not1 I548_636(w_548_636, w_515_657);
  not1 I548_843(w_548_843, w_004_028);
  nand2 I548_923(w_548_923, w_458_073, w_528_041);
  nand2 I549_164(w_549_164, w_062_605, w_075_096);
  and2 I549_222(w_549_222, w_512_374, w_307_008);
  or2  I549_244(w_549_244, w_349_052, w_151_587);
  and2 I549_284(w_549_284, w_120_002, w_365_858);
  not1 I549_352(w_549_352, w_168_259);
  and2 I550_785(w_550_785, w_151_380, w_281_393);
  and2 I551_082(w_551_082, w_542_308, w_119_798);
  not1 I551_271(w_551_271, w_538_363);
  and2 I551_365(w_551_365, w_174_048, w_204_674);
  nand2 I551_674(w_551_674, w_528_110, w_365_832);
  not1 I551_929(w_551_929, w_295_369);
  and2 I551_1193(w_551_1193, w_239_566, w_192_359);
  or2  I552_027(w_552_027, w_416_600, w_026_125);
  not1 I554_288(w_554_288, w_235_791);
  or2  I554_319(w_554_319, w_514_053, w_141_106);
  not1 I555_332(w_555_332, w_330_958);
  not1 I555_481(w_555_481, w_047_404);
  and2 I555_1052(w_555_1052, w_406_554, w_331_550);
  nand2 I555_1335(w_555_1335, w_354_460, w_387_720);
  and2 I555_1534(w_555_1534, w_250_222, w_306_1228);
  and2 I556_147(w_556_147, w_494_945, w_471_553);
  not1 I556_235(w_556_235, w_229_1253);
  not1 I556_258(w_556_258, w_180_352);
  and2 I556_272(w_556_272, w_375_1233, w_458_412);
  or2  I557_485(w_557_485, w_034_189, w_369_346);
  not1 I557_825(w_557_825, w_534_1231);
  nand2 I557_1075(w_557_1075, w_376_209, w_113_910);
  nand2 I559_669(w_559_669, w_337_369, w_154_181);
  and2 I559_922(w_559_922, w_011_172, w_280_389);
  nand2 I560_327(w_560_327, w_340_114, w_121_390);
  not1 I560_345(w_560_345, w_540_182);
  nand2 I560_1113(w_560_1113, w_474_412, w_089_578);
  nand2 I560_1382(w_560_1382, w_307_271, w_046_029);
  and2 I561_252(w_561_252, w_104_1263, w_410_008);
  nand2 I561_339(w_561_339, w_496_797, w_463_433);
  or2  I562_017(w_562_017, w_060_063, w_538_357);
  nand2 I563_139(w_563_139, w_473_1043, w_407_182);
  not1 I563_242(w_563_242, w_543_594);
  nand2 I563_721(w_563_721, w_040_407, w_204_064);
  nand2 I563_905(w_563_905, w_408_005, w_046_049);
  not1 I563_959(w_563_961, w_563_960);
  nand2 I563_960(w_563_962, w_563_961, w_014_646);
  or2  I563_961(w_563_963, w_435_916, w_563_962);
  and2 I563_962(w_563_960, w_130_508, w_563_963);
  nand2 I564_071(w_564_071, w_332_177, w_406_471);
  not1 I566_066(w_566_066, w_500_1299);
  nand2 I566_957(w_566_957, w_531_121, w_554_288);
  or2  I568_047(w_568_047, w_482_839, w_477_104);
  and2 I568_596(w_568_596, w_365_064, w_529_180);
  or2  I568_913(w_568_913, w_387_967, w_520_667);
  not1 I569_388(w_569_388, w_196_555);
  or2  I570_560(w_570_560, w_312_054, w_480_062);
  nand2 I570_1461(w_570_1461, w_103_232, w_179_361);
  nand2 I571_034(w_571_034, w_175_080, w_080_019);
  nand2 I571_1088(w_571_1088, w_431_1031, w_562_017);
  not1 I575_205(w_575_205, w_278_052);
  or2  I575_519(w_575_519, w_397_1463, w_202_662);
  nand2 I575_539(w_575_539, w_551_082, w_566_957);
  or2  I576_511(w_576_511, w_138_111, w_227_009);
  not1 I576_846(w_576_846, w_074_584);
  not1 I576_1032(w_576_1032, w_228_090);
  or2  I578_287(w_578_287, w_154_066, w_468_214);
  not1 I578_425(w_578_425, w_274_071);
  nand2 I578_634(w_578_634, w_235_669, w_514_1390);
  and2 I579_134(w_579_134, w_546_1098, w_306_1195);
  nand2 I579_721(w_579_721, w_459_383, w_434_633);
  nand2 I579_1003(w_579_1003, w_198_923, w_235_892);
  not1 I579_1598(w_579_1598, w_504_564);
  and2 I582_1282(w_582_1282, w_395_657, w_135_114);
  nand2 I582_1357(w_582_1357, w_135_387, w_388_936);
  nand2 I583_066(w_583_066, w_167_010, w_004_1532);
  or2  I583_224(w_583_224, w_088_1340, w_270_531);
  not1 I583_291(w_583_291, w_576_1032);
  nand2 I584_730(w_584_730, w_269_453, w_133_739);
  not1 I584_893(w_584_893, w_274_070);
  and2 I585_214(w_585_214, w_028_647, w_183_438);
  or2  I585_360(w_585_360, w_147_076, w_292_461);
  and2 I586_135(w_586_135, w_512_823, w_037_1389);
  not1 I586_969(w_586_969, w_035_194);
  nand2 I586_1406(w_586_1406, w_555_1052, w_374_798);
  and2 I587_856(w_587_856, w_252_617, w_489_036);
  or2  I587_869(w_587_869, w_522_090, w_503_694);
  nand2 I588_356(w_588_356, w_136_080, w_512_1078);
  nand2 I589_707(w_589_707, w_381_179, w_440_709);
  or2  I590_780(w_590_780, w_248_354, w_188_329);
  and2 I590_1014(w_590_1014, w_402_998, w_528_145);
  not1 I591_300(w_591_300, w_441_750);
  and2 I591_762(w_591_762, w_446_722, w_499_1419);
  nand2 I591_1100(w_591_1100, w_542_089, w_388_219);
  or2  I592_086(w_592_086, w_055_104, w_358_1178);
  not1 I592_142(w_592_142, w_487_790);
  and2 I592_687(w_592_687, w_555_332, w_307_274);
  nand2 I593_207(w_593_207, w_187_243, w_466_005);
  nand2 I595_157(w_595_157, w_011_845, w_551_674);
  and2 I595_178(w_595_178, w_498_402, w_175_084);
  nand2 I595_321(w_595_321, w_323_312, w_505_342);
  not1 I596_124(w_596_124, w_075_055);
  nand2 I596_343(w_596_343, w_176_1327, w_555_1534);
  not1 I597_068(w_597_068, w_337_027);
  and2 I597_813(w_597_813, w_510_051, w_347_053);
  or2  I598_265(w_598_265, w_162_093, w_372_215);
  or2  I599_010(w_599_010, w_462_134, w_318_336);
  not1 I599_034(w_599_034, w_433_070);
  and2 I599_056(w_599_056, w_171_037, w_515_456);
  or2  I600_523(w_600_523, w_174_581, w_066_753);
  or2  I600_663(w_600_663, w_115_129, w_497_364);
  or2  I601_015(w_601_015, w_030_706, w_244_796);
  or2  I601_063(w_601_063, w_260_029, w_187_081);
  and2 I601_438(w_601_438, w_255_132, w_583_291);
  or2  I601_471(w_601_471, w_353_240, w_575_539);
  or2  I602_517(w_602_517, w_080_034, w_598_265);
  nand2 I606_070(w_606_070, w_436_1601, w_038_200);
  nand2 I607_622(w_607_622, w_145_007, w_225_802);
  and2 I607_675(w_607_675, w_243_1362, w_244_892);
  nand2 I609_034(w_609_034, w_568_047, w_315_444);
  and2 I609_330(w_609_330, w_525_1141, w_027_093);
  not1 I610_888(w_610_890, w_610_889);
  not1 I610_889(w_610_891, w_610_890);
  not1 I610_890(w_610_892, w_610_891);
  not1 I610_891(w_610_893, w_610_892);
  nand2 I610_892(w_610_894, w_610_893, w_041_158);
  not1 I610_893(w_610_895, w_610_894);
  and2 I610_894(w_610_896, w_463_172, w_610_895);
  not1 I610_895(w_610_897, w_610_896);
  and2 I610_896(w_610_898, w_610_897, w_089_1226);
  or2  I610_897(w_610_899, w_396_560, w_610_898);
  and2 I610_898(w_610_889, w_610_899, w_160_041);
  or2  I611_122(w_611_122, w_422_306, w_050_393);
  or2  I611_200(w_611_200, w_200_197, w_216_467);
  nand2 I611_393(w_611_393, w_199_1644, w_343_016);
  nand2 I613_092(w_613_092, w_379_829, w_400_224);
  and2 I613_379(w_613_379, w_103_1200, w_324_008);
  nand2 I613_1491(w_613_1491, w_399_563, w_579_721);
  not1 I614_162(w_614_162, w_503_299);
  or2  I614_388(w_614_388, w_379_043, w_140_548);
  not1 I614_500(w_614_500, w_399_1417);
  not1 I615_216(w_615_216, w_556_272);
  or2  I616_164(w_616_164, w_266_543, w_273_595);
  or2  I616_1323(w_616_1323, w_257_360, w_138_142);
  and2 I617_575(w_617_575, w_084_091, w_343_227);
  nand2 I617_871(w_617_871, w_452_775, w_551_929);
  nand2 I618_405(w_618_405, w_151_1310, w_355_226);
  nand2 I619_033(w_619_033, w_327_516, w_302_402);
  and2 I619_080(w_619_080, w_132_039, w_113_390);
  not1 I620_074(w_620_074, w_107_468);
  or2  I620_379(w_620_379, w_321_097, w_376_513);
  nand2 I621_071(w_621_071, w_091_176, w_067_872);
  nand2 I621_268(w_621_268, w_390_195, w_509_322);
  nand2 I622_749(w_622_749, w_198_1377, w_163_041);
  not1 I623_435(w_623_435, w_253_005);
  nand2 I623_635(w_623_635, w_613_1491, w_023_1208);
  nand2 I624_1288(w_624_1288, w_185_1161, w_128_031);
  not1 I625_1222(w_625_1222, w_337_266);
  not1 I626_212(w_626_212, w_185_1466);
  not1 I626_1103(w_626_1103, w_127_516);
  nand2 I627_1504(w_627_1504, w_077_596, w_158_375);
  not1 I628_148(w_628_148, w_193_095);
  and2 I628_999(w_628_999, w_295_1365, w_112_350);
  or2  I628_1376(w_628_1376, w_190_479, w_287_022);
  not1 I629_028(w_629_028, w_144_271);
  nand2 I629_318(w_629_318, w_057_145, w_004_325);
  and2 I629_760(w_629_760, w_114_302, w_101_594);
  and2 I630_083(w_630_083, w_226_665, w_020_722);
  nand2 I630_312(w_630_312, w_308_256, w_497_391);
  and2 I631_069(w_631_069, w_091_132, w_561_252);
  nand2 I632_266(w_632_266, w_164_888, w_560_327);
  or2  I633_068(w_633_068, w_478_293, w_398_1205);
  or2  I633_696(w_633_696, w_151_694, w_430_088);
  nand2 I634_237(w_634_237, w_046_254, w_587_856);
  or2  I635_326(w_635_326, w_219_020, w_024_1561);
  not1 I635_649(w_635_649, w_194_853);
  nand2 I636_262(w_636_262, w_550_785, w_377_072);
  or2  I636_299(w_636_299, w_324_145, w_257_235);
  not1 I637_159(w_637_159, w_045_199);
  nand2 I637_508(w_637_508, w_579_1598, w_116_959);
  not1 I638_432(w_638_432, w_218_388);
  and2 I638_1113(w_638_1113, w_184_002, w_490_1421);
  and2 I638_1129(w_638_1129, w_443_718, w_246_168);
  not1 I639_313(w_639_313, w_617_871);
  nand2 I639_1097(w_639_1097, w_198_1352, w_014_001);
  nand2 I639_1572(w_639_1572, w_330_693, w_250_116);
  not1 I639_1573(w_639_1573, w_247_604);
  nand2 I640_066(w_640_066, w_620_379, w_427_021);
  not1 I640_496(w_640_496, w_461_310);
  or2  I640_710(w_640_710, w_117_532, w_251_282);
  nand2 I641_262(w_641_262, w_359_526, w_443_305);
  not1 I641_515(w_641_515, w_590_1014);
  nand2 I641_594(w_641_594, w_614_162, w_599_056);
  or2  I641_787(w_641_787, w_096_134, w_411_987);
  nand2 I642_231(w_642_231, w_095_387, w_347_1219);
  nand2 I642_268(w_642_268, w_512_679, w_141_076);
  nand2 I644_837(w_644_837, w_312_162, w_227_002);
  and2 I644_866(w_644_866, w_170_819, w_422_351);
  or2  I645_049(w_645_049, w_337_234, w_256_436);
  or2  I645_091(w_645_091, w_595_178, w_359_650);
  and2 I645_105(w_645_105, w_130_333, w_371_098);
  or2  I646_094(w_646_094, w_520_598, w_537_388);
  nand2 I647_214(w_647_214, w_262_131, w_548_509);
  and2 I647_288(w_647_288, w_284_140, w_629_760);
  nand2 I648_062(w_648_062, w_469_351, w_188_082);
  nand2 I648_1062(w_648_1062, w_201_117, w_584_893);
  not1 I649_568(w_649_568, w_338_1435);
  nand2 I650_134(w_650_134, w_564_071, w_248_059);
  not1 I650_173(w_650_173, w_382_185);
  and2 I651_012(w_651_012, w_134_893, w_479_1024);
  and2 I651_352(w_651_352, w_198_481, w_121_710);
  or2  I651_1455(w_651_1455, w_544_028, w_476_073);
  and2 I651_1483(w_651_1483, w_132_015, w_142_237);
  not1 I652_003(w_652_003, w_298_1289);
  not1 I652_032(w_652_032, w_167_006);
  nand2 I652_064(w_652_064, w_625_1222, w_122_175);
  not1 I654_208(w_654_208, w_251_010);
  not1 I655_134(w_655_134, w_329_460);
  or2  I655_1625(w_655_1625, w_046_120, w_274_039);
  or2  I657_1324(w_657_1324, w_379_194, w_082_265);
  nand2 I658_866(w_658_866, w_043_070, w_241_299);
  and2 I659_522(w_659_522, w_476_379, w_164_782);
  or2  I660_005(w_660_005, w_456_731, w_029_1057);
  or2  I660_064(w_660_064, w_033_1577, w_471_265);
  not1 I660_207(w_660_207, w_524_1505);
  and2 I660_223(w_660_223, w_043_016, w_177_1601);
  not1 I660_298(w_660_298, w_579_134);
  or2  I662_540(w_662_540, w_433_592, w_433_394);
  or2  I663_732(w_663_732, w_632_266, w_048_742);
  and2 I664_091(w_664_091, w_248_028, w_087_1104);
  and2 I665_324(w_665_324, w_463_044, w_265_699);
  nand2 I665_335(w_665_335, w_357_293, w_188_178);
  or2  I667_474(w_667_474, w_285_314, w_023_046);
  nand2 I668_104(w_668_104, w_519_189, w_563_139);
  not1 I668_967(w_668_967, w_453_196);
  and2 I669_042(w_669_042, w_289_1199, w_195_041);
  nand2 I669_044(w_669_044, w_402_569, w_513_1030);
  nand2 I669_079(w_669_079, w_611_393, w_387_317);
  not1 I669_136(w_669_138, w_669_137);
  nand2 I669_137(w_669_139, w_669_138, w_064_639);
  and2 I669_138(w_669_140, w_288_172, w_669_139);
  not1 I669_139(w_669_141, w_669_140);
  or2  I669_140(w_669_142, w_383_377, w_669_141);
  or2  I669_141(w_669_143, w_481_093, w_669_142);
  not1 I669_142(w_669_144, w_669_143);
  and2 I669_143(w_669_145, w_669_144, w_641_515);
  and2 I669_144(w_669_137, w_556_235, w_669_145);
  nand2 I670_119(w_670_119, w_536_150, w_071_130);
  nand2 I670_353(w_670_353, w_371_387, w_178_455);
  nand2 I670_636(w_670_636, w_478_815, w_070_369);
  and2 I671_330(w_671_330, w_283_1461, w_410_103);
  not1 I673_061(w_673_061, w_636_262);
  and2 I674_038(w_674_038, w_129_747, w_394_030);
  nand2 I674_041(w_674_041, w_242_064, w_601_063);
  nand2 I674_050(w_674_050, w_180_336, w_454_043);
  nand2 I675_004(w_675_004, w_456_769, w_588_356);
  or2  I675_012(w_675_012, w_549_352, w_557_485);
  nand2 I676_349(w_676_349, w_378_565, w_084_041);
  not1 I676_1465(w_676_1465, w_084_275);
  nand2 I677_132(w_677_132, w_135_385, w_537_615);
  or2  I678_238(w_678_238, w_133_411, w_417_017);
  nand2 I678_759(w_678_759, w_089_179, w_243_657);
  not1 I678_781(w_678_781, w_283_1219);
  and2 I679_272(w_679_272, w_614_500, w_316_101);
  nand2 I679_506(w_679_506, w_532_271, w_336_141);
  or2  I681_026(w_681_026, w_047_372, w_046_220);
  or2  I681_1392(w_681_1392, w_301_1280, w_646_094);
  or2  I682_001(w_682_001, w_018_100, w_179_351);
  and2 I682_042(w_682_042, w_418_673, w_448_252);
  nand2 I682_097(w_682_097, w_261_075, w_369_1193);
  and2 I682_148(w_682_148, w_645_049, w_396_254);
  nand2 I683_161(w_683_161, w_162_242, w_183_362);
  and2 I683_164(w_683_164, w_286_538, w_674_038);
  nand2 I683_238(w_683_238, w_667_474, w_078_109);
  not1 I685_1698(w_685_1698, w_403_223);
  nand2 I686_073(w_686_073, w_123_832, w_682_042);
  nand2 I686_417(w_686_417, w_575_519, w_478_1092);
  or2  I687_290(w_687_290, w_514_848, w_108_381);
  and2 I687_540(w_687_540, w_524_1502, w_100_900);
  nand2 I687_1614(w_687_1614, w_044_538, w_505_1503);
  and2 I688_909(w_688_909, w_323_403, w_181_095);
  and2 I690_753(w_690_753, w_515_679, w_106_854);
  and2 I691_286(w_691_286, w_601_438, w_638_1129);
  and2 I691_509(w_691_509, w_647_288, w_231_1104);
  nand2 I692_115(w_692_115, w_467_689, w_419_069);
  or2  I694_687(w_694_687, w_044_466, w_582_1357);
  or2  I694_874(w_694_874, w_488_641, w_021_272);
  nand2 I696_103(w_696_103, w_670_636, w_121_711);
  and2 I696_418(w_696_418, w_382_163, w_278_1207);
  nand2 I696_431(w_696_431, w_287_148, w_118_650);
  and2 I697_644(w_697_644, w_024_915, w_333_070);
  and2 I697_733(w_697_733, w_021_161, w_629_028);
  or2  I697_939(w_697_939, w_495_1084, w_110_862);
  nand2 I697_1369(w_697_1369, w_353_720, w_657_1324);
  not1 I698_1173(w_698_1173, w_163_290);
  or2  I699_079(w_699_079, w_642_268, w_256_060);
  and2 I700_106(w_700_106, w_358_692, w_317_1544);
  nand2 I700_818(w_700_818, w_650_134, w_293_441);
  not1 I701_276(w_701_276, w_362_481);
  nand2 I703_042(w_703_042, w_383_219, w_218_302);
  not1 I703_183(w_703_183, w_515_186);
  and2 I703_312(w_703_312, w_476_313, w_683_164);
  or2  I704_087(w_704_087, w_374_145, w_131_538);
  not1 I704_803(w_704_803, w_571_034);
  nand2 I704_1453(w_704_1453, w_401_517, w_173_762);
  and2 I705_087(w_705_087, w_538_864, w_474_300);
  not1 I706_587(w_706_587, w_499_1719);
  or2  I706_1392(w_706_1392, w_492_128, w_489_1344);
  not1 I707_418(w_707_418, w_568_913);
  and2 I708_131(w_708_131, w_629_318, w_531_628);
  nand2 I708_987(w_708_987, w_619_080, w_300_1448);
  or2  I708_1216(w_708_1216, w_049_132, w_401_063);
  nand2 I709_060(w_709_060, w_035_1425, w_445_301);
  and2 I711_891(w_711_891, w_084_271, w_091_132);
  or2  I712_441(w_712_441, w_310_223, w_476_191);
  and2 I712_442(w_712_442, w_475_095, w_183_1069);
  and2 I712_634(w_712_634, w_468_249, w_441_128);
  not1 I713_104(w_713_104, w_663_732);
  and2 I713_131(w_713_131, w_124_381, w_586_969);
  or2  I713_146(w_713_146, w_008_085, w_277_056);
  or2  I713_203(w_713_203, w_330_1024, w_002_575);
  and2 I714_604(w_714_604, w_678_238, w_252_349);
  and2 I715_306(w_715_306, w_361_238, w_083_004);
  or2  I715_605(w_715_605, w_236_391, w_149_076);
  and2 I715_843(w_715_843, w_664_091, w_195_311);
  not1 I716_110(w_716_110, w_691_286);
  not1 I716_135(w_716_135, w_170_1270);
  and2 I716_416(w_716_416, w_079_502, w_365_534);
  nand2 I716_418(w_716_418, w_534_1008, w_210_1199);
  nand2 I717_1135(w_717_1135, w_709_060, w_355_525);
  not1 I717_1608(w_717_1608, w_150_128);
  nand2 I719_461(w_719_461, w_675_012, w_162_795);
  nand2 I722_1277(w_722_1277, w_074_422, w_273_880);
  not1 I722_1323(w_722_1323, w_056_1172);
  and2 I722_1620(w_722_1622, w_611_122, w_722_1621);
  and2 I722_1621(w_722_1623, w_316_915, w_722_1622);
  or2  I722_1622(w_722_1624, w_184_004, w_722_1623);
  not1 I722_1623(w_722_1625, w_722_1624);
  nand2 I722_1624(w_722_1626, w_670_353, w_722_1625);
  nand2 I722_1625(w_722_1627, w_722_1626, w_298_828);
  or2  I722_1626(w_722_1628, w_722_1627, w_246_1608);
  or2  I722_1627(w_722_1621, w_320_484, w_722_1628);
  nand2 I723_166(w_723_166, w_478_367, w_506_135);
  and2 I724_167(w_724_167, w_430_014, w_660_207);
  and2 I724_444(w_724_444, w_193_173, w_584_730);
  nand2 I724_1149(w_724_1149, w_461_280, w_282_305);
  not1 I726_1725(w_726_1725, w_424_022);
  and2 I727_690(w_727_690, w_470_456, w_060_019);
  not1 I728_220(w_728_220, w_130_152);
  or2  I728_1474(w_728_1474, w_462_025, w_308_235);
  nand2 I729_404(w_729_404, w_246_112, w_534_014);
  not1 I730_029(w_730_029, w_001_1573);
  nand2 I730_695(w_730_695, w_546_258, w_215_1078);
  and2 I731_027(w_731_027, w_516_699, w_230_237);
  and2 I731_059(w_731_059, w_290_217, w_509_386);
  or2  I733_210(w_733_210, w_382_672, w_669_044);
  or2  I733_461(w_733_461, w_436_1391, w_560_1113);
  or2  I737_163(w_737_163, w_446_605, w_316_288);
  nand2 I739_100(w_739_100, w_232_385, w_641_594);
  nand2 I740_1463(w_740_1463, w_159_858, w_134_019);
  and2 I741_660(w_741_660, w_660_005, w_423_206);
  or2  I741_921(w_741_921, w_290_254, w_624_1288);
  or2  I742_065(w_742_065, w_357_401, w_416_1113);
  or2  I742_176(w_742_176, w_128_197, w_469_046);
  and2 I743_219(w_743_219, w_234_1075, w_246_986);
  not1 I744_084(w_744_084, w_609_330);
  and2 I744_349(w_744_349, w_289_1017, w_290_110);
  and2 I745_034(w_745_034, w_067_434, w_330_248);
  nand2 I745_1779(w_745_1779, w_347_1601, w_445_361);
  and2 I748_059(w_748_059, w_744_084, w_437_1574);
  and2 I748_137(w_748_137, w_052_037, w_279_205);
  not1 I748_352(w_748_352, w_344_141);
  nand2 I749_443(w_749_443, w_204_438, w_716_110);
  nand2 I749_660(w_749_660, w_704_1453, w_714_604);
  or2  I751_026(w_751_026, w_655_1625, w_694_874);
  not1 I752_789(w_752_789, w_368_1696);
  or2  I752_1842(w_752_1842, w_679_272, w_551_271);
  and2 I755_1157(w_755_1157, w_343_1177, w_297_041);
  or2  I756_029(w_756_029, w_642_231, w_652_064);
  or2  I756_402(w_756_402, w_075_109, w_284_987);
  not1 I758_301(w_758_301, w_430_130);
  nand2 I758_721(w_758_721, w_476_096, w_086_049);
  and2 I759_359(w_759_359, w_487_032, w_370_1007);
  not1 I761_029(w_761_029, w_051_121);
  not1 I761_408(w_761_408, w_717_1135);
  not1 I762_873(w_762_873, w_310_065);
  nand2 I762_973(w_762_973, w_216_306, w_047_465);
  nand2 I763_252(w_763_252, w_046_159, w_559_922);
  and2 I764_117(w_764_117, w_503_261, w_621_071);
  nand2 I766_241(w_766_241, w_507_110, w_585_214);
  or2  I768_099(w_768_099, w_283_034, w_751_026);
  or2  I768_1400(w_768_1400, w_182_243, w_046_133);
  or2  I768_1574(w_768_1574, w_190_1082, w_640_066);
  nand2 I769_202(w_769_204, w_170_903, w_769_203);
  or2  I769_203(w_769_205, w_259_392, w_769_204);
  or2  I769_204(w_769_206, w_769_205, w_583_066);
  or2  I769_205(w_769_207, w_769_206, w_596_343);
  and2 I769_206(w_769_208, w_769_207, w_004_279);
  and2 I769_207(w_769_209, w_560_345, w_769_208);
  nand2 I769_208(w_769_203, w_769_209, w_668_104);
  nand2 I770_377(w_770_377, w_659_522, w_059_228);
  nand2 I771_455(w_771_455, w_452_108, w_547_082);
  or2  I773_045(w_773_045, w_514_1099, w_247_877);
  and2 I773_106(w_773_106, w_160_212, w_496_959);
  not1 I773_158(w_773_158, w_143_328);
  or2  I774_273(w_774_273, w_756_402, w_083_007);
  not1 I774_275(w_774_275, w_285_507);
  or2  I774_358(w_774_358, w_242_001, w_188_553);
  or2  I774_402(w_774_402, w_284_1530, w_682_097);
  not1 I777_1423(w_777_1423, w_042_093);
  nand2 I778_157(w_778_157, w_544_081, w_429_200);
  not1 I779_268(w_779_268, w_205_933);
  not1 I779_1214(w_779_1214, w_157_020);
  or2  I781_001(w_781_001, w_112_987, w_582_1282);
  and2 I781_1578(w_781_1578, w_261_278, w_226_655);
  and2 I781_1927(w_781_1927, w_255_230, w_132_001);
  nand2 I782_660(w_782_660, w_502_289, w_504_314);
  and2 I782_860(w_782_860, w_549_284, w_175_090);
  or2  I783_1101(w_783_1101, w_090_145, w_523_688);
  nand2 I784_448(w_784_448, w_427_082, w_774_358);
  not1 I786_960(w_786_960, w_675_004);
  or2  I786_1041(w_786_1041, w_700_818, w_515_094);
  or2  I788_162(w_788_162, w_628_148, w_280_045);
  and2 I789_059(w_789_059, w_590_780, w_160_220);
  and2 I790_373(w_790_373, w_030_471, w_713_203);
  not1 I790_894(w_790_894, w_248_051);
  or2  I790_1308(w_790_1308, w_596_124, w_631_069);
  not1 I791_162(w_791_162, w_618_405);
  and2 I792_882(w_792_882, w_478_1191, w_095_059);
  or2  I793_071(w_793_071, w_093_034, w_184_010);
  or2  I793_376(w_793_376, w_637_159, w_264_425);
  not1 I794_021(w_794_021, w_079_005);
  or2  I794_319(w_794_319, w_471_359, w_011_587);
  nand2 I795_080(w_795_080, w_492_085, w_639_1097);
  not1 I796_506(w_796_506, w_589_707);
  not1 I796_1386(w_796_1386, w_507_047);
  or2  I796_1672(w_796_1672, w_392_1327, w_668_967);
  nand2 I797_000(w_797_000, w_313_033, w_128_091);
  not1 I797_284(w_797_284, w_483_094);
  nand2 I798_333(w_798_333, w_287_020, w_626_212);
  nand2 I798_611(w_798_611, w_060_074, w_729_404);
  nand2 I799_494(w_799_494, w_640_496, w_363_507);
  or2  I799_847(w_799_849, w_799_848, w_496_495);
  or2  I799_848(w_799_850, w_674_050, w_799_849);
  or2  I799_849(w_799_851, w_773_158, w_799_850);
  nand2 I799_850(w_799_852, w_799_851, w_271_175);
  not1 I799_851(w_799_853, w_799_852);
  nand2 I799_852(w_799_854, w_799_853, w_024_882);
  and2 I799_853(w_799_855, w_799_854, w_799_865);
  not1 I799_854(w_799_856, w_799_855);
  nand2 I799_855(w_799_848, w_651_012, w_799_856);
  or2  I799_856(w_799_861, w_799_860, w_409_773);
  or2  I799_857(w_799_862, w_799_861, w_292_804);
  not1 I799_858(w_799_863, w_799_862);
  not1 I799_859(w_799_860, w_799_855);
  and2 I799_860(w_799_865, w_478_1446, w_799_863);
  nand2 I800_598(w_800_598, w_408_015, w_082_179);
  and2 I803_018(w_803_018, w_459_833, w_551_365);
  or2  I803_122(w_803_122, w_544_040, w_137_007);
  or2  I803_464(w_803_464, w_692_115, w_708_987);
  or2  I805_553(w_805_553, w_321_092, w_149_489);
  or2  I807_312(w_807_312, w_548_923, w_102_797);
  or2  I807_337(w_807_337, w_792_882, w_502_250);
  nand2 I808_008(w_808_008, w_687_290, w_525_1399);
  or2  I808_810(w_808_810, w_793_071, w_557_825);
  nand2 I808_986(w_808_986, w_325_1534, w_429_1594);
  and2 I809_122(w_809_122, w_313_025, w_210_412);
  nand2 I809_1170(w_809_1170, w_396_282, w_109_077);
  not1 I810_657(w_810_657, w_469_529);
  nand2 I810_754(w_810_754, w_730_029, w_727_690);
  and2 I810_824(w_810_824, w_479_1741, w_084_474);
  nand2 I811_1068(w_811_1068, w_092_426, w_098_494);
  nand2 I811_1380(w_811_1380, w_733_461, w_315_232);
  or2  I811_1552(w_811_1552, w_138_031, w_633_696);
  nand2 I811_1655(w_811_1657, w_811_1656, w_800_598);
  nand2 I811_1656(w_811_1658, w_811_1657, w_353_181);
  and2 I811_1657(w_811_1656, w_811_1670, w_811_1658);
  not1 I811_1658(w_811_1663, w_811_1662);
  and2 I811_1659(w_811_1664, w_811_1663, w_674_041);
  not1 I811_1660(w_811_1665, w_811_1664);
  or2  I811_1661(w_811_1666, w_232_480, w_811_1665);
  not1 I811_1662(w_811_1667, w_811_1666);
  not1 I811_1663(w_811_1668, w_811_1667);
  not1 I811_1664(w_811_1662, w_811_1656);
  and2 I811_1665(w_811_1670, w_194_797, w_811_1668);
  not1 I813_1102(w_813_1102, w_442_759);
  or2  I814_632(w_814_632, w_046_012, w_600_663);
  and2 I815_878(w_815_878, w_141_720, w_499_181);
  or2  I817_481(w_817_481, w_427_172, w_146_071);
  and2 I817_484(w_817_484, w_073_031, w_768_1400);
  or2  I818_030(w_818_030, w_698_1173, w_368_986);
  and2 I818_157(w_818_157, w_509_148, w_814_632);
  and2 I819_177(w_819_177, w_231_1772, w_274_054);
  nand2 I819_178(w_819_178, w_636_299, w_613_379);
  not1 I819_190(w_819_190, w_488_278);
  nand2 I820_230(w_820_230, w_368_1526, w_811_1068);
  and2 I820_664(w_820_664, w_711_891, w_181_306);
  nand2 I821_012(w_821_012, w_808_008, w_724_444);
  or2  I825_278(w_825_278, w_509_110, w_583_224);
  nand2 I826_369(w_826_369, w_237_638, w_277_085);
  or2  I826_436(w_826_438, w_826_437, w_105_1459);
  or2  I826_437(w_826_439, w_826_438, w_161_455);
  and2 I826_438(w_826_440, w_826_439, w_826_452);
  nand2 I826_439(w_826_437, w_826_440, w_796_506);
  and2 I826_440(w_826_445, w_826_444, w_181_1114);
  or2  I826_441(w_826_446, w_826_445, w_016_013);
  nand2 I826_442(w_826_447, w_501_352, w_826_446);
  nand2 I826_443(w_826_448, w_826_447, w_807_337);
  and2 I826_444(w_826_449, w_826_448, w_277_292);
  and2 I826_445(w_826_450, w_826_449, w_059_023);
  not1 I826_446(w_826_444, w_826_440);
  and2 I826_447(w_826_452, w_506_138, w_826_450);
  nand2 I827_021(w_827_021, w_001_1685, w_239_601);
  or2  I827_820(w_827_820, w_791_162, w_645_105);
  or2  I828_066(w_828_066, w_578_287, w_278_414);
  or2  I828_715(w_828_715, w_299_691, w_433_560);
  and2 I829_391(w_829_391, w_686_417, w_748_137);
  or2  I830_022(w_830_022, w_749_443, w_440_814);
  or2  I831_1052(w_831_1052, w_818_030, w_135_346);
  not1 I832_266(w_832_266, w_576_846);
  and2 I833_562(w_833_562, w_388_751, w_648_1062);
  nand2 I834_1377(w_834_1377, w_180_239, w_361_317);
  nand2 I835_622(w_835_622, w_697_1369, w_476_389);
  nand2 I836_246(w_836_246, w_669_042, w_283_1149);
  nand2 I838_1026(w_838_1026, w_070_212, w_461_696);
  or2  I841_642(w_841_642, w_360_542, w_258_378);
  or2  I841_1177(w_841_1177, w_827_021, w_818_157);
  or2  I841_1412(w_841_1412, w_090_606, w_421_311);
  or2  I841_1480(w_841_1480, w_493_441, w_192_382);
  not1 I842_151(w_842_151, w_743_219);
  not1 I843_173(w_843_173, w_036_875);
  nand2 I843_278(w_843_278, w_655_134, w_703_312);
  nand2 I844_323(w_844_323, w_820_230, w_808_810);
  and2 I845_041(w_845_041, w_323_461, w_548_356);
  nand2 I847_251(w_847_251, w_510_261, w_682_001);
  nand2 I847_421(w_847_421, w_617_575, w_006_157);
  and2 I848_264(w_848_264, w_554_319, w_055_473);
  not1 I848_349(w_848_349, w_344_139);
  nand2 I848_565(w_848_565, w_679_506, w_358_1499);
  and2 I848_723(w_848_723, w_069_1776, w_156_041);
  nand2 I849_242(w_849_242, w_203_384, w_623_635);
  and2 I850_1264(w_850_1264, w_540_326, w_198_1667);
  not1 I851_1287(w_851_1289, w_851_1288);
  and2 I851_1288(w_851_1290, w_851_1289, w_169_068);
  and2 I851_1289(w_851_1291, w_239_367, w_851_1290);
  nand2 I851_1290(w_851_1292, w_851_1291, w_019_438);
  not1 I851_1291(w_851_1293, w_851_1292);
  nand2 I851_1292(w_851_1294, w_851_1293, w_040_590);
  not1 I851_1293(w_851_1295, w_851_1294);
  not1 I851_1294(w_851_1296, w_851_1295);
  and2 I851_1295(w_851_1297, w_851_1296, w_755_1157);
  or2  I851_1296(w_851_1288, w_851_1297, w_778_157);
  or2  I852_269(w_852_269, w_487_1147, w_114_116);
  not1 I855_166(w_855_166, w_566_066);
  not1 I855_946(w_855_946, w_214_754);
  and2 I856_1410(w_856_1410, w_312_133, w_276_145);
  and2 I858_124(w_858_124, w_611_200, w_045_255);
  and2 I858_381(w_858_381, w_826_369, w_556_258);
  or2  I860_017(w_860_017, w_628_1376, w_304_1341);
  and2 I860_405(w_860_405, w_084_233, w_041_278);
  or2  I860_903(w_860_903, w_571_1088, w_756_029);
  nand2 I860_1045(w_860_1045, w_439_508, w_328_005);
  and2 I862_052(w_862_052, w_111_343, w_286_530);
  nand2 I863_096(w_863_096, w_670_119, w_848_565);
  and2 I863_292(w_863_292, w_328_005, w_317_649);
  nand2 I863_388(w_863_390, w_520_1416, w_863_389);
  or2  I863_389(w_863_391, w_121_114, w_863_390);
  not1 I863_390(w_863_392, w_863_391);
  and2 I863_391(w_863_393, w_185_333, w_863_392);
  or2  I863_392(w_863_394, w_563_721, w_863_393);
  or2  I863_393(w_863_389, w_863_411, w_863_394);
  not1 I863_394(w_863_399, w_863_398);
  or2  I863_395(w_863_400, w_863_399, w_547_437);
  not1 I863_396(w_863_401, w_863_400);
  and2 I863_397(w_863_402, w_863_401, w_224_413);
  nand2 I863_398(w_863_403, w_863_402, w_697_733);
  nand2 I863_399(w_863_404, w_863_403, w_484_362);
  not1 I863_400(w_863_405, w_863_404);
  or2  I863_401(w_863_406, w_863_405, w_290_399);
  not1 I863_402(w_863_407, w_863_406);
  and2 I863_403(w_863_408, w_212_332, w_863_407);
  not1 I863_404(w_863_409, w_863_408);
  not1 I863_405(w_863_398, w_863_389);
  and2 I863_406(w_863_411, w_432_171, w_863_409);
  not1 I864_076(w_864_076, w_064_1438);
  or2  I865_178(w_865_178, w_833_562, w_121_517);
  or2  I866_722(w_866_722, w_848_349, w_863_096);
  or2  I866_1044(w_866_1044, w_135_258, w_362_483);
  or2  I868_223(w_868_223, w_027_198, w_404_266);
  or2  I871_000(w_871_000, w_374_1192, w_525_175);
  or2  I874_219(w_874_219, w_302_195, w_081_377);
  or2  I876_063(w_876_063, w_708_1216, w_496_1215);
  and2 I876_1135(w_876_1135, w_295_422, w_706_587);
  nand2 I877_566(w_877_566, w_774_402, w_166_597);
  nand2 I877_632(w_877_632, w_701_276, w_786_960);
  and2 I880_1190(w_880_1190, w_448_423, w_794_319);
  not1 I882_384(w_882_384, w_346_528);
  not1 I882_737(w_882_737, w_586_135);
  or2  I885_1687(w_885_1687, w_774_275, w_607_675);
  and2 I886_088(w_886_088, w_551_1193, w_599_034);
  not1 I888_1871(w_888_1871, w_524_121);
  nand2 I889_030(w_889_030, w_377_193, w_409_138);
  not1 I889_097(w_889_097, w_389_1637);
  not1 I890_411(w_890_411, w_219_172);
  or2  I890_822(w_890_822, w_283_1410, w_392_480);
  and2 I892_214(w_892_214, w_681_1392, w_216_540);
  not1 I893_056(w_893_056, w_175_091);
  not1 I894_393(w_894_393, w_326_383);
  and2 I894_585(w_894_587, w_894_586, w_570_1461);
  and2 I894_586(w_894_588, w_489_1324, w_894_587);
  and2 I894_587(w_894_589, w_116_454, w_894_588);
  or2  I894_588(w_894_590, w_164_146, w_894_589);
  nand2 I894_589(w_894_591, w_894_590, w_083_015);
  and2 I894_590(w_894_586, w_894_591, w_894_607);
  not1 I894_591(w_894_596, w_894_595);
  not1 I894_592(w_894_597, w_894_596);
  and2 I894_593(w_894_598, w_894_597, w_525_366);
  and2 I894_594(w_894_599, w_894_598, w_178_586);
  nand2 I894_595(w_894_600, w_252_382, w_894_599);
  not1 I894_596(w_894_601, w_894_600);
  or2  I894_597(w_894_602, w_894_601, w_451_632);
  nand2 I894_598(w_894_603, w_144_763, w_894_602);
  nand2 I894_599(w_894_604, w_762_973, w_894_603);
  or2  I894_600(w_894_605, w_894_604, w_789_059);
  not1 I894_601(w_894_595, w_894_586);
  and2 I894_602(w_894_607, w_479_643, w_894_605);
  nand2 I895_037(w_895_037, w_373_471, w_813_1102);
  and2 I897_1328(w_897_1330, w_211_212, w_897_1329);
  and2 I897_1329(w_897_1331, w_897_1330, w_093_070);
  or2  I897_1330(w_897_1332, w_897_1331, w_354_1250);
  not1 I897_1331(w_897_1333, w_897_1332);
  nand2 I897_1332(w_897_1334, w_897_1333, w_650_173);
  nand2 I897_1333(w_897_1335, w_214_230, w_897_1334);
  and2 I897_1334(w_897_1336, w_184_002, w_897_1335);
  and2 I897_1335(w_897_1337, w_897_1336, w_087_1494);
  or2  I897_1336(w_897_1338, w_249_423, w_897_1337);
  and2 I897_1337(w_897_1329, w_897_1338, w_163_147);
  nand2 I901_088(w_901_088, w_509_068, w_616_164);
  nand2 I901_574(w_901_574, w_162_130, w_607_622);
  and2 I901_607(w_901_607, w_035_1112, w_315_556);
  nand2 I902_415(w_902_415, w_424_025, w_868_223);
  nand2 I903_455(w_903_455, w_681_026, w_724_1149);
  not1 I905_262(w_905_262, w_623_435);
  nand2 I907_426(w_907_426, w_669_079, w_847_421);
  and2 I908_1300(w_908_1300, w_198_1676, w_431_239);
  nand2 I910_116(w_910_116, w_803_122, w_328_013);
  nand2 I911_069(w_911_069, w_124_466, w_134_414);
  and2 I912_120(w_912_120, w_421_143, w_615_216);
  nand2 I912_152(w_912_152, w_696_418, w_733_210);
  or2  I912_239(w_912_239, w_288_321, w_660_298);
  and2 I912_1012(w_912_1012, w_770_377, w_803_464);
  nand2 I915_132(w_915_132, w_025_1134, w_819_178);
  nand2 I915_948(w_915_948, w_540_341, w_200_317);
  and2 I916_191(w_916_191, w_235_106, w_708_131);
  and2 I916_732(w_916_732, w_424_021, w_793_376);
  nand2 I919_1870(w_919_1872, w_919_1871, w_406_870);
  or2  I919_1871(w_919_1873, w_919_1872, w_431_218);
  and2 I919_1872(w_919_1874, w_919_1873, w_478_665);
  and2 I919_1873(w_919_1875, w_919_1874, w_601_015);
  nand2 I919_1874(w_919_1876, w_412_028, w_919_1875);
  nand2 I919_1875(w_919_1877, w_919_1876, w_597_813);
  and2 I919_1876(w_919_1878, w_110_981, w_919_1877);
  not1 I919_1877(w_919_1871, w_919_1878);
  nand2 I921_020(w_921_020, w_712_441, w_217_197);
  nand2 I922_1398(w_922_1398, w_592_086, w_843_278);
  nand2 I922_1533(w_922_1533, w_049_962, w_098_276);
  nand2 I924_311(w_924_311, w_651_1455, w_715_306);
  or2  I925_563(w_925_563, w_059_572, w_449_347);
  nand2 I925_784(w_925_784, w_270_271, w_266_478);
  and2 I928_200(w_928_200, w_116_395, w_848_723);
  and2 I932_294(w_932_294, w_467_390, w_196_432);
  or2  I932_853(w_932_853, w_654_208, w_744_349);
  and2 I936_1058(w_936_1058, w_730_695, w_912_239);
  and2 I937_329(w_937_329, w_141_720, w_014_437);
  not1 I939_556(w_939_556, w_328_006);
  nand2 I940_013(w_940_013, w_635_649, w_758_721);
  and2 I940_080(w_940_080, w_013_132, w_035_1619);
  not1 I940_140(w_940_140, w_557_1075);
  not1 I941_1117(w_941_1119, w_941_1118);
  not1 I941_1118(w_941_1120, w_941_1119);
  and2 I941_1119(w_941_1118, w_838_1026, w_941_1120);
  not1 I942_113(w_942_113, w_168_399);
  not1 I949_751(w_949_751, w_786_1041);
  and2 I951_471(w_951_471, w_155_1257, w_758_301);
  or2  I952_247(w_952_247, w_433_631, w_901_088);
  and2 I957_171(w_957_171, w_442_118, w_088_1214);
  or2  I962_105(w_962_105, w_741_660, w_085_146);
  not1 I963_263(w_963_263, w_267_476);
  and2 I966_336(w_966_336, w_821_012, w_348_167);
  nand2 I966_460(w_966_462, w_966_461, w_966_480);
  nand2 I966_461(w_966_463, w_830_022, w_966_462);
  or2  I966_462(w_966_464, w_487_1069, w_966_463);
  nand2 I966_463(w_966_465, w_966_464, w_267_432);
  and2 I966_464(w_966_466, w_966_465, w_876_063);
  and2 I966_465(w_966_461, w_032_140, w_966_466);
  or2  I966_466(w_966_471, w_966_470, w_047_545);
  and2 I966_467(w_966_472, w_690_753, w_966_471);
  nand2 I966_468(w_966_473, w_966_472, w_259_070);
  or2  I966_469(w_966_474, w_966_473, w_510_180);
  and2 I966_470(w_966_475, w_966_474, w_016_028);
  and2 I966_471(w_966_476, w_966_475, w_512_268);
  or2  I966_472(w_966_477, w_966_476, w_481_1485);
  or2  I966_473(w_966_478, w_213_512, w_966_477);
  not1 I966_474(w_966_470, w_966_462);
  and2 I966_475(w_966_480, w_752_1842, w_966_478);
  not1 I968_263(w_968_263, w_699_079);
  not1 I968_742(w_968_742, w_871_000);
  nand2 I969_298(w_969_298, w_545_1157, w_763_252);
  not1 I975_392(w_975_392, w_046_276);
  and2 I975_669(w_975_669, w_200_137, w_439_531);
  or2  I975_1237(w_975_1237, w_406_964, w_456_283);
  or2  I976_215(w_976_215, w_858_381, w_299_100);
  not1 I976_286(w_976_288, w_976_287);
  and2 I976_287(w_976_289, w_341_249, w_976_288);
  or2  I976_288(w_976_290, w_976_289, w_164_498);
  and2 I976_289(w_976_291, w_137_112, w_976_290);
  nand2 I976_290(w_976_292, w_976_291, w_834_1377);
  or2  I976_291(w_976_293, w_299_113, w_976_292);
  or2  I976_292(w_976_294, w_599_010, w_976_293);
  nand2 I976_293(w_976_295, w_976_303, w_976_294);
  and2 I976_294(w_976_287, w_427_055, w_976_295);
  or2  I976_295(w_976_300, w_271_056, w_976_299);
  nand2 I976_296(w_976_301, w_976_300, w_660_223);
  not1 I976_297(w_976_299, w_976_295);
  and2 I976_298(w_976_303, w_660_064, w_976_301);
  not1 I978_267(w_978_267, w_302_122);
  and2 I979_555(w_979_555, w_299_740, w_255_136);
  not1 I979_812(w_979_812, w_415_207);
  nand2 I980_107(w_980_107, w_281_975, w_639_313);
  nand2 I981_087(w_981_087, w_894_393, w_586_1406);
  or2  I987_771(w_987_771, w_414_110, w_364_185);
  and2 I988_096(w_988_096, w_575_205, w_463_473);
  and2 I991_026(w_991_026, w_922_1398, w_052_173);
  not1 I996_217(w_996_217, w_795_080);
  or2  I996_1459(w_996_1461, w_996_1460, w_797_284);
  or2  I996_1460(w_996_1462, w_996_1461, w_356_068);
  not1 I996_1461(w_996_1463, w_996_1462);
  not1 I996_1462(w_996_1464, w_996_1463);
  or2  I996_1463(w_996_1465, w_996_1482, w_996_1464);
  not1 I996_1464(w_996_1466, w_996_1465);
  or2  I996_1465(w_996_1467, w_252_658, w_996_1466);
  or2  I996_1466(w_996_1460, w_696_431, w_996_1467);
  nand2 I996_1467(w_996_1472, w_373_465, w_996_1471);
  not1 I996_1468(w_996_1473, w_996_1472);
  or2  I996_1469(w_996_1474, w_996_1473, w_691_509);
  not1 I996_1470(w_996_1475, w_996_1474);
  nand2 I996_1471(w_996_1476, w_817_481, w_996_1475);
  not1 I996_1472(w_996_1477, w_996_1476);
  and2 I996_1473(w_996_1478, w_996_1477, w_797_000);
  not1 I996_1474(w_996_1479, w_996_1478);
  or2  I996_1475(w_996_1480, w_996_1479, w_311_453);
  not1 I996_1476(w_996_1471, w_996_1465);
  and2 I996_1477(w_996_1482, w_741_921, w_996_1480);
  and2 I999_921(w_999_921, w_020_858, w_052_1907);
  not1 I1002_108(w_1002_108, w_841_1177);
  not1 I1002_191(w_1002_191, w_742_176);
  not1 I1004_487(w_1004_487, w_019_428);
  not1 I1005_1726(w_1005_1726, w_391_048);
  nand2 I1006_1160(w_1006_1160, w_167_054, w_200_386);
  not1 I1010_649(w_1010_649, w_688_909);
  not1 I1011_314(w_1011_314, w_841_1412);
  and2 I1012_147(w_1012_147, w_902_415, w_483_425);
  nand2 I1012_353(w_1012_353, w_848_264, w_293_535);
  and2 I1013_326(w_1013_326, w_142_340, w_912_1012);
  not1 I1017_151(w_1017_151, w_460_906);
  and2 I1017_222(w_1017_222, w_446_536, w_705_087);
  or2  I1018_190(w_1018_190, w_256_421, w_401_383);
  not1 I1018_418(w_1018_418, w_097_473);
  or2  I1018_633(w_1018_633, w_541_073, w_210_1039);
  or2  I1019_850(w_1019_850, w_517_039, w_477_098);
  nand2 I1025_1532(w_1025_1532, w_639_1572, w_492_086);
  and2 I1030_528(w_1030_528, w_015_188, w_424_016);
  and2 I1033_020(w_1033_020, w_232_153, w_999_921);
  nand2 I1034_506(w_1034_506, w_860_405, w_115_434);
  not1 I1035_002(w_1035_002, w_764_117);
  or2  I1035_074(w_1035_074, w_895_037, w_460_1204);
  not1 I1036_151(w_1036_151, w_815_878);
  or2  I1036_805(w_1036_805, w_294_499, w_309_001);
  not1 I1038_1382(w_1038_1382, w_497_331);
  not1 I1041_374(w_1041_374, w_803_018);
  not1 I1044_059(w_1044_059, w_728_220);
  nand2 I1045_096(w_1045_096, w_996_217, w_362_212);
  or2  I1047_1404(w_1047_1404, w_719_461, w_228_032);
  and2 I1049_021(w_1049_021, w_1002_191, w_351_028);
  not1 I1050_082(w_1050_082, w_703_183);
  not1 I1053_806(w_1053_806, w_740_1463);
  or2  I1055_134(w_1055_134, w_506_472, w_292_892);
  nand2 I1055_452(w_1055_454, w_1055_453, w_728_1474);
  and2 I1055_453(w_1055_455, w_1055_454, w_556_147);
  not1 I1055_454(w_1055_456, w_1055_455);
  or2  I1055_455(w_1055_457, w_1055_456, w_788_162);
  not1 I1055_456(w_1055_458, w_1055_457);
  or2  I1055_457(w_1055_459, w_936_1058, w_1055_458);
  not1 I1055_458(w_1055_460, w_1055_459);
  and2 I1055_459(w_1055_461, w_135_221, w_1055_460);
  or2  I1055_460(w_1055_462, w_289_281, w_1055_461);
  and2 I1055_461(w_1055_463, w_088_1150, w_1055_462);
  or2  I1055_462(w_1055_464, w_628_999, w_1055_463);
  and2 I1055_463(w_1055_453, w_1055_464, w_940_080);
  and2 I1056_111(w_1056_111, w_888_1871, w_126_220);
  and2 I1057_865(w_1057_865, w_724_167, w_639_1573);
  nand2 I1060_189(w_1060_189, w_880_1190, w_112_770);
  nand2 I1064_040(w_1064_040, w_345_1056, w_652_032);
  not1 I1065_185(w_1065_185, w_024_1579);
  and2 I1065_229(w_1065_229, w_713_131, w_361_090);
  and2 I1065_406(w_1065_406, w_175_066, w_270_079);
  nand2 I1066_974(w_1066_974, w_782_660, w_665_324);
  and2 I1069_285(w_1069_285, w_395_966, w_652_003);
  and2 I1069_553(w_1069_553, w_179_1221, w_828_066);
  not1 I1069_579(w_1069_579, w_407_014);
  not1 I1072_321(w_1072_321, w_1036_151);
  not1 I1075_1903(w_1075_1905, w_1075_1904);
  not1 I1075_1904(w_1075_1906, w_1075_1905);
  and2 I1075_1905(w_1075_1907, w_781_1927, w_1075_1906);
  nand2 I1075_1906(w_1075_1908, w_357_083, w_1075_1907);
  and2 I1075_1907(w_1075_1909, w_1075_1908, w_087_1603);
  nand2 I1075_1908(w_1075_1910, w_1075_1924, w_1075_1909);
  not1 I1075_1909(w_1075_1911, w_1075_1910);
  and2 I1075_1910(w_1075_1904, w_1075_1911, w_697_644);
  and2 I1075_1911(w_1075_1916, w_925_563, w_1075_1915);
  and2 I1075_1912(w_1075_1917, w_1075_1916, w_809_1170);
  nand2 I1075_1913(w_1075_1918, w_1041_374, w_1075_1917);
  or2  I1075_1914(w_1075_1919, w_671_330, w_1075_1918);
  and2 I1075_1915(w_1075_1920, w_1075_1919, w_827_820);
  not1 I1075_1916(w_1075_1921, w_1075_1920);
  nand2 I1075_1917(w_1075_1922, w_570_560, w_1075_1921);
  not1 I1075_1918(w_1075_1915, w_1075_1910);
  and2 I1075_1919(w_1075_1924, w_597_068, w_1075_1922);
  nand2 I1076_206(w_1076_206, w_538_713, w_032_244);
  not1 I1078_045(w_1078_045, w_247_1659);
  and2 I1078_080(w_1078_082, w_1078_081, w_845_041);
  or2  I1078_081(w_1078_083, w_1018_190, w_1078_082);
  nand2 I1078_082(w_1078_084, w_549_164, w_1078_083);
  not1 I1078_083(w_1078_085, w_1078_084);
  not1 I1078_084(w_1078_086, w_1078_085);
  or2  I1078_085(w_1078_087, w_1078_086, w_026_1287);
  not1 I1078_086(w_1078_088, w_1078_087);
  or2  I1078_087(w_1078_089, w_1078_088, w_1069_579);
  or2  I1078_088(w_1078_090, w_1078_089, w_638_1113);
  and2 I1078_089(w_1078_091, w_1078_090, w_498_636);
  and2 I1078_090(w_1078_092, w_1078_091, w_1017_151);
  not1 I1078_091(w_1078_081, w_1078_092);
  nand2 I1080_723(w_1080_723, w_102_462, w_336_1049);
  or2  I1083_094(w_1083_094, w_418_1325, w_047_194);
  and2 I1087_369(w_1087_369, w_863_292, w_649_568);
  or2  I1088_775(w_1088_775, w_630_312, w_874_219);
  nand2 I1088_842(w_1088_842, w_078_053, w_048_312);
  not1 I1092_449(w_1092_449, w_430_067);
  not1 I1093_019(w_1093_019, w_979_812);
  not1 I1093_049(w_1093_049, w_1092_449);
  not1 I1095_044(w_1095_044, w_139_516);
  not1 I1097_525(w_1097_525, w_493_225);
  or2  I1097_1090(w_1097_1090, w_1083_094, w_901_574);
  not1 I1099_048(w_1099_048, w_097_119);
  and2 I1104_019(w_1104_019, w_685_1698, w_156_193);
  and2 I1108_010(w_1108_010, w_299_1020, w_1099_048);
  nand2 I1109_060(w_1109_060, w_969_298, w_779_268);
  or2  I1111_1175(w_1111_1175, w_707_418, w_055_422);
  nand2 I1112_1168(w_1112_1168, w_235_947, w_731_027);
  and2 I1112_1747(w_1112_1749, w_1087_369, w_1112_1748);
  not1 I1112_1748(w_1112_1750, w_1112_1749);
  not1 I1112_1749(w_1112_1751, w_1112_1750);
  and2 I1112_1750(w_1112_1752, w_057_632, w_1112_1751);
  not1 I1112_1751(w_1112_1753, w_1112_1752);
  nand2 I1112_1752(w_1112_1754, w_1112_1753, w_499_436);
  nand2 I1112_1753(w_1112_1755, w_1055_134, w_1112_1754);
  or2  I1112_1754(w_1112_1756, w_1112_1755, w_276_134);
  and2 I1112_1755(w_1112_1748, w_1112_1756, w_591_1100);
  and2 I1114_194(w_1114_194, w_443_369, w_291_793);
  or2  I1117_515(w_1117_515, w_1044_059, w_641_787);
  nand2 I1118_533(w_1118_533, w_021_074, w_563_242);
  or2  I1118_1454(w_1118_1456, w_560_1382, w_1118_1455);
  or2  I1118_1455(w_1118_1457, w_1118_1456, w_420_1439);
  and2 I1118_1456(w_1118_1458, w_794_021, w_1118_1457);
  not1 I1118_1457(w_1118_1459, w_1118_1458);
  nand2 I1118_1458(w_1118_1460, w_1118_1459, w_811_1380);
  nand2 I1118_1459(w_1118_1461, w_135_304, w_1118_1460);
  or2  I1118_1460(w_1118_1462, w_1118_1461, w_510_260);
  not1 I1118_1461(w_1118_1463, w_1118_1462);
  not1 I1118_1462(w_1118_1464, w_1118_1463);
  or2  I1118_1463(w_1118_1455, w_1118_1464, w_916_191);
  or2  I1124_1428(w_1124_1428, w_326_363, w_745_1779);
  or2  I1126_121(w_1126_121, w_592_687, w_850_1264);
  or2  I1128_466(w_1128_466, w_427_169, w_446_247);
  and2 I1131_656(w_1131_656, w_005_910, w_561_339);
  and2 I1131_664(w_1131_664, w_882_737, w_1124_1428);
  and2 I1132_1116(w_1132_1118, w_1132_1117, w_259_272);
  not1 I1132_1117(w_1132_1119, w_1132_1118);
  and2 I1132_1118(w_1132_1120, w_1132_1119, w_287_271);
  or2  I1132_1119(w_1132_1121, w_796_1386, w_1132_1120);
  not1 I1132_1120(w_1132_1122, w_1132_1121);
  and2 I1132_1121(w_1132_1123, w_416_364, w_1132_1122);
  nand2 I1132_1122(w_1132_1117, w_745_034, w_1132_1123);
  and2 I1133_1692(w_1133_1692, w_483_314, w_396_001);
  or2  I1134_1163(w_1134_1163, w_366_011, w_716_418);
  or2  I1137_216(w_1137_216, w_647_214, w_336_1116);
  and2 I1139_1355(w_1139_1355, w_104_776, w_042_141);
  or2  I1142_154(w_1142_154, w_043_041, w_268_357);
  not1 I1148_133(w_1148_133, w_1128_466);
  and2 I1157_360(w_1157_360, w_444_113, w_171_1112);
  and2 I1158_191(w_1158_191, w_715_605, w_1065_406);
  not1 I1161_784(w_1161_784, w_321_082);
  not1 I1162_232(w_1162_232, w_495_1004);
  not1 I1165_045(w_1165_045, w_064_749);
  not1 I1166_032(w_1166_032, w_252_005);
  or2  I1168_039(w_1168_039, w_067_225, w_045_213);
  not1 I1169_327(w_1169_327, w_592_142);
  or2  I1173_1388(w_1173_1388, w_678_759, w_774_273);
  and2 I1176_1250(w_1176_1252, w_290_007, w_1176_1251);
  nand2 I1176_1251(w_1176_1253, w_1176_1252, w_217_203);
  nand2 I1176_1252(w_1176_1254, w_1176_1253, w_798_333);
  nand2 I1176_1253(w_1176_1255, w_293_1017, w_1176_1254);
  nand2 I1176_1254(w_1176_1256, w_189_024, w_1176_1255);
  or2  I1176_1255(w_1176_1257, w_1176_1256, w_276_134);
  not1 I1176_1256(w_1176_1258, w_1176_1257);
  nand2 I1176_1257(w_1176_1259, w_860_903, w_1176_1258);
  nand2 I1176_1258(w_1176_1260, w_1176_1259, w_218_637);
  or2  I1176_1259(w_1176_1261, w_513_409, w_1176_1260);
  and2 I1176_1260(w_1176_1262, w_843_173, w_1176_1261);
  nand2 I1176_1261(w_1176_1251, w_1176_1262, w_1093_019);
  nand2 I1178_104(w_1178_104, w_825_278, w_777_1423);
  and2 I1181_634(w_1181_634, w_122_002, w_373_1800);
  nand2 I1181_769(w_1181_769, w_876_1135, w_1080_723);
  not1 I1183_177(w_1183_177, w_645_091);
  and2 I1190_258(w_1190_258, w_712_442, w_696_103);
  nand2 I1192_779(w_1192_779, w_915_132, w_1060_189);
  nand2 I1194_032(w_1194_032, w_911_069, w_237_138);
  not1 I1194_157(w_1194_157, w_1011_314);
  not1 I1199_581(w_1199_581, w_749_660);
  not1 I1199_1953(w_1199_1955, w_1199_1954);
  nand2 I1199_1954(w_1199_1956, w_1199_1955, w_236_182);
  or2  I1199_1955(w_1199_1954, w_1199_1956, w_1199_1973);
  not1 I1199_1956(w_1199_1961, w_1199_1960);
  not1 I1199_1957(w_1199_1962, w_1199_1961);
  not1 I1199_1958(w_1199_1963, w_1199_1962);
  or2  I1199_1959(w_1199_1964, w_1012_353, w_1199_1963);
  and2 I1199_1960(w_1199_1965, w_1199_1964, w_783_1101);
  not1 I1199_1961(w_1199_1966, w_1199_1965);
  nand2 I1199_1962(w_1199_1967, w_1199_1966, w_784_448);
  nand2 I1199_1963(w_1199_1968, w_1199_1967, w_295_616);
  and2 I1199_1964(w_1199_1969, w_416_198, w_1199_1968);
  not1 I1199_1965(w_1199_1970, w_1199_1969);
  and2 I1199_1966(w_1199_1971, w_1199_1970, w_922_1533);
  not1 I1199_1967(w_1199_1960, w_1199_1954);
  and2 I1199_1968(w_1199_1973, w_127_372, w_1199_1971);
  not1 I1200_704(w_1200_704, w_189_010);
  not1 I1203_345(w_1203_345, w_912_120);
  and2 I1204_137(w_1204_137, w_713_146, w_399_191);
  and2 I1208_1034(w_1208_1034, w_1072_321, w_158_162);
  not1 I1209_041(w_1209_041, w_223_221);
  or2  I1212_003(w_1212_003, w_238_073, w_094_058);
  not1 I1212_232(w_1212_232, w_301_1225);
  not1 I1213_087(w_1213_087, w_105_1403);
  not1 I1213_239(w_1213_239, w_1013_326);
  or2  I1215_855(w_1215_855, w_651_352, w_682_148);
  or2  I1224_1447(w_1224_1447, w_932_294, w_074_1109);
  nand2 I1226_737(w_1226_737, w_366_011, w_400_067);
  or2  I1226_1459(w_1226_1459, w_593_207, w_686_073);
  or2  I1227_414(w_1227_414, w_544_100, w_609_034);
  and2 I1230_964(w_1230_966, w_066_007, w_1230_965);
  or2  I1230_965(w_1230_967, w_1230_966, w_563_905);
  nand2 I1230_966(w_1230_968, w_1230_967, w_010_376);
  not1 I1230_967(w_1230_969, w_1230_968);
  and2 I1230_968(w_1230_970, w_1227_414, w_1230_969);
  nand2 I1230_969(w_1230_965, w_1230_970, w_585_360);
  not1 I1231_107(w_1231_107, w_422_251);
  and2 I1231_150(w_1231_150, w_365_620, w_799_494);
  and2 I1235_950(w_1235_950, w_737_163, w_687_1614);
  nand2 I1235_1006(w_1235_1006, w_1181_634, w_273_350);
  or2  I1236_1603(w_1236_1603, w_154_124, w_613_092);
  and2 I1239_311(w_1239_311, w_630_083, w_1111_1175);
  nand2 I1239_502(w_1239_502, w_389_1252, w_1065_185);
  and2 I1240_471(w_1240_471, w_552_027, w_877_566);
  not1 I1244_049(w_1244_049, w_405_284);
  or2  I1246_814(w_1246_814, w_097_354, w_466_271);
  nand2 I1252_023(w_1252_023, w_099_677, w_752_789);
  not1 I1253_704(w_1253_704, w_674_050);
  and2 I1253_710(w_1253_710, w_903_455, w_963_263);
  and2 I1258_009(w_1258_009, w_957_171, w_835_622);
  or2  I1258_040(w_1258_040, w_436_667, w_968_263);
  or2  I1259_894(w_1259_894, w_676_349, w_1231_107);
  or2  I1267_451(w_1267_451, w_627_1504, w_033_730);
  and2 I1270_723(w_1270_723, w_842_151, w_549_244);
  nand2 I1274_815(w_1274_815, w_866_1044, w_001_127);
  nand2 I1275_1431(w_1275_1433, w_1148_133, w_1275_1432);
  not1 I1275_1432(w_1275_1434, w_1275_1433);
  or2  I1275_1433(w_1275_1435, w_1275_1434, w_641_262);
  nand2 I1275_1434(w_1275_1436, w_1275_1435, w_1275_1456);
  not1 I1275_1435(w_1275_1437, w_1275_1436);
  nand2 I1275_1436(w_1275_1438, w_1275_1437, w_249_123);
  nand2 I1275_1437(w_1275_1439, w_968_742, w_1275_1438);
  not1 I1275_1438(w_1275_1440, w_1275_1439);
  nand2 I1275_1439(w_1275_1432, w_1275_1440, w_862_052);
  and2 I1275_1440(w_1275_1445, w_1275_1444, w_504_152);
  and2 I1275_1441(w_1275_1446, w_1275_1445, w_063_1040);
  nand2 I1275_1442(w_1275_1447, w_942_113, w_1275_1446);
  or2  I1275_1443(w_1275_1448, w_1275_1447, w_011_702);
  not1 I1275_1444(w_1275_1449, w_1275_1448);
  not1 I1275_1445(w_1275_1450, w_1275_1449);
  or2  I1275_1446(w_1275_1451, w_1275_1450, w_1246_814);
  nand2 I1275_1447(w_1275_1452, w_1275_1451, w_626_1103);
  or2  I1275_1448(w_1275_1453, w_421_269, w_1275_1452);
  not1 I1275_1449(w_1275_1454, w_1275_1453);
  not1 I1275_1450(w_1275_1444, w_1275_1436);
  and2 I1275_1451(w_1275_1456, w_135_160, w_1275_1454);
  or2  I1276_796(w_1276_796, w_169_1320, w_419_087);
  nand2 I1281_436(w_1281_436, w_365_536, w_716_135);
  nand2 I1288_1601(w_1288_1603, w_1288_1602, w_1033_020);
  and2 I1288_1602(w_1288_1604, w_1288_1603, w_1288_1622);
  nand2 I1288_1603(w_1288_1605, w_576_511, w_1288_1604);
  not1 I1288_1604(w_1288_1606, w_1288_1605);
  not1 I1288_1605(w_1288_1607, w_1288_1606);
  not1 I1288_1606(w_1288_1602, w_1288_1607);
  or2  I1288_1607(w_1288_1612, w_658_866, w_1288_1611);
  and2 I1288_1608(w_1288_1613, w_1288_1612, w_408_011);
  not1 I1288_1609(w_1288_1614, w_1288_1613);
  and2 I1288_1610(w_1288_1615, w_1288_1614, w_852_269);
  and2 I1288_1611(w_1288_1616, w_1288_1615, w_1142_154);
  nand2 I1288_1612(w_1288_1617, w_1288_1616, w_1253_710);
  nand2 I1288_1613(w_1288_1618, w_1288_1617, w_866_722);
  and2 I1288_1614(w_1288_1619, w_890_822, w_1288_1618);
  or2  I1288_1615(w_1288_1620, w_543_374, w_1288_1619);
  not1 I1288_1616(w_1288_1611, w_1288_1604);
  and2 I1288_1617(w_1288_1622, w_722_1277, w_1288_1620);
  not1 I1289_284(w_1289_284, w_424_002);
  nand2 I1289_456(w_1289_457, w_1289_456, w_620_074);
  not1 I1289_457(w_1289_458, w_1289_457);
  nand2 I1289_458(w_1289_459, w_1289_458, w_549_222);
  or2  I1289_459(w_1289_460, w_1289_459, w_036_355);
  not1 I1289_460(w_1289_461, w_1289_460);
  nand2 I1289_461(w_1289_462, w_860_1045, w_1289_461);
  and2 I1289_462(w_1289_463, w_1289_462, w_606_070);
  or2  I1289_463(w_1289_456, w_326_737, w_1289_463);
  not1 I1293_1762(w_1293_1762, w_1239_311);
  or2  I1297_202(w_1297_202, w_1064_040, w_1018_633);
  and2 I1298_517(w_1298_519, w_1298_518, w_258_413);
  or2  I1298_518(w_1298_520, w_113_708, w_1298_519);
  and2 I1298_519(w_1298_518, w_1298_529, w_1298_520);
  nand2 I1298_520(w_1298_525, w_1298_524, w_978_267);
  nand2 I1298_521(w_1298_526, w_310_019, w_1298_525);
  or2  I1298_522(w_1298_527, w_1298_526, w_855_946);
  not1 I1298_523(w_1298_524, w_1298_518);
  and2 I1298_524(w_1298_529, w_1235_950, w_1298_527);
  and2 I1299_668(w_1299_668, w_1289_284, w_088_279);
  and2 I1301_098(w_1301_098, w_600_523, w_309_086);
  or2  I1303_222(w_1303_222, w_673_061, w_704_087);
  and2 I1304_708(w_1304_708, w_1104_019, w_144_703);
  or2  I1305_025(w_1305_025, w_962_105, w_1065_229);
  nand2 I1305_036(w_1305_036, w_1200_704, w_365_198);
  or2  I1308_360(w_1308_362, w_1308_361, w_1308_384);
  not1 I1308_361(w_1308_363, w_1308_362);
  not1 I1308_362(w_1308_364, w_1308_363);
  nand2 I1308_363(w_1308_365, w_1308_364, w_332_063);
  not1 I1308_364(w_1308_366, w_1308_365);
  nand2 I1308_365(w_1308_367, w_1308_366, w_877_632);
  not1 I1308_366(w_1308_368, w_1308_367);
  and2 I1308_367(w_1308_369, w_1308_368, w_1117_515);
  nand2 I1308_368(w_1308_370, w_1308_369, w_1212_003);
  not1 I1308_369(w_1308_371, w_1308_370);
  or2  I1308_370(w_1308_372, w_1308_371, w_204_1002);
  not1 I1308_371(w_1308_361, w_1308_372);
  or2  I1308_372(w_1308_377, w_1308_376, w_107_888);
  not1 I1308_373(w_1308_378, w_1308_377);
  and2 I1308_374(w_1308_379, w_326_1155, w_1308_378);
  and2 I1308_375(w_1308_380, w_1308_379, w_1203_345);
  not1 I1308_376(w_1308_381, w_1308_380);
  and2 I1308_377(w_1308_382, w_633_068, w_1308_381);
  not1 I1308_378(w_1308_376, w_1308_362);
  and2 I1308_379(w_1308_384, w_882_384, w_1308_382);
  nand2 I1312_968(w_1312_970, w_1312_969, w_030_542);
  or2  I1312_969(w_1312_971, w_1312_970, w_492_043);
  not1 I1312_970(w_1312_972, w_1312_971);
  not1 I1312_971(w_1312_973, w_1312_972);
  nand2 I1312_972(w_1312_974, w_889_097, w_1312_973);
  not1 I1312_973(w_1312_975, w_1312_974);
  and2 I1312_974(w_1312_976, w_1312_975, w_270_265);
  nand2 I1312_975(w_1312_977, w_1312_976, w_156_447);
  and2 I1312_976(w_1312_978, w_726_1725, w_1312_977);
  and2 I1312_977(w_1312_979, w_1312_978, w_1005_1726);
  or2  I1312_978(w_1312_980, w_889_030, w_1312_979);
  or2  I1312_979(w_1312_969, w_1312_988, w_1312_980);
  and2 I1312_980(w_1312_985, w_1312_984, w_530_1605);
  or2  I1312_981(w_1312_986, w_1312_985, w_614_388);
  not1 I1312_982(w_1312_984, w_1312_969);
  and2 I1312_983(w_1312_988, w_908_1300, w_1312_986);
  not1 I1316_035(w_1316_035, w_141_542);
  or2  I1320_000(w_1320_000, w_428_864, w_622_749);
  and2 I1321_169(w_1321_169, w_805_553, w_004_731);
  and2 I1329_047(w_1329_047, w_697_939, w_1133_1692);
  nand2 I1329_157(w_1329_157, w_635_326, w_1066_974);
  nand2 I1329_196(w_1329_196, w_225_962, w_644_837);
  nand2 I1330_429(w_1330_429, w_503_023, w_819_177);
  nand2 I1331_343(w_1331_343, w_067_019, w_182_439);
  nand2 I1335_651(w_1335_651, w_1213_087, w_1208_1034);
  not1 I1339_1486(w_1339_1486, w_390_434);
  or2  I1354_916(w_1354_916, w_417_456, w_981_087);
  and2 I1362_599(w_1362_599, w_132_007, w_482_410);
  and2 I1363_168(w_1363_168, w_336_577, w_619_033);
  nand2 I1367_1256(w_1367_1256, w_234_011, w_766_241);
  and2 I1369_038(w_1369_038, w_521_852, w_458_1066);
  or2  I1375_1357(w_1375_1357, w_1236_1603, w_893_056);
  not1 I1376_518(w_1376_518, w_665_335);
  or2  I1378_503(w_1378_503, w_694_687, w_122_082);
  and2 I1380_542(w_1380_542, w_119_400, w_640_710);
  and2 I1381_336(w_1381_336, w_485_176, w_951_471);
  or2  I1391_245(w_1391_245, w_1047_1404, w_1363_168);
  or2  I1392_360(w_1392_360, w_915_948, w_324_742);
  or2  I1395_110(w_1395_110, w_779_1214, w_1274_815);
  nand2 I1396_1004(w_1396_1004, w_376_677, w_912_152);
  and2 I1399_334(w_1399_334, w_1258_009, w_546_078);
  not1 I1400_522(w_1400_522, w_1088_775);
  and2 I1403_125(w_1403_125, w_199_127, w_1331_343);
  and2 I1410_066(w_1410_066, w_651_1483, w_334_261);
  not1 I1410_086(w_1410_086, w_248_024);
  and2 I1422_539(w_1422_541, w_342_1028, w_1422_540);
  not1 I1422_540(w_1422_542, w_1422_541);
  or2  I1422_541(w_1422_543, w_1422_542, w_411_668);
  nand2 I1422_542(w_1422_544, w_1422_543, w_370_1459);
  or2  I1422_543(w_1422_540, w_1422_544, w_051_127);
  or2  I1423_461(w_1423_463, w_1423_462, w_116_386);
  or2  I1423_462(w_1423_464, w_1423_463, w_233_083);
  and2 I1423_463(w_1423_465, w_027_303, w_1423_464);
  not1 I1423_464(w_1423_466, w_1423_465);
  not1 I1423_465(w_1423_467, w_1423_466);
  and2 I1423_466(w_1423_468, w_134_477, w_1423_467);
  and2 I1423_467(w_1423_469, w_1423_468, w_683_161);
  nand2 I1423_468(w_1423_470, w_706_1392, w_1423_469);
  or2  I1423_469(w_1423_471, w_1069_285, w_1423_470);
  and2 I1423_470(w_1423_472, w_1423_471, w_1403_125);
  not1 I1423_471(w_1423_462, w_1423_472);
  nand2 I1427_403(w_1427_403, w_1301_098, w_251_204);
  and2 I1428_144(w_1428_144, w_1095_044, w_568_596);
  or2  I1429_723(w_1429_723, w_508_018, w_1281_436);
  nand2 I1433_189(w_1433_189, w_1226_1459, w_905_262);
  not1 I1440_698(w_1440_698, w_811_1552);
  nand2 I1446_545(w_1446_545, w_1109_060, w_498_507);
  nand2 I1449_388(w_1449_388, w_716_416, w_932_853);
  nand2 I1449_428(w_1449_428, w_1410_066, w_810_824);
  or2  I1449_505(w_1449_507, w_1165_045, w_1449_506);
  or2  I1449_506(w_1449_508, w_832_266, w_1449_507);
  nand2 I1449_507(w_1449_509, w_105_1248, w_1449_508);
  or2  I1449_508(w_1449_506, w_1449_509, w_555_1335);
  or2  I1454_158(w_1454_158, w_781_001, w_796_1672);
  and2 I1455_105(w_1455_105, w_355_213, w_388_339);
  and2 I1463_378(w_1463_378, w_762_873, w_1400_522);
  not1 I1463_482(w_1463_482, w_449_1041);
  nand2 I1468_475(w_1468_475, w_152_177, w_446_752);
  and2 I1486_226(w_1486_226, w_980_107, w_257_1467);
  nand2 I1492_357(w_1492_357, w_910_116, w_1056_111);
  nand2 I1494_332(w_1494_332, w_578_425, w_1157_360);
  and2 I1496_083(w_1496_083, w_704_803, w_099_140);
  and2 I1502_1051(w_1502_1051, w_1244_049, w_768_099);
  nand2 I1503_257(w_1503_257, w_591_762, w_174_742);
  or2  I1505_029(w_1505_029, w_886_088, w_1399_334);
  and2 I1510_151(w_1510_151, w_855_166, w_280_365);
  and2 I1511_527(w_1511_527, w_677_132, w_518_204);
  or2  I1513_018(w_1513_018, w_810_754, w_259_081);
  and2 I1524_069(w_1524_069, w_548_843, w_415_058);
  or2  I1529_1173(w_1529_1173, w_683_238, w_1212_232);
  and2 I1530_672(w_1530_672, w_248_147, w_1492_357);
  not1 I1534_349(w_1534_349, w_1097_525);
  not1 I1538_208(w_1538_208, w_398_086);
  or2  I1539_021(w_1539_021, w_1069_553, w_1305_025);
  or2  I1542_076(w_1542_076, w_907_426, w_062_072);
  and2 I1549_655(w_1549_655, w_212_762, w_1017_222);
  or2  I1550_140(w_1550_140, w_621_268, w_381_531);
  not1 I1560_137(w_1560_137, w_1169_327);
  or2  I1560_289(w_1560_289, w_1235_1006, w_559_669);
  nand2 I1561_166(w_1561_166, w_700_106, w_413_194);
  not1 I1563_104(w_1563_104, w_637_508);
  nand2 I1577_015(w_1577_015, w_885_1687, w_1194_032);
  nand2 I1578_109(w_1578_109, w_334_567, w_147_030);
  nand2 I1579_1707(w_1579_1709, w_1579_1708, w_1213_239);
  nand2 I1579_1708(w_1579_1710, w_1579_1709, w_1354_916);
  not1 I1579_1709(w_1579_1711, w_1579_1710);
  or2  I1579_1710(w_1579_1712, w_1579_1711, w_1226_737);
  nand2 I1579_1711(w_1579_1713, w_1579_1712, w_1258_040);
  and2 I1579_1712(w_1579_1714, w_1446_545, w_1579_1713);
  and2 I1579_1713(w_1579_1715, w_1579_1714, w_502_002);
  and2 I1579_1714(w_1579_1708, w_1579_1715, w_662_540);
  not1 I1580_224(w_1580_224, w_1173_1388);
  nand2 I1586_998(w_1586_998, w_616_1323, w_1563_104);
  or2  I1586_1357(w_1586_1357, w_916_732, w_294_813);
  not1 I1589_1440(w_1589_1440, w_723_166);
  or2  I1590_840(w_1590_840, w_648_062, w_1162_232);
  not1 I1594_878(w_1594_878, w_952_247);
  or2  I1596_216(w_1596_216, w_555_481, w_739_100);
  and2 I1598_1874(w_1598_1876, w_828_715, w_1598_1875);
  and2 I1598_1875(w_1598_1877, w_1598_1876, w_703_042);
  nand2 I1598_1876(w_1598_1878, w_1270_723, w_1598_1877);
  or2  I1598_1877(w_1598_1879, w_1598_1878, w_1376_518);
  not1 I1598_1878(w_1598_1880, w_1598_1879);
  nand2 I1598_1879(w_1598_1881, w_374_304, w_1598_1880);
  and2 I1598_1880(w_1598_1882, w_1598_1881, w_1093_049);
  not1 I1598_1881(w_1598_1883, w_1598_1882);
  and2 I1598_1882(w_1598_1884, w_121_723, w_1598_1883);
  nand2 I1598_1883(w_1598_1885, w_1502_1051, w_1598_1884);
  not1 I1598_1884(w_1598_1875, w_1598_1885);
  not1 I1601_112(w_1601_114, w_1601_113);
  or2  I1601_113(w_1601_115, w_1601_127, w_1601_114);
  not1 I1601_114(w_1601_113, w_1601_115);
  nand2 I1601_115(w_1601_120, w_1601_119, w_466_103);
  or2  I1601_116(w_1601_121, w_1601_120, w_975_669);
  and2 I1601_117(w_1601_122, w_1601_121, w_1468_475);
  or2  I1601_118(w_1601_123, w_1601_122, w_1534_349);
  and2 I1601_119(w_1601_124, w_1601_123, w_1259_894);
  nand2 I1601_120(w_1601_125, w_1601_124, w_901_607);
  not1 I1601_121(w_1601_119, w_1601_115);
  and2 I1601_122(w_1601_127, w_1025_1532, w_1601_125);
  and2 I1603_907(w_1603_907, w_644_866, w_1183_177);
  not1 I1603_1223(w_1603_1223, w_847_251);
  nand2 I1603_1583(w_1603_1583, w_1224_1447, w_464_379);
  or2  I1605_144(w_1605_144, w_1455_105, w_759_359);
  and2 I1609_218(w_1609_218, w_1494_332, w_1578_109);
  nand2 I1615_1009(w_1615_1009, w_988_096, w_1589_1440);
  nand2 I1622_078(w_1622_078, w_523_021, w_1433_189);
  and2 I1629_026(w_1629_026, w_1034_506, w_1036_805);
  or2  I1635_431(w_1635_431, w_264_257, w_1524_069);
  or2  I1652_404(w_1652_404, w_1329_157, w_748_059);
  and2 I1656_1926(w_1656_1928, w_1381_336, w_1656_1927);
  not1 I1656_1927(w_1656_1929, w_1656_1928);
  not1 I1656_1928(w_1656_1930, w_1656_1929);
  and2 I1656_1929(w_1656_1927, w_1656_1930, w_924_311);
  and2 I1666_1996(w_1666_1998, w_1666_1997, w_1605_144);
  nand2 I1666_1997(w_1666_1999, w_1666_1998, w_267_329);
  and2 I1666_1998(w_1666_2000, w_1666_1999, w_921_020);
  nand2 I1666_1999(w_1666_2001, w_768_1574, w_1666_2000);
  or2  I1666_2000(w_1666_2002, w_1666_2016, w_1666_2001);
  nand2 I1666_2001(w_1666_2003, w_1666_2002, w_1622_078);
  nand2 I1666_2002(w_1666_2004, w_1666_2003, w_939_556);
  nand2 I1666_2003(w_1666_2005, w_773_106, w_1666_2004);
  nand2 I1666_2004(w_1666_2006, w_1652_404, w_1666_2005);
  and2 I1666_2005(w_1666_2007, w_1666_2006, w_493_430);
  and2 I1666_2006(w_1666_2008, w_1666_2007, w_1267_451);
  or2  I1666_2007(w_1666_1997, w_1666_2008, w_1510_151);
  nand2 I1666_2008(w_1666_2013, w_1666_2012, w_1088_842);
  and2 I1666_2009(w_1666_2014, w_676_1465, w_1666_2013);
  not1 I1666_2010(w_1666_2012, w_1666_2002);
  and2 I1666_2011(w_1666_2016, w_356_335, w_1666_2014);
  and2 I1673_151(w_1673_151, w_949_751, w_150_715);
  not1 I1687_828(w_1687_828, w_748_352);
  and2 I1688_1680(w_1688_1682, w_1688_1681, w_524_464);
  and2 I1688_1681(w_1688_1683, w_1688_1682, w_1530_672);
  or2  I1688_1682(w_1688_1684, w_1688_1683, w_712_634);
  not1 I1688_1683(w_1688_1685, w_1688_1684);
  nand2 I1688_1684(w_1688_1686, w_1688_1685, w_304_846);
  or2  I1688_1685(w_1688_1687, w_1688_1686, w_1316_035);
  or2  I1688_1686(w_1688_1688, w_1688_1687, w_1586_1357);
  or2  I1688_1687(w_1688_1681, w_058_038, w_1688_1688);
  and2 I1692_078(w_1692_078, w_1580_224, w_085_439);
  not1 I1692_765(w_1692_767, w_1692_766);
  and2 I1692_766(w_1692_768, w_1692_767, w_940_140);
  or2  I1692_767(w_1692_769, w_1692_782, w_1692_768);
  or2  I1692_768(w_1692_770, w_1692_769, w_068_030);
  nand2 I1692_769(w_1692_766, w_1692_770, w_461_171);
  or2  I1692_770(w_1692_775, w_1692_774, w_1239_502);
  or2  I1692_771(w_1692_776, w_1629_026, w_1692_775);
  not1 I1692_772(w_1692_777, w_1692_776);
  and2 I1692_773(w_1692_778, w_186_165, w_1692_777);
  and2 I1692_774(w_1692_779, w_1692_778, w_336_1630);
  not1 I1692_775(w_1692_780, w_1692_779);
  not1 I1692_776(w_1692_774, w_1692_769);
  and2 I1692_777(w_1692_782, w_1134_1163, w_1692_780);
  or2  I1701_010(w_1701_010, w_841_1480, w_687_540);
  nand2 I1716_1335(w_1716_1335, w_1561_166, w_500_891);
  nand2 I1721_407(w_1721_407, w_1692_078, w_831_1052);
  nand2 I1721_863(w_1721_863, w_1010_649, w_807_312);
  not1 I1726_437(w_1726_437, w_578_634);
  and2 I1727_092(w_1727_092, w_1549_655, w_1112_1168);
  not1 I1732_311(w_1732_311, w_171_654);
  not1 I1734_083(w_1734_083, w_1727_092);
  and2 I1754_1116(w_1754_1116, w_1449_428, w_103_1257);
  not1 I1755_243(w_1755_243, w_602_517);
  nand2 I1760_002(w_1760_002, w_1428_144, w_496_101);
  or2  I1760_054(w_1760_054, w_1078_045, w_1178_104);
  not1 I1774_625(w_1774_625, w_782_860);
  or2  I1777_499(w_1777_499, w_447_169, w_1429_723);
  and2 I1787_1409(w_1787_1409, w_1018_418, w_1050_082);
  or2  I1800_369(w_1800_369, w_1006_1160, w_1754_1116);
  and2 I1801_026(w_1801_026, w_1392_360, w_595_157);
  and2 I1806_215(w_1806_215, w_179_397, w_1166_032);
  or2  I1810_274(w_1810_274, w_809_122, w_209_1088);
  or2  I1811_265(w_1811_265, w_1330_429, w_773_045);
  not1 I1816_144(w_1816_144, w_027_407);
  nand2 I1818_358(w_1818_360, w_1818_359, w_256_622);
  nand2 I1818_359(w_1818_361, w_1594_878, w_1818_360);
  not1 I1818_360(w_1818_362, w_1818_361);
  nand2 I1818_361(w_1818_359, w_1818_362, w_1560_289);
  not1 I1819_036(w_1819_036, w_411_1244);
  not1 I1820_561(w_1820_561, w_849_242);
  and2 I1821_247(w_1821_249, w_1252_023, w_1821_248);
  nand2 I1821_248(w_1821_250, w_514_955, w_1821_249);
  nand2 I1821_249(w_1821_251, w_1821_250, w_1821_268);
  or2  I1821_250(w_1821_252, w_1821_251, w_054_544);
  and2 I1821_251(w_1821_253, w_819_190, w_1821_252);
  nand2 I1821_252(w_1821_248, w_1821_253, w_820_664);
  or2  I1821_253(w_1821_258, w_1821_257, w_352_672);
  not1 I1821_254(w_1821_259, w_1821_258);
  and2 I1821_255(w_1821_260, w_310_477, w_1821_259);
  and2 I1821_256(w_1821_261, w_1463_482, w_1821_260);
  not1 I1821_257(w_1821_262, w_1821_261);
  not1 I1821_258(w_1821_263, w_1821_262);
  not1 I1821_259(w_1821_264, w_1821_263);
  nand2 I1821_260(w_1821_265, w_1199_581, w_1821_264);
  and2 I1821_261(w_1821_266, w_1821_265, w_731_059);
  not1 I1821_262(w_1821_257, w_1821_251);
  and2 I1821_263(w_1821_268, w_790_1308, w_1821_266);
  nand2 I1824_1451(w_1824_1453, w_1824_1452, w_966_336);
  nand2 I1824_1452(w_1824_1454, w_1824_1453, w_1158_191);
  and2 I1824_1453(w_1824_1452, w_1586_998, w_1824_1454);
  or2  I1833_629(w_1833_629, w_829_391, w_638_432);
  not1 I1836_1756(w_1836_1758, w_1836_1757);
  nand2 I1836_1757(w_1836_1759, w_238_272, w_1836_1758);
  nand2 I1836_1758(w_1836_1760, w_1836_1759, w_1304_708);
  or2  I1836_1759(w_1836_1761, w_397_673, w_1836_1760);
  nand2 I1836_1760(w_1836_1762, w_1836_1761, w_286_076);
  not1 I1836_1761(w_1836_1763, w_1836_1762);
  and2 I1836_1762(w_1836_1764, w_1836_1763, w_1303_222);
  not1 I1836_1763(w_1836_1765, w_1836_1764);
  and2 I1836_1764(w_1836_1766, w_341_302, w_1836_1765);
  and2 I1836_1765(w_1836_1767, w_1836_1766, w_403_097);
  and2 I1836_1766(w_1836_1768, w_1836_1778, w_1836_1767);
  or2  I1836_1767(w_1836_1757, w_1836_1768, w_1819_036);
  not1 I1836_1768(w_1836_1773, w_1836_1772);
  or2  I1836_1769(w_1836_1774, w_975_392, w_1836_1773);
  or2  I1836_1770(w_1836_1775, w_1836_1774, w_781_1578);
  or2  I1836_1771(w_1836_1776, w_1609_218, w_1836_1775);
  not1 I1836_1772(w_1836_1772, w_1836_1768);
  and2 I1836_1773(w_1836_1778, w_1538_208, w_1836_1776);
  not1 I1848_116(w_1848_118, w_1848_117);
  not1 I1848_117(w_1848_119, w_1848_118);
  not1 I1848_118(w_1848_120, w_1848_119);
  not1 I1848_119(w_1848_117, w_1848_120);
  not1 I1871_787(w_1871_787, w_199_620);
  or2  I1873_820(w_1873_820, w_979_555, w_761_408);
  not1 I1885_477(w_1885_477, w_1038_1382);
  not1 I1890_797(w_1890_797, w_1168_039);
  nand2 I1891_031(w_1891_031, w_1049_021, w_1721_863);
  and2 I1904_1675(w_1904_1675, w_311_386, w_548_325);
  and2 I1905_377(w_1905_377, w_858_124, w_1505_029);
  not1 I1911_1095(w_1911_1097, w_1911_1096);
  not1 I1911_1096(w_1911_1098, w_1911_1097);
  nand2 I1911_1097(w_1911_1099, w_1801_026, w_1911_1098);
  nand2 I1911_1098(w_1911_1100, w_810_657, w_1911_1099);
  nand2 I1911_1099(w_1911_1101, w_1911_1100, w_798_611);
  nand2 I1911_1100(w_1911_1102, w_1911_1101, w_1503_257);
  or2  I1911_1101(w_1911_1103, w_1911_1102, w_510_177);
  not1 I1911_1102(w_1911_1104, w_1911_1103);
  or2  I1911_1103(w_1911_1105, w_051_992, w_1911_1104);
  nand2 I1911_1104(w_1911_1106, w_1687_828, w_1911_1105);
  not1 I1911_1105(w_1911_1107, w_1911_1106);
  or2  I1911_1106(w_1911_1096, w_1787_1409, w_1911_1107);
  not1 I1916_638(w_1916_638, w_890_411);
  not1 I1927_525(w_1927_525, w_1890_797);
  or2  I1937_085(w_1937_085, w_434_621, w_975_1237);
  and2 I1940_595(w_1940_595, w_1002_108, w_1004_487);
  not1 I1943_034(w_1943_034, w_545_1135);
  not1 I1964_004(w_1964_004, w_488_978);
  nand2 I1983_007(w_1983_007, w_1542_076, w_247_657);
  or2  I1986_071(w_1986_071, w_120_172, w_722_1323);
  not1 I1986_421(w_1986_421, w_1486_226);
  not1 I1990_1658(w_1990_1658, w_1367_1256);
  or2  I1994_186(w_1994_186, w_147_066, w_1983_007);
  not1 I1997_662(w_1997_662, w_442_1693);
  not1 I2000_000(w_2000_000, w_206_621);
  and2 I2000_001(w_2000_001, w_1811_265, w_1209_041);
  and2 I2000_002(w_2000_002, w_1603_1583, w_1131_656);
  and2 I2000_003(w_2000_003, w_1990_1658, w_222_411);
  or2  I2000_004(w_2000_004, w_334_650, w_1299_668);
  or2  I2000_005(w_2000_005, w_1560_137, w_1454_158);
  and2 I2000_006(w_2000_006, w_281_131, w_1590_840);
  nand2 I2000_007(w_2000_007, w_1335_651, w_401_544);
  or2  I2000_008(w_2000_008, w_1777_499, w_488_908);
  not1 I2000_009(w_2000_009, w_1820_561);
  and2 I2000_010(w_2000_010, w_042_009, w_493_157);
  nand2 I2000_011(w_2000_011, w_144_044, w_000_1704);
  not1 I2000_012(w_2000_012, w_1806_215);
  not1 I2000_013(w_2000_013, w_088_698);
  or2  I2000_014(w_2000_014, w_928_200, w_1940_595);
  nand2 I2000_015(w_2000_015, w_836_246, w_1716_1335);
  and2 I2000_016(w_2000_016, w_976_215, w_1496_083);
  or2  I2000_017(w_2000_017, w_1891_031, w_171_971);
  not1 I2000_018(w_2000_018, w_315_720);
  not1 I2000_019(w_2000_019, w_020_579);
  or2  I2000_020(w_2000_020, w_587_869, w_1321_169);
  not1 I2000_021(w_2000_021, w_601_471);
  not1 I2000_022(w_2000_022, w_532_410);
  not1 I2000_023(w_2000_023, w_1369_038);
  or2  I2000_024(w_2000_024, w_1045_096, w_790_894);
  or2  I2000_025(w_2000_025, w_467_1137, w_1916_638);
  and2 I2000_026(w_2000_026, w_991_026, w_1181_769);
  not1 I2000_027(w_2000_027, w_1035_002);
  or2  I2000_028(w_2000_028, w_1904_1675, w_1550_140);
  and2 I2000_029(w_2000_029, w_374_1496, w_1161_784);
  not1 I2000_030(w_2000_030, w_530_1263);
  nand2 I2000_031(w_2000_031, w_1927_525, w_1529_1173);
  not1 I2000_032(w_2000_032, w_1997_662);
  nand2 I2000_033(w_2000_033, w_987_771, w_362_293);
  and2 I2000_034(w_2000_034, w_1131_664, w_1339_1486);
  and2 I2000_035(w_2000_035, w_1596_216, w_139_1326);
  not1 I2000_036(w_2000_036, w_865_178);
  nand2 I2000_037(w_2000_037, w_001_921, w_1833_629);
  or2  I2000_038(w_2000_038, w_1760_054, w_1190_258);
  and2 I2000_039(w_2000_039, w_1539_021, w_1511_527);
  nand2 I2000_040(w_2000_040, w_1873_820, w_1375_1357);
  and2 I2000_041(w_2000_041, w_715_843, w_1732_311);
  and2 I2000_042(w_2000_042, w_1871_787, w_146_232);
  and2 I2000_043(w_2000_043, w_1097_1090, w_1734_083);
  not1 I2000_044(w_2000_044, w_1395_110);
  and2 I2000_045(w_2000_045, w_937_329, w_1885_477);
  or2  I2000_046(w_2000_046, w_1396_1004, w_1701_010);
  and2 I2000_047(w_2000_047, w_1076_206, w_1320_000);
  not1 I2000_048(w_2000_048, w_1053_806);
  not1 I2000_049(w_2000_049, w_1276_796);
  or2  I2000_050(w_2000_050, w_717_1608, w_1774_625);
  not1 I2000_051(w_2000_051, w_1057_865);
  or2  I2000_052(w_2000_052, w_100_610, w_379_781);
  nand2 I2000_053(w_2000_053, w_856_1410, w_595_321);
  nand2 I2000_054(w_2000_054, w_569_388, w_892_214);
  or2  I2000_055(w_2000_055, w_1035_074, w_1114_194);
  or2  I2000_056(w_2000_056, w_742_065, w_1986_071);
  not1 I2000_057(w_2000_057, w_1760_002);
  or2  I2000_058(w_2000_058, w_817_484, w_086_1269);
  not1 I2000_059(w_2000_059, w_465_050);
  or2  I2000_060(w_2000_060, w_1673_151, w_1240_471);
  and2 I2000_061(w_2000_061, w_1810_274, w_1816_144);
  nand2 I2000_062(w_2000_062, w_1204_137, w_1449_388);
  not1 I2000_063(w_2000_063, w_543_740);
  and2 I2000_064(w_2000_064, w_003_042, w_1192_779);
  nand2 I2000_065(w_2000_065, w_362_105, w_1126_121);
  nand2 I2000_066(w_2000_066, w_1943_034, w_548_636);
  nand2 I2000_067(w_2000_067, w_141_046, w_771_455);
  and2 I2000_068(w_2000_068, w_940_013, w_463_144);
  not1 I2000_069(w_2000_069, w_264_181);
  and2 I2000_070(w_2000_070, w_808_986, w_1380_542);
  and2 I2000_071(w_2000_071, w_925_784, w_068_062);
  not1 I2000_072(w_2000_072, w_1194_157);
  or2  I2000_073(w_2000_073, w_1137_216, w_046_254);
  nand2 I2000_074(w_2000_074, w_187_075, w_275_490);
  or2  I2000_075(w_2000_075, w_1215_855, w_1905_377);
  not1 I2000_076(w_2000_076, w_169_507);
  not1 I2000_077(w_2000_077, w_1329_047);
  nand2 I2000_078(w_2000_078, w_844_323, w_1964_004);
  nand2 I2000_079(w_2000_079, w_1603_1223, w_1937_085);
  and2 I2000_080(w_2000_080, w_1427_403, w_1118_533);
  or2  I2000_081(w_2000_081, w_1305_036, w_1012_147);
  and2 I2000_082(w_2000_082, w_579_1003, w_841_642);
  or2  I2000_083(w_2000_083, w_1362_599, w_371_092);
  not1 I2000_084(w_2000_084, w_1410_086);
  not1 I2000_085(w_2000_085, w_1726_437);
  or2  I2000_086(w_2000_086, w_1329_196, w_1603_907);
  or2  I2000_087(w_2000_087, w_1030_528, w_1635_431);
  not1 I2000_088(w_2000_088, w_1293_1762);
  nand2 I2000_089(w_2000_089, w_1440_698, w_118_795);
  nand2 I2000_090(w_2000_090, w_761_029, w_1253_704);
  and2 I2000_091(w_2000_091, w_297_083, w_1994_186);
  or2  I2000_092(w_2000_092, w_1721_407, w_546_065);
  and2 I2000_093(w_2000_093, w_149_309, w_369_1531);
  not1 I2000_094(w_2000_094, w_004_1447);
  or2  I2000_095(w_2000_095, w_1297_202, w_516_317);
  nand2 I2000_096(w_2000_096, w_634_237, w_150_1395);
  not1 I2000_097(w_2000_097, w_1755_243);
  not1 I2000_098(w_2000_098, w_053_077);
  and2 I2000_099(w_2000_099, w_591_300, w_397_1350);
  not1 I2000_100(w_2000_100, w_1800_369);
  and2 I2000_101(w_2000_101, w_461_047, w_1231_150);
  and2 I2000_102(w_2000_102, w_678_781, w_1577_015);
  or2  I2000_103(w_2000_103, w_1019_850, w_1391_245);
  and2 I2000_104(w_2000_104, w_1139_1355, w_1108_010);
  or2  I2000_105(w_2000_105, w_1513_018, w_713_104);
  not1 I2000_106(w_2000_106, w_1463_378);
  and2 I2000_107(w_2000_107, w_1615_1009, w_864_076);
  and2 I2000_108(w_2000_108, w_096_195, w_860_017);
  or2  I2000_109(w_2000_109, w_790_373, w_1986_421);
  and2 I2000_110(w_2000_110, w_1378_503, w_273_869);

  initial begin
    $get_module_info();
  end
endmodule

// ****** Combined Logic Module Defination ******

// ****** TestBench Module Defination ******

/*
module tb();
  wire  w_000_000, w_000_001, w_000_002, w_000_003, w_000_004, w_000_005, w_000_006, w_000_007, w_000_008, w_000_009, w_000_010, w_000_011, w_000_012, w_000_013, w_000_014, w_000_015, w_000_016, w_000_017, w_000_018, w_000_019, w_000_020, w_000_021, w_000_022, w_000_023, w_000_024, w_000_025, w_000_026, w_000_027, w_000_028, w_000_029, w_000_030, w_000_031, w_000_032, w_000_033, w_000_034, w_000_035, w_000_036, w_000_037, w_000_038, w_000_039, w_000_040, w_000_041, w_000_042, w_000_043, w_000_044, w_000_045, w_000_046, w_000_047, w_000_048, w_000_049, w_000_050, w_000_051, w_000_052, w_000_053, w_000_054, w_000_055, w_000_056, w_000_057, w_000_058, w_000_059, w_000_060, w_000_061, w_000_062, w_000_063, w_000_065, w_000_066, w_000_067, w_000_068, w_000_069, w_000_070, w_000_071, w_000_072, w_000_073, w_000_074, w_000_075, w_000_076, w_000_077, w_000_078, w_000_079, w_000_080, w_000_081, w_000_082, w_000_083, w_000_084, w_000_085, w_000_086, w_000_087, w_000_088, w_000_089, w_000_090, w_000_091, w_000_092, w_000_093, w_000_094, w_000_095, w_000_096, w_000_097, w_000_098, w_000_099, w_000_100, w_000_101, w_000_102, w_000_103, w_000_104, w_000_105, w_000_106, w_000_107, w_000_108, w_000_109, w_000_110, w_000_111, w_000_112, w_000_113, w_000_114, w_000_115, w_000_116, w_000_117, w_000_118, w_000_119, w_000_120, w_000_121, w_000_122, w_000_123, w_000_124, w_000_125, w_000_126, w_000_127, w_000_128, w_000_129, w_000_130, w_000_131, w_000_132, w_000_133, w_000_134, w_000_135, w_000_136, w_000_137, w_000_138, w_000_139, w_000_140, w_000_141, w_000_142, w_000_143, w_000_144, w_000_145, w_000_146, w_000_147, w_000_148, w_000_149, w_000_150, w_000_151, w_000_152, w_000_153, w_000_154, w_000_155, w_000_156, w_000_157, w_000_158, w_000_159, w_000_160, w_000_161, w_000_162, w_000_163, w_000_164, w_000_165, w_000_166, w_000_167, w_000_168, w_000_169, w_000_170, w_000_171, w_000_172, w_000_173, w_000_174, w_000_175, w_000_176, w_000_177, w_000_178, w_000_179, w_000_180, w_000_181, w_000_182, w_000_183, w_000_184, w_000_185, w_000_186, w_000_187, w_000_188, w_000_189, w_000_190, w_000_191, w_000_192, w_000_193, w_000_194, w_000_195, w_000_196, w_000_197, w_000_198, w_000_199, w_000_200, w_000_201, w_000_202, w_000_203, w_000_204, w_000_205, w_000_206, w_000_207, w_000_208, w_000_209, w_000_210, w_000_211, w_000_212, w_000_213, w_000_214, w_000_215, w_000_216, w_000_217, w_000_218, w_000_219, w_000_220, w_000_221, w_000_222, w_000_223, w_000_224, w_000_225, w_000_226, w_000_227, w_000_228, w_000_229, w_000_230, w_000_231, w_000_232, w_000_233, w_000_234, w_000_235, w_000_236, w_000_237, w_000_238, w_000_239, w_000_240, w_000_241, w_000_242, w_000_243, w_000_244, w_000_245, w_000_246, w_000_247, w_000_248, w_000_249, w_000_250, w_000_251, w_000_252, w_000_253, w_000_254, w_000_255, w_000_256, w_000_257, w_000_258, w_000_259, w_000_260, w_000_261, w_000_262, w_000_263, w_000_264, w_000_265, w_000_266, w_000_267, w_000_268, w_000_269, w_000_270, w_000_271, w_000_272, w_000_273, w_000_274, w_000_275, w_000_276, w_000_277, w_000_278, w_000_279, w_000_280, w_000_281, w_000_282, w_000_283, w_000_284, w_000_285, w_000_286, w_000_287, w_000_289, w_000_290, w_000_291, w_000_292, w_000_293, w_000_294, w_000_295, w_000_296, w_000_297, w_000_298, w_000_299, w_000_300, w_000_301, w_000_302, w_000_303, w_000_304, w_000_305, w_000_306, w_000_307, w_000_308, w_000_309, w_000_310, w_000_311, w_000_312, w_000_313, w_000_314, w_000_315, w_000_316, w_000_317, w_000_318, w_000_319, w_000_320, w_000_321, w_000_322, w_000_323, w_000_324, w_000_325, w_000_326, w_000_327, w_000_328, w_000_329, w_000_330, w_000_331, w_000_332, w_000_333, w_000_334, w_000_335, w_000_336, w_000_337, w_000_338, w_000_339, w_000_340, w_000_341, w_000_342, w_000_343, w_000_344, w_000_345, w_000_346, w_000_347, w_000_348, w_000_349, w_000_350, w_000_351, w_000_352, w_000_353, w_000_354, w_000_355, w_000_356, w_000_357, w_000_358, w_000_359, w_000_360, w_000_361, w_000_362, w_000_363, w_000_364, w_000_365, w_000_366, w_000_367, w_000_368, w_000_369, w_000_370, w_000_371, w_000_372, w_000_373, w_000_374, w_000_375, w_000_376, w_000_377, w_000_378, w_000_379, w_000_380, w_000_381, w_000_382, w_000_383, w_000_384, w_000_385, w_000_386, w_000_387, w_000_388, w_000_389, w_000_390, w_000_391, w_000_392, w_000_393, w_000_394, w_000_395, w_000_396, w_000_397, w_000_398, w_000_399, w_000_400, w_000_401, w_000_402, w_000_403, w_000_404, w_000_405, w_000_406, w_000_407, w_000_408, w_000_409, w_000_410, w_000_411, w_000_412, w_000_413, w_000_414, w_000_415, w_000_416, w_000_417, w_000_418, w_000_419, w_000_420, w_000_421, w_000_422, w_000_423, w_000_424, w_000_425, w_000_426, w_000_427, w_000_428, w_000_429, w_000_430, w_000_431, w_000_432, w_000_433, w_000_434, w_000_435, w_000_436, w_000_437, w_000_438, w_000_439, w_000_440, w_000_441, w_000_442, w_000_443, w_000_444, w_000_445, w_000_446, w_000_447, w_000_448, w_000_449, w_000_450, w_000_451, w_000_452, w_000_453, w_000_454, w_000_455, w_000_456, w_000_457, w_000_458, w_000_459, w_000_460, w_000_461, w_000_462, w_000_463, w_000_464, w_000_465, w_000_466, w_000_467, w_000_468, w_000_469, w_000_470, w_000_471, w_000_472, w_000_473, w_000_474, w_000_475, w_000_476, w_000_477, w_000_478, w_000_479, w_000_480, w_000_481, w_000_482, w_000_483, w_000_484, w_000_485, w_000_486, w_000_487, w_000_488, w_000_489, w_000_490, w_000_491, w_000_492, w_000_493, w_000_494, w_000_495, w_000_496, w_000_498, w_000_499, w_000_500, w_000_501, w_000_502, w_000_503, w_000_504, w_000_505, w_000_506, w_000_507, w_000_508, w_000_509, w_000_510, w_000_511, w_000_512, w_000_513, w_000_514, w_000_515, w_000_516, w_000_517, w_000_518, w_000_519, w_000_520, w_000_521, w_000_522, w_000_523, w_000_524, w_000_525, w_000_526, w_000_527, w_000_528, w_000_529, w_000_530, w_000_531, w_000_532, w_000_533, w_000_534, w_000_535, w_000_536, w_000_537, w_000_538, w_000_539, w_000_540, w_000_541, w_000_542, w_000_543, w_000_544, w_000_545, w_000_546, w_000_547, w_000_548, w_000_549, w_000_550, w_000_551, w_000_552, w_000_553, w_000_554, w_000_555, w_000_556, w_000_557, w_000_558, w_000_559, w_000_560, w_000_561, w_000_562, w_000_563, w_000_564, w_000_565, w_000_566, w_000_567, w_000_568, w_000_569, w_000_570, w_000_571, w_000_572, w_000_573, w_000_575, w_000_576, w_000_577, w_000_578, w_000_579, w_000_580, w_000_581, w_000_582, w_000_583, w_000_584, w_000_585, w_000_586, w_000_587, w_000_588, w_000_589, w_000_590, w_000_591, w_000_592, w_000_593, w_000_594, w_000_595, w_000_596, w_000_597, w_000_598, w_000_599, w_000_600, w_000_601, w_000_602, w_000_603, w_000_604, w_000_605, w_000_606, w_000_607, w_000_608, w_000_609, w_000_610, w_000_611, w_000_612, w_000_613, w_000_614, w_000_615, w_000_616, w_000_617, w_000_618, w_000_619, w_000_620, w_000_621, w_000_622, w_000_623, w_000_624, w_000_625, w_000_626, w_000_627, w_000_628, w_000_629, w_000_630, w_000_631, w_000_632, w_000_633, w_000_634, w_000_635, w_000_636, w_000_638, w_000_639, w_000_640, w_000_641, w_000_643, w_000_644, w_000_645, w_000_646, w_000_647, w_000_648, w_000_649, w_000_650, w_000_651, w_000_652, w_000_653, w_000_654, w_000_655, w_000_656, w_000_657, w_000_658, w_000_659, w_000_660, w_000_661, w_000_662, w_000_663, w_000_664, w_000_665, w_000_667, w_000_668, w_000_669, w_000_670, w_000_671, w_000_672, w_000_673, w_000_674, w_000_675, w_000_676, w_000_677, w_000_678, w_000_679, w_000_680, w_000_681, w_000_682, w_000_683, w_000_684, w_000_685, w_000_686, w_000_687, w_000_688, w_000_689, w_000_690, w_000_691, w_000_692, w_000_693, w_000_694, w_000_695, w_000_696, w_000_697, w_000_698, w_000_699, w_000_700, w_000_701, w_000_702, w_000_703, w_000_704, w_000_705, w_000_706, w_000_707, w_000_708, w_000_709, w_000_710, w_000_711, w_000_712, w_000_713, w_000_714, w_000_715, w_000_716, w_000_717, w_000_718, w_000_719, w_000_720, w_000_721, w_000_722, w_000_723, w_000_724, w_000_725, w_000_726, w_000_727, w_000_728, w_000_729, w_000_730, w_000_731, w_000_732, w_000_733, w_000_734, w_000_735, w_000_736, w_000_737, w_000_738, w_000_739, w_000_740, w_000_741, w_000_742, w_000_743, w_000_744, w_000_745, w_000_746, w_000_747, w_000_748, w_000_749, w_000_750, w_000_751, w_000_752, w_000_753, w_000_754, w_000_755, w_000_756, w_000_757, w_000_758, w_000_759, w_000_760, w_000_761, w_000_762, w_000_763, w_000_764, w_000_765, w_000_766, w_000_767, w_000_768, w_000_769, w_000_770, w_000_771, w_000_772, w_000_773, w_000_774, w_000_775, w_000_776, w_000_777, w_000_778, w_000_779, w_000_780, w_000_781, w_000_782, w_000_783, w_000_784, w_000_785, w_000_786, w_000_787, w_000_788, w_000_789, w_000_790, w_000_791, w_000_792, w_000_793, w_000_794, w_000_795, w_000_796, w_000_797, w_000_798, w_000_799, w_000_800, w_000_801, w_000_802, w_000_803, w_000_804, w_000_805, w_000_806, w_000_807, w_000_808, w_000_809, w_000_810, w_000_811, w_000_812, w_000_813, w_000_814, w_000_815, w_000_816, w_000_817, w_000_818, w_000_819, w_000_820, w_000_821, w_000_822, w_000_823, w_000_824, w_000_825, w_000_826, w_000_827, w_000_828, w_000_829, w_000_830, w_000_831, w_000_832, w_000_833, w_000_835, w_000_836, w_000_837, w_000_838, w_000_839, w_000_840, w_000_841, w_000_842, w_000_843, w_000_844, w_000_845, w_000_846, w_000_847, w_000_848, w_000_849, w_000_850, w_000_851, w_000_852, w_000_853, w_000_854, w_000_855, w_000_856, w_000_857, w_000_858, w_000_859, w_000_860, w_000_861, w_000_862, w_000_863, w_000_864, w_000_865, w_000_866, w_000_867, w_000_868, w_000_869, w_000_870, w_000_871, w_000_872, w_000_873, w_000_874, w_000_875, w_000_876, w_000_877, w_000_878, w_000_879, w_000_880, w_000_881, w_000_882, w_000_883, w_000_884, w_000_885, w_000_886, w_000_887, w_000_888, w_000_889, w_000_890, w_000_891, w_000_892, w_000_893, w_000_894, w_000_895, w_000_896, w_000_897, w_000_898, w_000_899, w_000_900, w_000_901, w_000_902, w_000_903, w_000_904, w_000_905, w_000_906, w_000_907, w_000_908, w_000_909, w_000_910, w_000_911, w_000_912, w_000_913, w_000_914, w_000_915, w_000_916, w_000_917, w_000_918, w_000_919, w_000_920, w_000_921, w_000_922, w_000_923, w_000_924, w_000_925, w_000_926, w_000_927, w_000_928, w_000_929, w_000_930, w_000_931, w_000_932, w_000_933, w_000_935, w_000_936, w_000_937, w_000_938, w_000_939, w_000_940, w_000_941, w_000_942, w_000_943, w_000_944, w_000_945, w_000_946, w_000_947, w_000_948, w_000_949, w_000_950, w_000_951, w_000_952, w_000_953, w_000_954, w_000_955, w_000_956, w_000_957, w_000_958, w_000_959, w_000_960, w_000_961, w_000_962, w_000_963, w_000_964, w_000_965, w_000_966, w_000_967, w_000_968, w_000_969, w_000_970, w_000_971, w_000_972, w_000_973, w_000_974, w_000_975, w_000_976, w_000_977, w_000_978, w_000_979, w_000_980, w_000_981, w_000_982, w_000_983, w_000_984, w_000_985, w_000_986, w_000_987, w_000_988, w_000_989, w_000_990, w_000_991, w_000_992, w_000_993, w_000_994, w_000_995, w_000_996, w_000_997, w_000_998, w_000_999, w_000_1000, w_000_1001, w_000_1002, w_000_1003, w_000_1004, w_000_1005, w_000_1006, w_000_1007, w_000_1008, w_000_1009, w_000_1010, w_000_1011, w_000_1012, w_000_1013, w_000_1014, w_000_1015, w_000_1016, w_000_1017, w_000_1018, w_000_1019, w_000_1020, w_000_1021, w_000_1022, w_000_1023, w_000_1024, w_000_1025, w_000_1026, w_000_1027, w_000_1028, w_000_1029, w_000_1030, w_000_1031, w_000_1032, w_000_1033, w_000_1034, w_000_1035, w_000_1036, w_000_1037, w_000_1038, w_000_1039, w_000_1040, w_000_1041, w_000_1042, w_000_1043, w_000_1044, w_000_1045, w_000_1046, w_000_1047, w_000_1048, w_000_1049, w_000_1050, w_000_1051, w_000_1052, w_000_1053, w_000_1054, w_000_1055, w_000_1056, w_000_1057, w_000_1058, w_000_1060, w_000_1061, w_000_1062, w_000_1063, w_000_1064, w_000_1065, w_000_1066, w_000_1067, w_000_1068, w_000_1069, w_000_1070, w_000_1071, w_000_1072, w_000_1073, w_000_1074, w_000_1075, w_000_1076, w_000_1077, w_000_1078, w_000_1079, w_000_1080, w_000_1081, w_000_1082, w_000_1083, w_000_1084, w_000_1085, w_000_1086, w_000_1087, w_000_1088, w_000_1089, w_000_1090, w_000_1091, w_000_1093, w_000_1094, w_000_1095, w_000_1096, w_000_1097, w_000_1098, w_000_1099, w_000_1101, w_000_1102, w_000_1103, w_000_1104, w_000_1105, w_000_1106, w_000_1107, w_000_1108, w_000_1109, w_000_1110, w_000_1111, w_000_1112, w_000_1113, w_000_1114, w_000_1115, w_000_1116, w_000_1117, w_000_1118, w_000_1119, w_000_1120, w_000_1121, w_000_1122, w_000_1123, w_000_1124, w_000_1125, w_000_1126, w_000_1127, w_000_1128, w_000_1129, w_000_1130, w_000_1131, w_000_1132, w_000_1133, w_000_1134, w_000_1136, w_000_1137, w_000_1138, w_000_1139, w_000_1140, w_000_1141, w_000_1142, w_000_1143, w_000_1144, w_000_1145, w_000_1146, w_000_1147, w_000_1148, w_000_1149, w_000_1150, w_000_1151, w_000_1152, w_000_1153, w_000_1154, w_000_1155, w_000_1156, w_000_1157, w_000_1158, w_000_1159, w_000_1160, w_000_1161, w_000_1162, w_000_1163, w_000_1165, w_000_1166, w_000_1168, w_000_1169, w_000_1171, w_000_1172, w_000_1173, w_000_1174, w_000_1175, w_000_1176, w_000_1177, w_000_1178, w_000_1179, w_000_1180, w_000_1181, w_000_1182, w_000_1183, w_000_1184, w_000_1185, w_000_1186, w_000_1187, w_000_1188, w_000_1189, w_000_1190, w_000_1191, w_000_1192, w_000_1193, w_000_1194, w_000_1195, w_000_1196, w_000_1197, w_000_1198, w_000_1199, w_000_1200, w_000_1201, w_000_1202, w_000_1203, w_000_1204, w_000_1205, w_000_1206, w_000_1207, w_000_1208, w_000_1209, w_000_1210, w_000_1211, w_000_1212, w_000_1213, w_000_1214, w_000_1215, w_000_1216, w_000_1217, w_000_1218, w_000_1219, w_000_1220, w_000_1221, w_000_1222, w_000_1223, w_000_1224, w_000_1225, w_000_1226, w_000_1227, w_000_1228, w_000_1229, w_000_1230, w_000_1231, w_000_1232, w_000_1233, w_000_1234, w_000_1235, w_000_1236, w_000_1237, w_000_1238, w_000_1239, w_000_1240, w_000_1241, w_000_1242, w_000_1243, w_000_1244, w_000_1245, w_000_1246, w_000_1247, w_000_1248, w_000_1249, w_000_1250, w_000_1251, w_000_1252, w_000_1253, w_000_1254, w_000_1255, w_000_1256, w_000_1257, w_000_1258, w_000_1259, w_000_1260, w_000_1261, w_000_1262, w_000_1264, w_000_1265, w_000_1266, w_000_1267, w_000_1268, w_000_1270, w_000_1271, w_000_1272, w_000_1274, w_000_1275, w_000_1276, w_000_1277, w_000_1278, w_000_1279, w_000_1282, w_000_1283, w_000_1284, w_000_1285, w_000_1286, w_000_1287, w_000_1288, w_000_1289, w_000_1290, w_000_1291, w_000_1293, w_000_1294, w_000_1295, w_000_1296, w_000_1297, w_000_1298, w_000_1299, w_000_1300, w_000_1301, w_000_1302, w_000_1303, w_000_1304, w_000_1305, w_000_1306, w_000_1307, w_000_1308, w_000_1309, w_000_1310, w_000_1311, w_000_1312, w_000_1313, w_000_1314, w_000_1315, w_000_1316, w_000_1317, w_000_1318, w_000_1320, w_000_1321, w_000_1322, w_000_1323, w_000_1324, w_000_1325, w_000_1326, w_000_1327, w_000_1328, w_000_1329, w_000_1330, w_000_1331, w_000_1332, w_000_1333, w_000_1334, w_000_1335, w_000_1338, w_000_1339, w_000_1340, w_000_1341, w_000_1342, w_000_1343, w_000_1344, w_000_1345, w_000_1346, w_000_1347, w_000_1348, w_000_1349, w_000_1350, w_000_1351, w_000_1352, w_000_1353, w_000_1354, w_000_1355, w_000_1356, w_000_1357, w_000_1358, w_000_1359, w_000_1360, w_000_1361, w_000_1362, w_000_1363, w_000_1365, w_000_1366, w_000_1367, w_000_1368, w_000_1369, w_000_1370, w_000_1371, w_000_1372, w_000_1373, w_000_1374, w_000_1375, w_000_1376, w_000_1377, w_000_1378, w_000_1379, w_000_1380, w_000_1381, w_000_1382, w_000_1383, w_000_1385, w_000_1386, w_000_1387, w_000_1388, w_000_1389, w_000_1390, w_000_1391, w_000_1392, w_000_1393, w_000_1394, w_000_1395, w_000_1396, w_000_1397, w_000_1398, w_000_1399, w_000_1400, w_000_1401, w_000_1402, w_000_1403, w_000_1405, w_000_1406, w_000_1407, w_000_1408, w_000_1409, w_000_1410, w_000_1411, w_000_1412, w_000_1413, w_000_1414, w_000_1415, w_000_1417, w_000_1418, w_000_1419, w_000_1421, w_000_1422, w_000_1423, w_000_1424, w_000_1425, w_000_1426, w_000_1427, w_000_1428, w_000_1429, w_000_1430, w_000_1431, w_000_1432, w_000_1433, w_000_1434, w_000_1435, w_000_1436, w_000_1437, w_000_1438, w_000_1439, w_000_1440, w_000_1441, w_000_1442, w_000_1443, w_000_1444, w_000_1445, w_000_1447, w_000_1448, w_000_1449, w_000_1450, w_000_1451, w_000_1452, w_000_1453, w_000_1454, w_000_1455, w_000_1457, w_000_1458, w_000_1459, w_000_1460, w_000_1461, w_000_1462, w_000_1463, w_000_1464, w_000_1465, w_000_1466, w_000_1467, w_000_1469, w_000_1470, w_000_1471, w_000_1472, w_000_1473, w_000_1474, w_000_1475, w_000_1476, w_000_1477, w_000_1478, w_000_1480, w_000_1481, w_000_1482, w_000_1483, w_000_1484, w_000_1485, w_000_1486, w_000_1487, w_000_1488, w_000_1489, w_000_1490, w_000_1491, w_000_1492, w_000_1493, w_000_1494, w_000_1495, w_000_1496, w_000_1497, w_000_1498, w_000_1499, w_000_1500, w_000_1501, w_000_1502, w_000_1503, w_000_1504, w_000_1505, w_000_1506, w_000_1507, w_000_1508, w_000_1509, w_000_1510, w_000_1511, w_000_1512, w_000_1513, w_000_1514, w_000_1515, w_000_1516, w_000_1518, w_000_1519, w_000_1520, w_000_1521, w_000_1522, w_000_1523, w_000_1524, w_000_1525, w_000_1526, w_000_1527, w_000_1528, w_000_1529, w_000_1530, w_000_1531, w_000_1532, w_000_1533, w_000_1534, w_000_1535, w_000_1536, w_000_1537, w_000_1538, w_000_1539, w_000_1540, w_000_1541, w_000_1542, w_000_1543, w_000_1544, w_000_1545, w_000_1546, w_000_1547, w_000_1548, w_000_1549, w_000_1550, w_000_1551, w_000_1552, w_000_1553, w_000_1554, w_000_1555, w_000_1556, w_000_1557, w_000_1558, w_000_1559, w_000_1560, w_000_1561, w_000_1562, w_000_1563, w_000_1564, w_000_1565, w_000_1566, w_000_1567, w_000_1568, w_000_1569, w_000_1570, w_000_1571, w_000_1572, w_000_1573, w_000_1574, w_000_1575, w_000_1576, w_000_1577, w_000_1578, w_000_1579, w_000_1580, w_000_1581, w_000_1583, w_000_1584, w_000_1585, w_000_1586, w_000_1587, w_000_1588, w_000_1589, w_000_1590, w_000_1591, w_000_1592, w_000_1593, w_000_1594, w_000_1595, w_000_1596, w_000_1597, w_000_1598, w_000_1599, w_000_1600, w_000_1601, w_000_1602, w_000_1603, w_000_1604, w_000_1605, w_000_1606, w_000_1607, w_000_1608, w_000_1609, w_000_1610, w_000_1611, w_000_1612, w_000_1613, w_000_1614, w_000_1615, w_000_1616, w_000_1617, w_000_1618, w_000_1619, w_000_1620, w_000_1621, w_000_1622, w_000_1623, w_000_1624, w_000_1625, w_000_1626, w_000_1627, w_000_1628, w_000_1629, w_000_1630, w_000_1631, w_000_1632, w_000_1633, w_000_1634, w_000_1635, w_000_1636, w_000_1637, w_000_1638, w_000_1639, w_000_1640, w_000_1641, w_000_1642, w_000_1643, w_000_1644, w_000_1645, w_000_1646, w_000_1647, w_000_1648, w_000_1649, w_000_1650, w_000_1651, w_000_1652, w_000_1653, w_000_1654, w_000_1655, w_000_1656, w_000_1657, w_000_1658, w_000_1659, w_000_1660, w_000_1661, w_000_1662, w_000_1663, w_000_1664, w_000_1665, w_000_1666, w_000_1667, w_000_1669, w_000_1671, w_000_1672, w_000_1673, w_000_1674, w_000_1675, w_000_1676, w_000_1677, w_000_1678, w_000_1679, w_000_1680, w_000_1682, w_000_1683, w_000_1684, w_000_1685, w_000_1686, w_000_1687, w_000_1688, w_000_1690, w_000_1691, w_000_1692, w_000_1693, w_000_1694, w_000_1695, w_000_1696, w_000_1698, w_000_1699, w_000_1700, w_000_1701, w_000_1702, w_000_1703, w_000_1704, w_000_1705, w_000_1706, w_000_1707, w_000_1709, w_000_1710, w_000_1711, w_000_1712, w_000_1713, w_000_1716, w_000_1717, w_000_1719, w_000_1720, w_000_1722, w_000_1723, w_000_1725, w_000_1726, w_000_1727, w_000_1728, w_000_1729, w_000_1730, w_000_1732, w_000_1733, w_000_1734, w_000_1736, w_000_1737, w_000_1739, w_000_1740, w_000_1741, w_000_1742, w_000_1744, w_000_1745, w_000_1746, w_000_1747, w_000_1748, w_000_1749, w_000_1752, w_000_1753, w_000_1754, w_000_1755, w_000_1756, w_000_1757, w_000_1758, w_000_1759, w_000_1760, w_000_1761, w_000_1762, w_000_1763, w_000_1764, w_000_1765, w_000_1766, w_000_1768, w_000_1769, w_000_1770, w_000_1771, w_000_1772, w_000_1774, w_000_1775, w_000_1776, w_000_1778, w_000_1779, w_000_1780, w_000_1781, w_000_1782, w_000_1783, w_000_1784, w_000_1785, w_000_1787, w_000_1788, w_000_1789, w_000_1790, w_000_1791, w_000_1792, w_000_1794, w_000_1795, w_000_1796, w_000_1797, w_000_1800, w_000_1801, w_000_1802, w_000_1803, w_000_1804, w_000_1805, w_000_1806, w_000_1807, w_000_1808, w_000_1809, w_000_1810, w_000_1811, w_000_1812, w_000_1813, w_000_1814, w_000_1815, w_000_1816, w_000_1817, w_000_1818, w_000_1819, w_000_1820, w_000_1821, w_000_1822, w_000_1823, w_000_1824, w_000_1826, w_000_1827, w_000_1828, w_000_1829, w_000_1830, w_000_1831, w_000_1832, w_000_1833, w_000_1834, w_000_1835, w_000_1836, w_000_1837, w_000_1838, w_000_1839, w_000_1840, w_000_1841, w_000_1842, w_000_1843, w_000_1844, w_000_1845, w_000_1846, w_000_1847, w_000_1848, w_000_1849, w_000_1850, w_000_1851, w_000_1852, w_000_1857, w_000_1859, w_000_1861, w_000_1862, w_000_1863, w_000_1864, w_000_1865, w_000_1866, w_000_1868, w_000_1869, w_000_1870, w_000_1871, w_000_1873, w_000_1875, w_000_1876, w_000_1877, w_000_1878, w_000_1879, w_000_1880, w_000_1881, w_000_1882, w_000_1883, w_000_1885, w_000_1886, w_000_1887, w_000_1888, w_000_1889, w_000_1890, w_000_1893, w_000_1894, w_000_1895, w_000_1896, w_000_1899, w_000_1900, w_000_1902, w_000_1904, w_000_1905, w_000_1906, w_000_1907, w_000_1908, w_000_1909, w_000_1910, w_000_1912, w_000_1913, w_000_1914, w_000_1916, w_000_1917, w_000_1921, w_000_1922, w_000_1923, w_000_1924, w_000_1925, w_000_1926, w_000_1929, w_000_1931, w_000_1932, w_000_1935, w_000_1939, w_000_1942, w_000_1943, w_000_1946, w_000_1947, w_000_1949, w_000_1951, w_000_1962, w_000_1969, w_000_1971, w_000_1975, w_000_1977, w_2000_000, w_2000_001, w_2000_002, w_2000_003, w_2000_004, w_2000_005, w_2000_006, w_2000_007, w_2000_008, w_2000_009, w_2000_010, w_2000_011, w_2000_012, w_2000_013, w_2000_014, w_2000_015, w_2000_016, w_2000_017, w_2000_018, w_2000_019, w_2000_020, w_2000_021, w_2000_022, w_2000_023, w_2000_024, w_2000_025, w_2000_026, w_2000_027, w_2000_028, w_2000_029, w_2000_030, w_2000_031, w_2000_032, w_2000_033, w_2000_034, w_2000_035, w_2000_036, w_2000_037, w_2000_038, w_2000_039, w_2000_040, w_2000_041, w_2000_042, w_2000_043, w_2000_044, w_2000_045, w_2000_046, w_2000_047, w_2000_048, w_2000_049, w_2000_050, w_2000_051, w_2000_052, w_2000_053, w_2000_054, w_2000_055, w_2000_056, w_2000_057, w_2000_058, w_2000_059, w_2000_060, w_2000_061, w_2000_062, w_2000_063, w_2000_064, w_2000_065, w_2000_066, w_2000_067, w_2000_068, w_2000_069, w_2000_070, w_2000_071, w_2000_072, w_2000_073, w_2000_074, w_2000_075, w_2000_076, w_2000_077, w_2000_078, w_2000_079, w_2000_080, w_2000_081, w_2000_082, w_2000_083, w_2000_084, w_2000_085, w_2000_086, w_2000_087, w_2000_088, w_2000_089, w_2000_090, w_2000_091, w_2000_092, w_2000_093, w_2000_094, w_2000_095, w_2000_096, w_2000_097, w_2000_098, w_2000_099, w_2000_100, w_2000_101, w_2000_102, w_2000_103, w_2000_104, w_2000_105, w_2000_106, w_2000_107, w_2000_108, w_2000_109, w_2000_110 ;
  combLogic I0(  w_000_000, w_000_001, w_000_002, w_000_003, w_000_004, w_000_005, w_000_006, w_000_007, w_000_008, w_000_009, w_000_010, w_000_011, w_000_012, w_000_013, w_000_014, w_000_015, w_000_016, w_000_017, w_000_018, w_000_019, w_000_020, w_000_021, w_000_022, w_000_023, w_000_024, w_000_025, w_000_026, w_000_027, w_000_028, w_000_029, w_000_030, w_000_031, w_000_032, w_000_033, w_000_034, w_000_035, w_000_036, w_000_037, w_000_038, w_000_039, w_000_040, w_000_041, w_000_042, w_000_043, w_000_044, w_000_045, w_000_046, w_000_047, w_000_048, w_000_049, w_000_050, w_000_051, w_000_052, w_000_053, w_000_054, w_000_055, w_000_056, w_000_057, w_000_058, w_000_059, w_000_060, w_000_061, w_000_062, w_000_063, w_000_065, w_000_066, w_000_067, w_000_068, w_000_069, w_000_070, w_000_071, w_000_072, w_000_073, w_000_074, w_000_075, w_000_076, w_000_077, w_000_078, w_000_079, w_000_080, w_000_081, w_000_082, w_000_083, w_000_084, w_000_085, w_000_086, w_000_087, w_000_088, w_000_089, w_000_090, w_000_091, w_000_092, w_000_093, w_000_094, w_000_095, w_000_096, w_000_097, w_000_098, w_000_099, w_000_100, w_000_101, w_000_102, w_000_103, w_000_104, w_000_105, w_000_106, w_000_107, w_000_108, w_000_109, w_000_110, w_000_111, w_000_112, w_000_113, w_000_114, w_000_115, w_000_116, w_000_117, w_000_118, w_000_119, w_000_120, w_000_121, w_000_122, w_000_123, w_000_124, w_000_125, w_000_126, w_000_127, w_000_128, w_000_129, w_000_130, w_000_131, w_000_132, w_000_133, w_000_134, w_000_135, w_000_136, w_000_137, w_000_138, w_000_139, w_000_140, w_000_141, w_000_142, w_000_143, w_000_144, w_000_145, w_000_146, w_000_147, w_000_148, w_000_149, w_000_150, w_000_151, w_000_152, w_000_153, w_000_154, w_000_155, w_000_156, w_000_157, w_000_158, w_000_159, w_000_160, w_000_161, w_000_162, w_000_163, w_000_164, w_000_165, w_000_166, w_000_167, w_000_168, w_000_169, w_000_170, w_000_171, w_000_172, w_000_173, w_000_174, w_000_175, w_000_176, w_000_177, w_000_178, w_000_179, w_000_180, w_000_181, w_000_182, w_000_183, w_000_184, w_000_185, w_000_186, w_000_187, w_000_188, w_000_189, w_000_190, w_000_191, w_000_192, w_000_193, w_000_194, w_000_195, w_000_196, w_000_197, w_000_198, w_000_199, w_000_200, w_000_201, w_000_202, w_000_203, w_000_204, w_000_205, w_000_206, w_000_207, w_000_208, w_000_209, w_000_210, w_000_211, w_000_212, w_000_213, w_000_214, w_000_215, w_000_216, w_000_217, w_000_218, w_000_219, w_000_220, w_000_221, w_000_222, w_000_223, w_000_224, w_000_225, w_000_226, w_000_227, w_000_228, w_000_229, w_000_230, w_000_231, w_000_232, w_000_233, w_000_234, w_000_235, w_000_236, w_000_237, w_000_238, w_000_239, w_000_240, w_000_241, w_000_242, w_000_243, w_000_244, w_000_245, w_000_246, w_000_247, w_000_248, w_000_249, w_000_250, w_000_251, w_000_252, w_000_253, w_000_254, w_000_255, w_000_256, w_000_257, w_000_258, w_000_259, w_000_260, w_000_261, w_000_262, w_000_263, w_000_264, w_000_265, w_000_266, w_000_267, w_000_268, w_000_269, w_000_270, w_000_271, w_000_272, w_000_273, w_000_274, w_000_275, w_000_276, w_000_277, w_000_278, w_000_279, w_000_280, w_000_281, w_000_282, w_000_283, w_000_284, w_000_285, w_000_286, w_000_287, w_000_289, w_000_290, w_000_291, w_000_292, w_000_293, w_000_294, w_000_295, w_000_296, w_000_297, w_000_298, w_000_299, w_000_300, w_000_301, w_000_302, w_000_303, w_000_304, w_000_305, w_000_306, w_000_307, w_000_308, w_000_309, w_000_310, w_000_311, w_000_312, w_000_313, w_000_314, w_000_315, w_000_316, w_000_317, w_000_318, w_000_319, w_000_320, w_000_321, w_000_322, w_000_323, w_000_324, w_000_325, w_000_326, w_000_327, w_000_328, w_000_329, w_000_330, w_000_331, w_000_332, w_000_333, w_000_334, w_000_335, w_000_336, w_000_337, w_000_338, w_000_339, w_000_340, w_000_341, w_000_342, w_000_343, w_000_344, w_000_345, w_000_346, w_000_347, w_000_348, w_000_349, w_000_350, w_000_351, w_000_352, w_000_353, w_000_354, w_000_355, w_000_356, w_000_357, w_000_358, w_000_359, w_000_360, w_000_361, w_000_362, w_000_363, w_000_364, w_000_365, w_000_366, w_000_367, w_000_368, w_000_369, w_000_370, w_000_371, w_000_372, w_000_373, w_000_374, w_000_375, w_000_376, w_000_377, w_000_378, w_000_379, w_000_380, w_000_381, w_000_382, w_000_383, w_000_384, w_000_385, w_000_386, w_000_387, w_000_388, w_000_389, w_000_390, w_000_391, w_000_392, w_000_393, w_000_394, w_000_395, w_000_396, w_000_397, w_000_398, w_000_399, w_000_400, w_000_401, w_000_402, w_000_403, w_000_404, w_000_405, w_000_406, w_000_407, w_000_408, w_000_409, w_000_410, w_000_411, w_000_412, w_000_413, w_000_414, w_000_415, w_000_416, w_000_417, w_000_418, w_000_419, w_000_420, w_000_421, w_000_422, w_000_423, w_000_424, w_000_425, w_000_426, w_000_427, w_000_428, w_000_429, w_000_430, w_000_431, w_000_432, w_000_433, w_000_434, w_000_435, w_000_436, w_000_437, w_000_438, w_000_439, w_000_440, w_000_441, w_000_442, w_000_443, w_000_444, w_000_445, w_000_446, w_000_447, w_000_448, w_000_449, w_000_450, w_000_451, w_000_452, w_000_453, w_000_454, w_000_455, w_000_456, w_000_457, w_000_458, w_000_459, w_000_460, w_000_461, w_000_462, w_000_463, w_000_464, w_000_465, w_000_466, w_000_467, w_000_468, w_000_469, w_000_470, w_000_471, w_000_472, w_000_473, w_000_474, w_000_475, w_000_476, w_000_477, w_000_478, w_000_479, w_000_480, w_000_481, w_000_482, w_000_483, w_000_484, w_000_485, w_000_486, w_000_487, w_000_488, w_000_489, w_000_490, w_000_491, w_000_492, w_000_493, w_000_494, w_000_495, w_000_496, w_000_498, w_000_499, w_000_500, w_000_501, w_000_502, w_000_503, w_000_504, w_000_505, w_000_506, w_000_507, w_000_508, w_000_509, w_000_510, w_000_511, w_000_512, w_000_513, w_000_514, w_000_515, w_000_516, w_000_517, w_000_518, w_000_519, w_000_520, w_000_521, w_000_522, w_000_523, w_000_524, w_000_525, w_000_526, w_000_527, w_000_528, w_000_529, w_000_530, w_000_531, w_000_532, w_000_533, w_000_534, w_000_535, w_000_536, w_000_537, w_000_538, w_000_539, w_000_540, w_000_541, w_000_542, w_000_543, w_000_544, w_000_545, w_000_546, w_000_547, w_000_548, w_000_549, w_000_550, w_000_551, w_000_552, w_000_553, w_000_554, w_000_555, w_000_556, w_000_557, w_000_558, w_000_559, w_000_560, w_000_561, w_000_562, w_000_563, w_000_564, w_000_565, w_000_566, w_000_567, w_000_568, w_000_569, w_000_570, w_000_571, w_000_572, w_000_573, w_000_575, w_000_576, w_000_577, w_000_578, w_000_579, w_000_580, w_000_581, w_000_582, w_000_583, w_000_584, w_000_585, w_000_586, w_000_587, w_000_588, w_000_589, w_000_590, w_000_591, w_000_592, w_000_593, w_000_594, w_000_595, w_000_596, w_000_597, w_000_598, w_000_599, w_000_600, w_000_601, w_000_602, w_000_603, w_000_604, w_000_605, w_000_606, w_000_607, w_000_608, w_000_609, w_000_610, w_000_611, w_000_612, w_000_613, w_000_614, w_000_615, w_000_616, w_000_617, w_000_618, w_000_619, w_000_620, w_000_621, w_000_622, w_000_623, w_000_624, w_000_625, w_000_626, w_000_627, w_000_628, w_000_629, w_000_630, w_000_631, w_000_632, w_000_633, w_000_634, w_000_635, w_000_636, w_000_638, w_000_639, w_000_640, w_000_641, w_000_643, w_000_644, w_000_645, w_000_646, w_000_647, w_000_648, w_000_649, w_000_650, w_000_651, w_000_652, w_000_653, w_000_654, w_000_655, w_000_656, w_000_657, w_000_658, w_000_659, w_000_660, w_000_661, w_000_662, w_000_663, w_000_664, w_000_665, w_000_667, w_000_668, w_000_669, w_000_670, w_000_671, w_000_672, w_000_673, w_000_674, w_000_675, w_000_676, w_000_677, w_000_678, w_000_679, w_000_680, w_000_681, w_000_682, w_000_683, w_000_684, w_000_685, w_000_686, w_000_687, w_000_688, w_000_689, w_000_690, w_000_691, w_000_692, w_000_693, w_000_694, w_000_695, w_000_696, w_000_697, w_000_698, w_000_699, w_000_700, w_000_701, w_000_702, w_000_703, w_000_704, w_000_705, w_000_706, w_000_707, w_000_708, w_000_709, w_000_710, w_000_711, w_000_712, w_000_713, w_000_714, w_000_715, w_000_716, w_000_717, w_000_718, w_000_719, w_000_720, w_000_721, w_000_722, w_000_723, w_000_724, w_000_725, w_000_726, w_000_727, w_000_728, w_000_729, w_000_730, w_000_731, w_000_732, w_000_733, w_000_734, w_000_735, w_000_736, w_000_737, w_000_738, w_000_739, w_000_740, w_000_741, w_000_742, w_000_743, w_000_744, w_000_745, w_000_746, w_000_747, w_000_748, w_000_749, w_000_750, w_000_751, w_000_752, w_000_753, w_000_754, w_000_755, w_000_756, w_000_757, w_000_758, w_000_759, w_000_760, w_000_761, w_000_762, w_000_763, w_000_764, w_000_765, w_000_766, w_000_767, w_000_768, w_000_769, w_000_770, w_000_771, w_000_772, w_000_773, w_000_774, w_000_775, w_000_776, w_000_777, w_000_778, w_000_779, w_000_780, w_000_781, w_000_782, w_000_783, w_000_784, w_000_785, w_000_786, w_000_787, w_000_788, w_000_789, w_000_790, w_000_791, w_000_792, w_000_793, w_000_794, w_000_795, w_000_796, w_000_797, w_000_798, w_000_799, w_000_800, w_000_801, w_000_802, w_000_803, w_000_804, w_000_805, w_000_806, w_000_807, w_000_808, w_000_809, w_000_810, w_000_811, w_000_812, w_000_813, w_000_814, w_000_815, w_000_816, w_000_817, w_000_818, w_000_819, w_000_820, w_000_821, w_000_822, w_000_823, w_000_824, w_000_825, w_000_826, w_000_827, w_000_828, w_000_829, w_000_830, w_000_831, w_000_832, w_000_833, w_000_835, w_000_836, w_000_837, w_000_838, w_000_839, w_000_840, w_000_841, w_000_842, w_000_843, w_000_844, w_000_845, w_000_846, w_000_847, w_000_848, w_000_849, w_000_850, w_000_851, w_000_852, w_000_853, w_000_854, w_000_855, w_000_856, w_000_857, w_000_858, w_000_859, w_000_860, w_000_861, w_000_862, w_000_863, w_000_864, w_000_865, w_000_866, w_000_867, w_000_868, w_000_869, w_000_870, w_000_871, w_000_872, w_000_873, w_000_874, w_000_875, w_000_876, w_000_877, w_000_878, w_000_879, w_000_880, w_000_881, w_000_882, w_000_883, w_000_884, w_000_885, w_000_886, w_000_887, w_000_888, w_000_889, w_000_890, w_000_891, w_000_892, w_000_893, w_000_894, w_000_895, w_000_896, w_000_897, w_000_898, w_000_899, w_000_900, w_000_901, w_000_902, w_000_903, w_000_904, w_000_905, w_000_906, w_000_907, w_000_908, w_000_909, w_000_910, w_000_911, w_000_912, w_000_913, w_000_914, w_000_915, w_000_916, w_000_917, w_000_918, w_000_919, w_000_920, w_000_921, w_000_922, w_000_923, w_000_924, w_000_925, w_000_926, w_000_927, w_000_928, w_000_929, w_000_930, w_000_931, w_000_932, w_000_933, w_000_935, w_000_936, w_000_937, w_000_938, w_000_939, w_000_940, w_000_941, w_000_942, w_000_943, w_000_944, w_000_945, w_000_946, w_000_947, w_000_948, w_000_949, w_000_950, w_000_951, w_000_952, w_000_953, w_000_954, w_000_955, w_000_956, w_000_957, w_000_958, w_000_959, w_000_960, w_000_961, w_000_962, w_000_963, w_000_964, w_000_965, w_000_966, w_000_967, w_000_968, w_000_969, w_000_970, w_000_971, w_000_972, w_000_973, w_000_974, w_000_975, w_000_976, w_000_977, w_000_978, w_000_979, w_000_980, w_000_981, w_000_982, w_000_983, w_000_984, w_000_985, w_000_986, w_000_987, w_000_988, w_000_989, w_000_990, w_000_991, w_000_992, w_000_993, w_000_994, w_000_995, w_000_996, w_000_997, w_000_998, w_000_999, w_000_1000, w_000_1001, w_000_1002, w_000_1003, w_000_1004, w_000_1005, w_000_1006, w_000_1007, w_000_1008, w_000_1009, w_000_1010, w_000_1011, w_000_1012, w_000_1013, w_000_1014, w_000_1015, w_000_1016, w_000_1017, w_000_1018, w_000_1019, w_000_1020, w_000_1021, w_000_1022, w_000_1023, w_000_1024, w_000_1025, w_000_1026, w_000_1027, w_000_1028, w_000_1029, w_000_1030, w_000_1031, w_000_1032, w_000_1033, w_000_1034, w_000_1035, w_000_1036, w_000_1037, w_000_1038, w_000_1039, w_000_1040, w_000_1041, w_000_1042, w_000_1043, w_000_1044, w_000_1045, w_000_1046, w_000_1047, w_000_1048, w_000_1049, w_000_1050, w_000_1051, w_000_1052, w_000_1053, w_000_1054, w_000_1055, w_000_1056, w_000_1057, w_000_1058, w_000_1060, w_000_1061, w_000_1062, w_000_1063, w_000_1064, w_000_1065, w_000_1066, w_000_1067, w_000_1068, w_000_1069, w_000_1070, w_000_1071, w_000_1072, w_000_1073, w_000_1074, w_000_1075, w_000_1076, w_000_1077, w_000_1078, w_000_1079, w_000_1080, w_000_1081, w_000_1082, w_000_1083, w_000_1084, w_000_1085, w_000_1086, w_000_1087, w_000_1088, w_000_1089, w_000_1090, w_000_1091, w_000_1093, w_000_1094, w_000_1095, w_000_1096, w_000_1097, w_000_1098, w_000_1099, w_000_1101, w_000_1102, w_000_1103, w_000_1104, w_000_1105, w_000_1106, w_000_1107, w_000_1108, w_000_1109, w_000_1110, w_000_1111, w_000_1112, w_000_1113, w_000_1114, w_000_1115, w_000_1116, w_000_1117, w_000_1118, w_000_1119, w_000_1120, w_000_1121, w_000_1122, w_000_1123, w_000_1124, w_000_1125, w_000_1126, w_000_1127, w_000_1128, w_000_1129, w_000_1130, w_000_1131, w_000_1132, w_000_1133, w_000_1134, w_000_1136, w_000_1137, w_000_1138, w_000_1139, w_000_1140, w_000_1141, w_000_1142, w_000_1143, w_000_1144, w_000_1145, w_000_1146, w_000_1147, w_000_1148, w_000_1149, w_000_1150, w_000_1151, w_000_1152, w_000_1153, w_000_1154, w_000_1155, w_000_1156, w_000_1157, w_000_1158, w_000_1159, w_000_1160, w_000_1161, w_000_1162, w_000_1163, w_000_1165, w_000_1166, w_000_1168, w_000_1169, w_000_1171, w_000_1172, w_000_1173, w_000_1174, w_000_1175, w_000_1176, w_000_1177, w_000_1178, w_000_1179, w_000_1180, w_000_1181, w_000_1182, w_000_1183, w_000_1184, w_000_1185, w_000_1186, w_000_1187, w_000_1188, w_000_1189, w_000_1190, w_000_1191, w_000_1192, w_000_1193, w_000_1194, w_000_1195, w_000_1196, w_000_1197, w_000_1198, w_000_1199, w_000_1200, w_000_1201, w_000_1202, w_000_1203, w_000_1204, w_000_1205, w_000_1206, w_000_1207, w_000_1208, w_000_1209, w_000_1210, w_000_1211, w_000_1212, w_000_1213, w_000_1214, w_000_1215, w_000_1216, w_000_1217, w_000_1218, w_000_1219, w_000_1220, w_000_1221, w_000_1222, w_000_1223, w_000_1224, w_000_1225, w_000_1226, w_000_1227, w_000_1228, w_000_1229, w_000_1230, w_000_1231, w_000_1232, w_000_1233, w_000_1234, w_000_1235, w_000_1236, w_000_1237, w_000_1238, w_000_1239, w_000_1240, w_000_1241, w_000_1242, w_000_1243, w_000_1244, w_000_1245, w_000_1246, w_000_1247, w_000_1248, w_000_1249, w_000_1250, w_000_1251, w_000_1252, w_000_1253, w_000_1254, w_000_1255, w_000_1256, w_000_1257, w_000_1258, w_000_1259, w_000_1260, w_000_1261, w_000_1262, w_000_1264, w_000_1265, w_000_1266, w_000_1267, w_000_1268, w_000_1270, w_000_1271, w_000_1272, w_000_1274, w_000_1275, w_000_1276, w_000_1277, w_000_1278, w_000_1279, w_000_1282, w_000_1283, w_000_1284, w_000_1285, w_000_1286, w_000_1287, w_000_1288, w_000_1289, w_000_1290, w_000_1291, w_000_1293, w_000_1294, w_000_1295, w_000_1296, w_000_1297, w_000_1298, w_000_1299, w_000_1300, w_000_1301, w_000_1302, w_000_1303, w_000_1304, w_000_1305, w_000_1306, w_000_1307, w_000_1308, w_000_1309, w_000_1310, w_000_1311, w_000_1312, w_000_1313, w_000_1314, w_000_1315, w_000_1316, w_000_1317, w_000_1318, w_000_1320, w_000_1321, w_000_1322, w_000_1323, w_000_1324, w_000_1325, w_000_1326, w_000_1327, w_000_1328, w_000_1329, w_000_1330, w_000_1331, w_000_1332, w_000_1333, w_000_1334, w_000_1335, w_000_1338, w_000_1339, w_000_1340, w_000_1341, w_000_1342, w_000_1343, w_000_1344, w_000_1345, w_000_1346, w_000_1347, w_000_1348, w_000_1349, w_000_1350, w_000_1351, w_000_1352, w_000_1353, w_000_1354, w_000_1355, w_000_1356, w_000_1357, w_000_1358, w_000_1359, w_000_1360, w_000_1361, w_000_1362, w_000_1363, w_000_1365, w_000_1366, w_000_1367, w_000_1368, w_000_1369, w_000_1370, w_000_1371, w_000_1372, w_000_1373, w_000_1374, w_000_1375, w_000_1376, w_000_1377, w_000_1378, w_000_1379, w_000_1380, w_000_1381, w_000_1382, w_000_1383, w_000_1385, w_000_1386, w_000_1387, w_000_1388, w_000_1389, w_000_1390, w_000_1391, w_000_1392, w_000_1393, w_000_1394, w_000_1395, w_000_1396, w_000_1397, w_000_1398, w_000_1399, w_000_1400, w_000_1401, w_000_1402, w_000_1403, w_000_1405, w_000_1406, w_000_1407, w_000_1408, w_000_1409, w_000_1410, w_000_1411, w_000_1412, w_000_1413, w_000_1414, w_000_1415, w_000_1417, w_000_1418, w_000_1419, w_000_1421, w_000_1422, w_000_1423, w_000_1424, w_000_1425, w_000_1426, w_000_1427, w_000_1428, w_000_1429, w_000_1430, w_000_1431, w_000_1432, w_000_1433, w_000_1434, w_000_1435, w_000_1436, w_000_1437, w_000_1438, w_000_1439, w_000_1440, w_000_1441, w_000_1442, w_000_1443, w_000_1444, w_000_1445, w_000_1447, w_000_1448, w_000_1449, w_000_1450, w_000_1451, w_000_1452, w_000_1453, w_000_1454, w_000_1455, w_000_1457, w_000_1458, w_000_1459, w_000_1460, w_000_1461, w_000_1462, w_000_1463, w_000_1464, w_000_1465, w_000_1466, w_000_1467, w_000_1469, w_000_1470, w_000_1471, w_000_1472, w_000_1473, w_000_1474, w_000_1475, w_000_1476, w_000_1477, w_000_1478, w_000_1480, w_000_1481, w_000_1482, w_000_1483, w_000_1484, w_000_1485, w_000_1486, w_000_1487, w_000_1488, w_000_1489, w_000_1490, w_000_1491, w_000_1492, w_000_1493, w_000_1494, w_000_1495, w_000_1496, w_000_1497, w_000_1498, w_000_1499, w_000_1500, w_000_1501, w_000_1502, w_000_1503, w_000_1504, w_000_1505, w_000_1506, w_000_1507, w_000_1508, w_000_1509, w_000_1510, w_000_1511, w_000_1512, w_000_1513, w_000_1514, w_000_1515, w_000_1516, w_000_1518, w_000_1519, w_000_1520, w_000_1521, w_000_1522, w_000_1523, w_000_1524, w_000_1525, w_000_1526, w_000_1527, w_000_1528, w_000_1529, w_000_1530, w_000_1531, w_000_1532, w_000_1533, w_000_1534, w_000_1535, w_000_1536, w_000_1537, w_000_1538, w_000_1539, w_000_1540, w_000_1541, w_000_1542, w_000_1543, w_000_1544, w_000_1545, w_000_1546, w_000_1547, w_000_1548, w_000_1549, w_000_1550, w_000_1551, w_000_1552, w_000_1553, w_000_1554, w_000_1555, w_000_1556, w_000_1557, w_000_1558, w_000_1559, w_000_1560, w_000_1561, w_000_1562, w_000_1563, w_000_1564, w_000_1565, w_000_1566, w_000_1567, w_000_1568, w_000_1569, w_000_1570, w_000_1571, w_000_1572, w_000_1573, w_000_1574, w_000_1575, w_000_1576, w_000_1577, w_000_1578, w_000_1579, w_000_1580, w_000_1581, w_000_1583, w_000_1584, w_000_1585, w_000_1586, w_000_1587, w_000_1588, w_000_1589, w_000_1590, w_000_1591, w_000_1592, w_000_1593, w_000_1594, w_000_1595, w_000_1596, w_000_1597, w_000_1598, w_000_1599, w_000_1600, w_000_1601, w_000_1602, w_000_1603, w_000_1604, w_000_1605, w_000_1606, w_000_1607, w_000_1608, w_000_1609, w_000_1610, w_000_1611, w_000_1612, w_000_1613, w_000_1614, w_000_1615, w_000_1616, w_000_1617, w_000_1618, w_000_1619, w_000_1620, w_000_1621, w_000_1622, w_000_1623, w_000_1624, w_000_1625, w_000_1626, w_000_1627, w_000_1628, w_000_1629, w_000_1630, w_000_1631, w_000_1632, w_000_1633, w_000_1634, w_000_1635, w_000_1636, w_000_1637, w_000_1638, w_000_1639, w_000_1640, w_000_1641, w_000_1642, w_000_1643, w_000_1644, w_000_1645, w_000_1646, w_000_1647, w_000_1648, w_000_1649, w_000_1650, w_000_1651, w_000_1652, w_000_1653, w_000_1654, w_000_1655, w_000_1656, w_000_1657, w_000_1658, w_000_1659, w_000_1660, w_000_1661, w_000_1662, w_000_1663, w_000_1664, w_000_1665, w_000_1666, w_000_1667, w_000_1669, w_000_1671, w_000_1672, w_000_1673, w_000_1674, w_000_1675, w_000_1676, w_000_1677, w_000_1678, w_000_1679, w_000_1680, w_000_1682, w_000_1683, w_000_1684, w_000_1685, w_000_1686, w_000_1687, w_000_1688, w_000_1690, w_000_1691, w_000_1692, w_000_1693, w_000_1694, w_000_1695, w_000_1696, w_000_1698, w_000_1699, w_000_1700, w_000_1701, w_000_1702, w_000_1703, w_000_1704, w_000_1705, w_000_1706, w_000_1707, w_000_1709, w_000_1710, w_000_1711, w_000_1712, w_000_1713, w_000_1716, w_000_1717, w_000_1719, w_000_1720, w_000_1722, w_000_1723, w_000_1725, w_000_1726, w_000_1727, w_000_1728, w_000_1729, w_000_1730, w_000_1732, w_000_1733, w_000_1734, w_000_1736, w_000_1737, w_000_1739, w_000_1740, w_000_1741, w_000_1742, w_000_1744, w_000_1745, w_000_1746, w_000_1747, w_000_1748, w_000_1749, w_000_1752, w_000_1753, w_000_1754, w_000_1755, w_000_1756, w_000_1757, w_000_1758, w_000_1759, w_000_1760, w_000_1761, w_000_1762, w_000_1763, w_000_1764, w_000_1765, w_000_1766, w_000_1768, w_000_1769, w_000_1770, w_000_1771, w_000_1772, w_000_1774, w_000_1775, w_000_1776, w_000_1778, w_000_1779, w_000_1780, w_000_1781, w_000_1782, w_000_1783, w_000_1784, w_000_1785, w_000_1787, w_000_1788, w_000_1789, w_000_1790, w_000_1791, w_000_1792, w_000_1794, w_000_1795, w_000_1796, w_000_1797, w_000_1800, w_000_1801, w_000_1802, w_000_1803, w_000_1804, w_000_1805, w_000_1806, w_000_1807, w_000_1808, w_000_1809, w_000_1810, w_000_1811, w_000_1812, w_000_1813, w_000_1814, w_000_1815, w_000_1816, w_000_1817, w_000_1818, w_000_1819, w_000_1820, w_000_1821, w_000_1822, w_000_1823, w_000_1824, w_000_1826, w_000_1827, w_000_1828, w_000_1829, w_000_1830, w_000_1831, w_000_1832, w_000_1833, w_000_1834, w_000_1835, w_000_1836, w_000_1837, w_000_1838, w_000_1839, w_000_1840, w_000_1841, w_000_1842, w_000_1843, w_000_1844, w_000_1845, w_000_1846, w_000_1847, w_000_1848, w_000_1849, w_000_1850, w_000_1851, w_000_1852, w_000_1857, w_000_1859, w_000_1861, w_000_1862, w_000_1863, w_000_1864, w_000_1865, w_000_1866, w_000_1868, w_000_1869, w_000_1870, w_000_1871, w_000_1873, w_000_1875, w_000_1876, w_000_1877, w_000_1878, w_000_1879, w_000_1880, w_000_1881, w_000_1882, w_000_1883, w_000_1885, w_000_1886, w_000_1887, w_000_1888, w_000_1889, w_000_1890, w_000_1893, w_000_1894, w_000_1895, w_000_1896, w_000_1899, w_000_1900, w_000_1902, w_000_1904, w_000_1905, w_000_1906, w_000_1907, w_000_1908, w_000_1909, w_000_1910, w_000_1912, w_000_1913, w_000_1914, w_000_1916, w_000_1917, w_000_1921, w_000_1922, w_000_1923, w_000_1924, w_000_1925, w_000_1926, w_000_1929, w_000_1931, w_000_1932, w_000_1935, w_000_1939, w_000_1942, w_000_1943, w_000_1946, w_000_1947, w_000_1949, w_000_1951, w_000_1962, w_000_1969, w_000_1971, w_000_1975, w_000_1977, w_2000_000, w_2000_001, w_2000_002, w_2000_003, w_2000_004, w_2000_005, w_2000_006, w_2000_007, w_2000_008, w_2000_009, w_2000_010, w_2000_011, w_2000_012, w_2000_013, w_2000_014, w_2000_015, w_2000_016, w_2000_017, w_2000_018, w_2000_019, w_2000_020, w_2000_021, w_2000_022, w_2000_023, w_2000_024, w_2000_025, w_2000_026, w_2000_027, w_2000_028, w_2000_029, w_2000_030, w_2000_031, w_2000_032, w_2000_033, w_2000_034, w_2000_035, w_2000_036, w_2000_037, w_2000_038, w_2000_039, w_2000_040, w_2000_041, w_2000_042, w_2000_043, w_2000_044, w_2000_045, w_2000_046, w_2000_047, w_2000_048, w_2000_049, w_2000_050, w_2000_051, w_2000_052, w_2000_053, w_2000_054, w_2000_055, w_2000_056, w_2000_057, w_2000_058, w_2000_059, w_2000_060, w_2000_061, w_2000_062, w_2000_063, w_2000_064, w_2000_065, w_2000_066, w_2000_067, w_2000_068, w_2000_069, w_2000_070, w_2000_071, w_2000_072, w_2000_073, w_2000_074, w_2000_075, w_2000_076, w_2000_077, w_2000_078, w_2000_079, w_2000_080, w_2000_081, w_2000_082, w_2000_083, w_2000_084, w_2000_085, w_2000_086, w_2000_087, w_2000_088, w_2000_089, w_2000_090, w_2000_091, w_2000_092, w_2000_093, w_2000_094, w_2000_095, w_2000_096, w_2000_097, w_2000_098, w_2000_099, w_2000_100, w_2000_101, w_2000_102, w_2000_103, w_2000_104, w_2000_105, w_2000_106, w_2000_107, w_2000_108, w_2000_109, w_2000_110  );

  reg r0, r1, r2, r3, r4, r5, r6, r7, r8, r9, r10, r11, r12, r13, r14, r15, r16, r17, r18, r19, r20, r21, r22, r23, r24, r25, r26, r27, r28, r29, r30, r31, r32, r33, r34, r35, r36, r37, r38, r39, r40, r41, r42, r43, r44, r45, r46, r47, r48, r49, r50, r51, r52, r53, r54, r55, r56, r57, r58, r59, r60, r61, r62, r63, r64, r65, r66, r67, r68, r69, r70, r71, r72, r73, r74, r75, r76, r77, r78, r79, r80, r81, r82, r83, r84, r85, r86, r87, r88, r89, r90, r91, r92, r93, r94, r95, r96, r97, r98, r99, r100, r101, r102, r103, r104, r105, r106, r107, r108, r109, r110, r111, r112, r113, r114, r115, r116, r117, r118, r119, r120, r121, r122, r123, r124, r125, r126, r127, r128, r129, r130, r131, r132, r133, r134, r135, r136, r137, r138, r139, r140, r141, r142, r143, r144, r145, r146, r147, r148, r149, r150, r151, r152, r153, r154, r155, r156, r157, r158, r159, r160, r161, r162, r163, r164, r165, r166, r167, r168, r169, r170, r171, r172, r173, r174, r175, r176, r177, r178, r179, r180, r181, r182, r183, r184, r185, r186, r187, r188, r189, r190, r191, r192, r193, r194, r195, r196, r197, r198, r199, r200, r201, r202, r203, r204, r205, r206, r207, r208, r209, r210, r211, r212, r213, r214, r215, r216, r217, r218, r219, r220, r221, r222, r223, r224, r225, r226, r227, r228, r229, r230, r231, r232, r233, r234, r235, r236, r237, r238, r239, r240, r241, r242, r243, r244, r245, r246, r247, r248, r249, r250, r251, r252, r253, r254, r255, r256, r257, r258, r259, r260, r261, r262, r263, r264, r265, r266, r267, r268, r269, r270, r271, r272, r273, r274, r275, r276, r277, r278, r279, r280, r281, r282, r283, r284, r285, r286, r287, r288, r289, r290, r291, r292, r293, r294, r295, r296, r297, r298, r299, r300, r301, r302, r303, r304, r305, r306, r307, r308, r309, r310, r311, r312, r313, r314, r315, r316, r317, r318, r319, r320, r321, r322, r323, r324, r325, r326, r327, r328, r329, r330, r331, r332, r333, r334, r335, r336, r337, r338, r339, r340, r341, r342, r343, r344, r345, r346, r347, r348, r349, r350, r351, r352, r353, r354, r355, r356, r357, r358, r359, r360, r361, r362, r363, r364, r365, r366, r367, r368, r369, r370, r371, r372, r373, r374, r375, r376, r377, r378, r379, r380, r381, r382, r383, r384, r385, r386, r387, r388, r389, r390, r391, r392, r393, r394, r395, r396, r397, r398, r399, r400, r401, r402, r403, r404, r405, r406, r407, r408, r409, r410, r411, r412, r413, r414, r415, r416, r417, r418, r419, r420, r421, r422, r423, r424, r425, r426, r427, r428, r429, r430, r431, r432, r433, r434, r435, r436, r437, r438, r439, r440, r441, r442, r443, r444, r445, r446, r447, r448, r449, r450, r451, r452, r453, r454, r455, r456, r457, r458, r459, r460, r461, r462, r463, r464, r465, r466, r467, r468, r469, r470, r471, r472, r473, r474, r475, r476, r477, r478, r479, r480, r481, r482, r483, r484, r485, r486, r487, r488, r489, r490, r491, r492, r493, r494, r495, r496, r497, r498, r499, r500, r501, r502, r503, r504, r505, r506, r507, r508, r509, r510, r511, r512, r513, r514, r515, r516, r517, r518, r519, r520, r521, r522, r523, r524, r525, r526, r527, r528, r529, r530, r531, r532, r533, r534, r535, r536, r537, r538, r539, r540, r541, r542, r543, r544, r545, r546, r547, r548, r549, r550, r551, r552, r553, r554, r555, r556, r557, r558, r559, r560, r561, r562, r563, r564, r565, r566, r567, r568, r569, r570, r571, r572, r573, r574, r575, r576, r577, r578, r579, r580, r581, r582, r583, r584, r585, r586, r587, r588, r589, r590, r591, r592, r593, r594, r595, r596, r597, r598, r599, r600, r601, r602, r603, r604, r605, r606, r607, r608, r609, r610, r611, r612, r613, r614, r615, r616, r617, r618, r619, r620, r621, r622, r623, r624, r625, r626, r627, r628, r629, r630, r631, r632, r633, r634, r635, r636, r637, r638, r639, r640, r641, r642, r643, r644, r645, r646, r647, r648, r649, r650, r651, r652, r653, r654, r655, r656, r657, r658, r659, r660, r661, r662, r663, r664, r665, r666, r667, r668, r669, r670, r671, r672, r673, r674, r675, r676, r677, r678, r679, r680, r681, r682, r683, r684, r685, r686, r687, r688, r689, r690, r691, r692, r693, r694, r695, r696, r697, r698, r699, r700, r701, r702, r703, r704, r705, r706, r707, r708, r709, r710, r711, r712, r713, r714, r715, r716, r717, r718, r719, r720, r721, r722, r723, r724, r725, r726, r727, r728, r729, r730, r731, r732, r733, r734, r735, r736, r737, r738, r739, r740, r741, r742, r743, r744, r745, r746, r747, r748, r749, r750, r751, r752, r753, r754, r755, r756, r757, r758, r759, r760, r761, r762, r763, r764, r765, r766, r767, r768, r769, r770, r771, r772, r773, r774, r775, r776, r777, r778, r779, r780, r781, r782, r783, r784, r785, r786, r787, r788, r789, r790, r791, r792, r793, r794, r795, r796, r797, r798, r799, r800, r801, r802, r803, r804, r805, r806, r807, r808, r809, r810, r811, r812, r813, r814, r815, r816, r817, r818, r819, r820, r821, r822, r823, r824, r825, r826, r827, r828, r829, r830, r831, r832, r833, r834, r835, r836, r837, r838, r839, r840, r841, r842, r843, r844, r845, r846, r847, r848, r849, r850, r851, r852, r853, r854, r855, r856, r857, r858, r859, r860, r861, r862, r863, r864, r865, r866, r867, r868, r869, r870, r871, r872, r873, r874, r875, r876, r877, r878, r879, r880, r881, r882, r883, r884, r885, r886, r887, r888, r889, r890, r891, r892, r893, r894, r895, r896, r897, r898, r899, r900, r901, r902, r903, r904, r905, r906, r907, r908, r909, r910, r911, r912, r913, r914, r915, r916, r917, r918, r919, r920, r921, r922, r923, r924, r925, r926, r927, r928, r929, r930, r931, r932, r933, r934, r935, r936, r937, r938, r939, r940, r941, r942, r943, r944, r945, r946, r947, r948, r949, r950, r951, r952, r953, r954, r955, r956, r957, r958, r959, r960, r961, r962, r963, r964, r965, r966, r967, r968, r969, r970, r971, r972, r973, r974, r975, r976, r977, r978, r979, r980, r981, r982, r983, r984, r985, r986, r987, r988, r989, r990, r991, r992, r993, r994, r995, r996, r997, r998, r999, r1000, r1001, r1002, r1003, r1004, r1005, r1006, r1007, r1008, r1009, r1010, r1011, r1012, r1013, r1014, r1015, r1016, r1017, r1018, r1019, r1020, r1021, r1022, r1023, r1024, r1025, r1026, r1027, r1028, r1029, r1030, r1031, r1032, r1033, r1034, r1035, r1036, r1037, r1038, r1039, r1040, r1041, r1042, r1043, r1044, r1045, r1046, r1047, r1048, r1049, r1050, r1051, r1052, r1053, r1054, r1055, r1056, r1057, r1058, r1059, r1060, r1061, r1062, r1063, r1064, r1065, r1066, r1067, r1068, r1069, r1070, r1071, r1072, r1073, r1074, r1075, r1076, r1077, r1078, r1079, r1080, r1081, r1082, r1083, r1084, r1085, r1086, r1087, r1088, r1089, r1090, r1091, r1092, r1093, r1094, r1095, r1096, r1097, r1098, r1099, r1100, r1101, r1102, r1103, r1104, r1105, r1106, r1107, r1108, r1109, r1110, r1111, r1112, r1113, r1114, r1115, r1116, r1117, r1118, r1119, r1120, r1121, r1122, r1123, r1124, r1125, r1126, r1127, r1128, r1129, r1130, r1131, r1132, r1133, r1134, r1135, r1136, r1137, r1138, r1139, r1140, r1141, r1142, r1143, r1144, r1145, r1146, r1147, r1148, r1149, r1150, r1151, r1152, r1153, r1154, r1155, r1156, r1157, r1158, r1159, r1160, r1161, r1162, r1163, r1164, r1165, r1166, r1167, r1168, r1169, r1170, r1171, r1172, r1173, r1174, r1175, r1176, r1177, r1178, r1179, r1180, r1181, r1182, r1183, r1184, r1185, r1186, r1187, r1188, r1189, r1190, r1191, r1192, r1193, r1194, r1195, r1196, r1197, r1198, r1199, r1200, r1201, r1202, r1203, r1204, r1205, r1206, r1207, r1208, r1209, r1210, r1211, r1212, r1213, r1214, r1215, r1216, r1217, r1218, r1219, r1220, r1221, r1222, r1223, r1224, r1225, r1226, r1227, r1228, r1229, r1230, r1231, r1232, r1233, r1234, r1235, r1236, r1237, r1238, r1239, r1240, r1241, r1242, r1243, r1244, r1245, r1246, r1247, r1248, r1249, r1250, r1251, r1252, r1253, r1254, r1255, r1256, r1257, r1258, r1259, r1260, r1261, r1262, r1263, r1264, r1265, r1266, r1267, r1268, r1269, r1270, r1271, r1272, r1273, r1274, r1275, r1276, r1277, r1278, r1279, r1280, r1281, r1282, r1283, r1284, r1285, r1286, r1287, r1288, r1289, r1290, r1291, r1292, r1293, r1294, r1295, r1296, r1297, r1298, r1299, r1300, r1301, r1302, r1303, r1304, r1305, r1306, r1307, r1308, r1309, r1310, r1311, r1312, r1313, r1314, r1315, r1316, r1317, r1318, r1319, r1320, r1321, r1322, r1323, r1324, r1325, r1326, r1327, r1328, r1329, r1330, r1331, r1332, r1333, r1334, r1335, r1336, r1337, r1338, r1339, r1340, r1341, r1342, r1343, r1344, r1345, r1346, r1347, r1348, r1349, r1350, r1351, r1352, r1353, r1354, r1355, r1356, r1357, r1358, r1359, r1360, r1361, r1362, r1363, r1364, r1365, r1366, r1367, r1368, r1369, r1370, r1371, r1372, r1373, r1374, r1375, r1376, r1377, r1378, r1379, r1380, r1381, r1382, r1383, r1384, r1385, r1386, r1387, r1388, r1389, r1390, r1391, r1392, r1393, r1394, r1395, r1396, r1397, r1398, r1399, r1400, r1401, r1402, r1403, r1404, r1405, r1406, r1407, r1408, r1409, r1410, r1411, r1412, r1413, r1414, r1415, r1416, r1417, r1418, r1419, r1420, r1421, r1422, r1423, r1424, r1425, r1426, r1427, r1428, r1429, r1430, r1431, r1432, r1433, r1434, r1435, r1436, r1437, r1438, r1439, r1440, r1441, r1442, r1443, r1444, r1445, r1446, r1447, r1448, r1449, r1450, r1451, r1452, r1453, r1454, r1455, r1456, r1457, r1458, r1459, r1460, r1461, r1462, r1463, r1464, r1465, r1466, r1467, r1468, r1469, r1470, r1471, r1472, r1473, r1474, r1475, r1476, r1477, r1478, r1479, r1480, r1481, r1482, r1483, r1484, r1485, r1486, r1487, r1488, r1489, r1490, r1491, r1492, r1493, r1494, r1495, r1496, r1497, r1498, r1499, r1500, r1501, r1502, r1503, r1504, r1505, r1506, r1507, r1508, r1509, r1510, r1511, r1512, r1513, r1514, r1515, r1516, r1517, r1518, r1519, r1520, r1521, r1522, r1523, r1524, r1525, r1526, r1527, r1528, r1529, r1530, r1531, r1532, r1533, r1534, r1535, r1536, r1537, r1538, r1539, r1540, r1541, r1542, r1543, r1544, r1545, r1546, r1547, r1548, r1549, r1550, r1551, r1552, r1553, r1554, r1555, r1556, r1557, r1558, r1559, r1560, r1561, r1562, r1563, r1564, r1565, r1566, r1567, r1568, r1569, r1570, r1571, r1572, r1573, r1574, r1575, r1576, r1577, r1578, r1579, r1580, r1581, r1582, r1583, r1584, r1585, r1586, r1587, r1588, r1589, r1590, r1591, r1592, r1593, r1594, r1595, r1596, r1597, r1598, r1599, r1600, r1601, r1602, r1603, r1604, r1605, r1606, r1607, r1608, r1609, r1610, r1611, r1612, r1613, r1614, r1615, r1616, r1617, r1618, r1619, r1620, r1621, r1622, r1623, r1624, r1625, r1626, r1627, r1628, r1629, r1630, r1631, r1632, r1633, r1634, r1635, r1636, r1637, r1638, r1639, r1640, r1641, r1642, r1643, r1644, r1645, r1646, r1647, r1648, r1649, r1650, r1651, r1652, r1653, r1654, r1655, r1656, r1657, r1658, r1659, r1660, r1661, r1662, r1663, r1664, r1665, r1666, r1667, r1668, r1669, r1670, r1671, r1672, r1673, r1674, r1675, r1676, r1677, r1678, r1679, r1680, r1681, r1682, r1683, r1684, r1685, r1686, r1687, r1688, r1689, r1690, r1691, r1692, r1693, r1694, r1695, r1696, r1697, r1698, r1699, r1700, r1701, r1702, r1703, r1704, r1705, r1706, r1707, r1708, r1709, r1710, r1711, r1712, r1713, r1714, r1715, r1716, r1717, r1718, r1719, r1720, r1721, r1722, r1723, r1724, r1725, r1726, r1727, r1728, r1729, r1730, r1731, r1732, r1733, r1734, r1735, r1736, r1737, r1738, r1739, r1740, r1741, r1742, r1743, r1744, r1745, r1746, r1747, r1748, r1749, r1750, r1751, r1752, r1753, r1754, r1755, r1756, r1757, r1758, r1759, r1760, r1761, r1762, r1763, r1764, r1765, r1766, r1767, r1768, r1769, r1770, r1771, r1772, r1773, r1774, r1775, r1776, r1777, r1778, r1779, r1780, r1781, r1782, r1783, r1784, r1785, r1786, r1787, r1788, r1789, r1790, r1791, r1792, r1793, r1794, r1795, r1796, r1797, r1798, r1799, r1800, r1801, r1802, r1803, r1804, r1805, r1806, r1807, r1808, r1809, r1810, r1811, r1812, r1813, r1814, r1815, r1816, r1817, r1818, r1819, r1820, r1821, r1822, r1823, r1824, r1825, r1826, r1827, r1828, r1829, r1830, r1831, r1832, r1833, r1834, r1835, r1836, r1837, r1838, r1839, r1840, r1841, r1842, r1843, r1844, r1845, r1846, r1847, r1848, r1849, r1850, r1851, r1852, r1853, r1854, r1855, r1856, r1857, r1858, r1859, r1860, r1861, r1862, r1863, r1864, r1865, r1866, r1867, r1868, r1869, r1870, r1871, r1872, r1873, r1874, r1875, r1876, r1877, r1878, r1879, r1880, r1881, r1882, r1883, r1884, r1885, r1886, r1887, r1888, r1889, r1890, r1891, r1892, r1893, r1894, r1895, r1896, r1897, r1898, r1899, r1900, r1901, r1902, r1903, r1904, r1905, r1906, r1907, r1908, r1909, r1910, r1911, r1912, r1913, r1914, r1915, r1916, r1917, r1918, r1919, r1920, r1921, r1922, r1923, r1924, r1925, r1926, r1927, r1928, r1929, r1930, r1931, r1932, r1933, r1934, r1935, r1936, r1937, r1938, r1939, r1940, r1941, r1942, r1943, r1944, r1945, r1946, r1947, r1948, r1949, r1950, r1951, r1952, r1953, r1954, r1955, r1956, r1957, r1958, r1959, r1960, r1961, r1962, r1963, r1964, r1965, r1966, r1967, r1968, r1969, r1970, r1971, r1972, r1973, r1974, r1975, r1976, r1977, r1978, r1979, r1980, r1981, r1982, r1983, r1984, r1985, r1986, r1987, r1988, r1989, r1990, r1991, r1992, r1993, r1994, r1995, r1996, r1997, rEnd; 

  assign w_000_000 = r0;
  assign w_000_001 = r1;
  assign w_000_002 = r2;
  assign w_000_003 = r3;
  assign w_000_004 = r4;
  assign w_000_005 = r5;
  assign w_000_006 = r6;
  assign w_000_007 = r7;
  assign w_000_008 = r8;
  assign w_000_009 = r9;
  assign w_000_010 = r10;
  assign w_000_011 = r11;
  assign w_000_012 = r12;
  assign w_000_013 = r13;
  assign w_000_014 = r14;
  assign w_000_015 = r15;
  assign w_000_016 = r16;
  assign w_000_017 = r17;
  assign w_000_018 = r18;
  assign w_000_019 = r19;
  assign w_000_020 = r20;
  assign w_000_021 = r21;
  assign w_000_022 = r22;
  assign w_000_023 = r23;
  assign w_000_024 = r24;
  assign w_000_025 = r25;
  assign w_000_026 = r26;
  assign w_000_027 = r27;
  assign w_000_028 = r28;
  assign w_000_029 = r29;
  assign w_000_030 = r30;
  assign w_000_031 = r31;
  assign w_000_032 = r32;
  assign w_000_033 = r33;
  assign w_000_034 = r34;
  assign w_000_035 = r35;
  assign w_000_036 = r36;
  assign w_000_037 = r37;
  assign w_000_038 = r38;
  assign w_000_039 = r39;
  assign w_000_040 = r40;
  assign w_000_041 = r41;
  assign w_000_042 = r42;
  assign w_000_043 = r43;
  assign w_000_044 = r44;
  assign w_000_045 = r45;
  assign w_000_046 = r46;
  assign w_000_047 = r47;
  assign w_000_048 = r48;
  assign w_000_049 = r49;
  assign w_000_050 = r50;
  assign w_000_051 = r51;
  assign w_000_052 = r52;
  assign w_000_053 = r53;
  assign w_000_054 = r54;
  assign w_000_055 = r55;
  assign w_000_056 = r56;
  assign w_000_057 = r57;
  assign w_000_058 = r58;
  assign w_000_059 = r59;
  assign w_000_060 = r60;
  assign w_000_061 = r61;
  assign w_000_062 = r62;
  assign w_000_063 = r63;
  assign w_000_064 = r64;
  assign w_000_065 = r65;
  assign w_000_066 = r66;
  assign w_000_067 = r67;
  assign w_000_068 = r68;
  assign w_000_069 = r69;
  assign w_000_070 = r70;
  assign w_000_071 = r71;
  assign w_000_072 = r72;
  assign w_000_073 = r73;
  assign w_000_074 = r74;
  assign w_000_075 = r75;
  assign w_000_076 = r76;
  assign w_000_077 = r77;
  assign w_000_078 = r78;
  assign w_000_079 = r79;
  assign w_000_080 = r80;
  assign w_000_081 = r81;
  assign w_000_082 = r82;
  assign w_000_083 = r83;
  assign w_000_084 = r84;
  assign w_000_085 = r85;
  assign w_000_086 = r86;
  assign w_000_087 = r87;
  assign w_000_088 = r88;
  assign w_000_089 = r89;
  assign w_000_090 = r90;
  assign w_000_091 = r91;
  assign w_000_092 = r92;
  assign w_000_093 = r93;
  assign w_000_094 = r94;
  assign w_000_095 = r95;
  assign w_000_096 = r96;
  assign w_000_097 = r97;
  assign w_000_098 = r98;
  assign w_000_099 = r99;
  assign w_000_100 = r100;
  assign w_000_101 = r101;
  assign w_000_102 = r102;
  assign w_000_103 = r103;
  assign w_000_104 = r104;
  assign w_000_105 = r105;
  assign w_000_106 = r106;
  assign w_000_107 = r107;
  assign w_000_108 = r108;
  assign w_000_109 = r109;
  assign w_000_110 = r110;
  assign w_000_111 = r111;
  assign w_000_112 = r112;
  assign w_000_113 = r113;
  assign w_000_114 = r114;
  assign w_000_115 = r115;
  assign w_000_116 = r116;
  assign w_000_117 = r117;
  assign w_000_118 = r118;
  assign w_000_119 = r119;
  assign w_000_120 = r120;
  assign w_000_121 = r121;
  assign w_000_122 = r122;
  assign w_000_123 = r123;
  assign w_000_124 = r124;
  assign w_000_125 = r125;
  assign w_000_126 = r126;
  assign w_000_127 = r127;
  assign w_000_128 = r128;
  assign w_000_129 = r129;
  assign w_000_130 = r130;
  assign w_000_131 = r131;
  assign w_000_132 = r132;
  assign w_000_133 = r133;
  assign w_000_134 = r134;
  assign w_000_135 = r135;
  assign w_000_136 = r136;
  assign w_000_137 = r137;
  assign w_000_138 = r138;
  assign w_000_139 = r139;
  assign w_000_140 = r140;
  assign w_000_141 = r141;
  assign w_000_142 = r142;
  assign w_000_143 = r143;
  assign w_000_144 = r144;
  assign w_000_145 = r145;
  assign w_000_146 = r146;
  assign w_000_147 = r147;
  assign w_000_148 = r148;
  assign w_000_149 = r149;
  assign w_000_150 = r150;
  assign w_000_151 = r151;
  assign w_000_152 = r152;
  assign w_000_153 = r153;
  assign w_000_154 = r154;
  assign w_000_155 = r155;
  assign w_000_156 = r156;
  assign w_000_157 = r157;
  assign w_000_158 = r158;
  assign w_000_159 = r159;
  assign w_000_160 = r160;
  assign w_000_161 = r161;
  assign w_000_162 = r162;
  assign w_000_163 = r163;
  assign w_000_164 = r164;
  assign w_000_165 = r165;
  assign w_000_166 = r166;
  assign w_000_167 = r167;
  assign w_000_168 = r168;
  assign w_000_169 = r169;
  assign w_000_170 = r170;
  assign w_000_171 = r171;
  assign w_000_172 = r172;
  assign w_000_173 = r173;
  assign w_000_174 = r174;
  assign w_000_175 = r175;
  assign w_000_176 = r176;
  assign w_000_177 = r177;
  assign w_000_178 = r178;
  assign w_000_179 = r179;
  assign w_000_180 = r180;
  assign w_000_181 = r181;
  assign w_000_182 = r182;
  assign w_000_183 = r183;
  assign w_000_184 = r184;
  assign w_000_185 = r185;
  assign w_000_186 = r186;
  assign w_000_187 = r187;
  assign w_000_188 = r188;
  assign w_000_189 = r189;
  assign w_000_190 = r190;
  assign w_000_191 = r191;
  assign w_000_192 = r192;
  assign w_000_193 = r193;
  assign w_000_194 = r194;
  assign w_000_195 = r195;
  assign w_000_196 = r196;
  assign w_000_197 = r197;
  assign w_000_198 = r198;
  assign w_000_199 = r199;
  assign w_000_200 = r200;
  assign w_000_201 = r201;
  assign w_000_202 = r202;
  assign w_000_203 = r203;
  assign w_000_204 = r204;
  assign w_000_205 = r205;
  assign w_000_206 = r206;
  assign w_000_207 = r207;
  assign w_000_208 = r208;
  assign w_000_209 = r209;
  assign w_000_210 = r210;
  assign w_000_211 = r211;
  assign w_000_212 = r212;
  assign w_000_213 = r213;
  assign w_000_214 = r214;
  assign w_000_215 = r215;
  assign w_000_216 = r216;
  assign w_000_217 = r217;
  assign w_000_218 = r218;
  assign w_000_219 = r219;
  assign w_000_220 = r220;
  assign w_000_221 = r221;
  assign w_000_222 = r222;
  assign w_000_223 = r223;
  assign w_000_224 = r224;
  assign w_000_225 = r225;
  assign w_000_226 = r226;
  assign w_000_227 = r227;
  assign w_000_228 = r228;
  assign w_000_229 = r229;
  assign w_000_230 = r230;
  assign w_000_231 = r231;
  assign w_000_232 = r232;
  assign w_000_233 = r233;
  assign w_000_234 = r234;
  assign w_000_235 = r235;
  assign w_000_236 = r236;
  assign w_000_237 = r237;
  assign w_000_238 = r238;
  assign w_000_239 = r239;
  assign w_000_240 = r240;
  assign w_000_241 = r241;
  assign w_000_242 = r242;
  assign w_000_243 = r243;
  assign w_000_244 = r244;
  assign w_000_245 = r245;
  assign w_000_246 = r246;
  assign w_000_247 = r247;
  assign w_000_248 = r248;
  assign w_000_249 = r249;
  assign w_000_250 = r250;
  assign w_000_251 = r251;
  assign w_000_252 = r252;
  assign w_000_253 = r253;
  assign w_000_254 = r254;
  assign w_000_255 = r255;
  assign w_000_256 = r256;
  assign w_000_257 = r257;
  assign w_000_258 = r258;
  assign w_000_259 = r259;
  assign w_000_260 = r260;
  assign w_000_261 = r261;
  assign w_000_262 = r262;
  assign w_000_263 = r263;
  assign w_000_264 = r264;
  assign w_000_265 = r265;
  assign w_000_266 = r266;
  assign w_000_267 = r267;
  assign w_000_268 = r268;
  assign w_000_269 = r269;
  assign w_000_270 = r270;
  assign w_000_271 = r271;
  assign w_000_272 = r272;
  assign w_000_273 = r273;
  assign w_000_274 = r274;
  assign w_000_275 = r275;
  assign w_000_276 = r276;
  assign w_000_277 = r277;
  assign w_000_278 = r278;
  assign w_000_279 = r279;
  assign w_000_280 = r280;
  assign w_000_281 = r281;
  assign w_000_282 = r282;
  assign w_000_283 = r283;
  assign w_000_284 = r284;
  assign w_000_285 = r285;
  assign w_000_286 = r286;
  assign w_000_287 = r287;
  assign w_000_288 = r288;
  assign w_000_289 = r289;
  assign w_000_290 = r290;
  assign w_000_291 = r291;
  assign w_000_292 = r292;
  assign w_000_293 = r293;
  assign w_000_294 = r294;
  assign w_000_295 = r295;
  assign w_000_296 = r296;
  assign w_000_297 = r297;
  assign w_000_298 = r298;
  assign w_000_299 = r299;
  assign w_000_300 = r300;
  assign w_000_301 = r301;
  assign w_000_302 = r302;
  assign w_000_303 = r303;
  assign w_000_304 = r304;
  assign w_000_305 = r305;
  assign w_000_306 = r306;
  assign w_000_307 = r307;
  assign w_000_308 = r308;
  assign w_000_309 = r309;
  assign w_000_310 = r310;
  assign w_000_311 = r311;
  assign w_000_312 = r312;
  assign w_000_313 = r313;
  assign w_000_314 = r314;
  assign w_000_315 = r315;
  assign w_000_316 = r316;
  assign w_000_317 = r317;
  assign w_000_318 = r318;
  assign w_000_319 = r319;
  assign w_000_320 = r320;
  assign w_000_321 = r321;
  assign w_000_322 = r322;
  assign w_000_323 = r323;
  assign w_000_324 = r324;
  assign w_000_325 = r325;
  assign w_000_326 = r326;
  assign w_000_327 = r327;
  assign w_000_328 = r328;
  assign w_000_329 = r329;
  assign w_000_330 = r330;
  assign w_000_331 = r331;
  assign w_000_332 = r332;
  assign w_000_333 = r333;
  assign w_000_334 = r334;
  assign w_000_335 = r335;
  assign w_000_336 = r336;
  assign w_000_337 = r337;
  assign w_000_338 = r338;
  assign w_000_339 = r339;
  assign w_000_340 = r340;
  assign w_000_341 = r341;
  assign w_000_342 = r342;
  assign w_000_343 = r343;
  assign w_000_344 = r344;
  assign w_000_345 = r345;
  assign w_000_346 = r346;
  assign w_000_347 = r347;
  assign w_000_348 = r348;
  assign w_000_349 = r349;
  assign w_000_350 = r350;
  assign w_000_351 = r351;
  assign w_000_352 = r352;
  assign w_000_353 = r353;
  assign w_000_354 = r354;
  assign w_000_355 = r355;
  assign w_000_356 = r356;
  assign w_000_357 = r357;
  assign w_000_358 = r358;
  assign w_000_359 = r359;
  assign w_000_360 = r360;
  assign w_000_361 = r361;
  assign w_000_362 = r362;
  assign w_000_363 = r363;
  assign w_000_364 = r364;
  assign w_000_365 = r365;
  assign w_000_366 = r366;
  assign w_000_367 = r367;
  assign w_000_368 = r368;
  assign w_000_369 = r369;
  assign w_000_370 = r370;
  assign w_000_371 = r371;
  assign w_000_372 = r372;
  assign w_000_373 = r373;
  assign w_000_374 = r374;
  assign w_000_375 = r375;
  assign w_000_376 = r376;
  assign w_000_377 = r377;
  assign w_000_378 = r378;
  assign w_000_379 = r379;
  assign w_000_380 = r380;
  assign w_000_381 = r381;
  assign w_000_382 = r382;
  assign w_000_383 = r383;
  assign w_000_384 = r384;
  assign w_000_385 = r385;
  assign w_000_386 = r386;
  assign w_000_387 = r387;
  assign w_000_388 = r388;
  assign w_000_389 = r389;
  assign w_000_390 = r390;
  assign w_000_391 = r391;
  assign w_000_392 = r392;
  assign w_000_393 = r393;
  assign w_000_394 = r394;
  assign w_000_395 = r395;
  assign w_000_396 = r396;
  assign w_000_397 = r397;
  assign w_000_398 = r398;
  assign w_000_399 = r399;
  assign w_000_400 = r400;
  assign w_000_401 = r401;
  assign w_000_402 = r402;
  assign w_000_403 = r403;
  assign w_000_404 = r404;
  assign w_000_405 = r405;
  assign w_000_406 = r406;
  assign w_000_407 = r407;
  assign w_000_408 = r408;
  assign w_000_409 = r409;
  assign w_000_410 = r410;
  assign w_000_411 = r411;
  assign w_000_412 = r412;
  assign w_000_413 = r413;
  assign w_000_414 = r414;
  assign w_000_415 = r415;
  assign w_000_416 = r416;
  assign w_000_417 = r417;
  assign w_000_418 = r418;
  assign w_000_419 = r419;
  assign w_000_420 = r420;
  assign w_000_421 = r421;
  assign w_000_422 = r422;
  assign w_000_423 = r423;
  assign w_000_424 = r424;
  assign w_000_425 = r425;
  assign w_000_426 = r426;
  assign w_000_427 = r427;
  assign w_000_428 = r428;
  assign w_000_429 = r429;
  assign w_000_430 = r430;
  assign w_000_431 = r431;
  assign w_000_432 = r432;
  assign w_000_433 = r433;
  assign w_000_434 = r434;
  assign w_000_435 = r435;
  assign w_000_436 = r436;
  assign w_000_437 = r437;
  assign w_000_438 = r438;
  assign w_000_439 = r439;
  assign w_000_440 = r440;
  assign w_000_441 = r441;
  assign w_000_442 = r442;
  assign w_000_443 = r443;
  assign w_000_444 = r444;
  assign w_000_445 = r445;
  assign w_000_446 = r446;
  assign w_000_447 = r447;
  assign w_000_448 = r448;
  assign w_000_449 = r449;
  assign w_000_450 = r450;
  assign w_000_451 = r451;
  assign w_000_452 = r452;
  assign w_000_453 = r453;
  assign w_000_454 = r454;
  assign w_000_455 = r455;
  assign w_000_456 = r456;
  assign w_000_457 = r457;
  assign w_000_458 = r458;
  assign w_000_459 = r459;
  assign w_000_460 = r460;
  assign w_000_461 = r461;
  assign w_000_462 = r462;
  assign w_000_463 = r463;
  assign w_000_464 = r464;
  assign w_000_465 = r465;
  assign w_000_466 = r466;
  assign w_000_467 = r467;
  assign w_000_468 = r468;
  assign w_000_469 = r469;
  assign w_000_470 = r470;
  assign w_000_471 = r471;
  assign w_000_472 = r472;
  assign w_000_473 = r473;
  assign w_000_474 = r474;
  assign w_000_475 = r475;
  assign w_000_476 = r476;
  assign w_000_477 = r477;
  assign w_000_478 = r478;
  assign w_000_479 = r479;
  assign w_000_480 = r480;
  assign w_000_481 = r481;
  assign w_000_482 = r482;
  assign w_000_483 = r483;
  assign w_000_484 = r484;
  assign w_000_485 = r485;
  assign w_000_486 = r486;
  assign w_000_487 = r487;
  assign w_000_488 = r488;
  assign w_000_489 = r489;
  assign w_000_490 = r490;
  assign w_000_491 = r491;
  assign w_000_492 = r492;
  assign w_000_493 = r493;
  assign w_000_494 = r494;
  assign w_000_495 = r495;
  assign w_000_496 = r496;
  assign w_000_497 = r497;
  assign w_000_498 = r498;
  assign w_000_499 = r499;
  assign w_000_500 = r500;
  assign w_000_501 = r501;
  assign w_000_502 = r502;
  assign w_000_503 = r503;
  assign w_000_504 = r504;
  assign w_000_505 = r505;
  assign w_000_506 = r506;
  assign w_000_507 = r507;
  assign w_000_508 = r508;
  assign w_000_509 = r509;
  assign w_000_510 = r510;
  assign w_000_511 = r511;
  assign w_000_512 = r512;
  assign w_000_513 = r513;
  assign w_000_514 = r514;
  assign w_000_515 = r515;
  assign w_000_516 = r516;
  assign w_000_517 = r517;
  assign w_000_518 = r518;
  assign w_000_519 = r519;
  assign w_000_520 = r520;
  assign w_000_521 = r521;
  assign w_000_522 = r522;
  assign w_000_523 = r523;
  assign w_000_524 = r524;
  assign w_000_525 = r525;
  assign w_000_526 = r526;
  assign w_000_527 = r527;
  assign w_000_528 = r528;
  assign w_000_529 = r529;
  assign w_000_530 = r530;
  assign w_000_531 = r531;
  assign w_000_532 = r532;
  assign w_000_533 = r533;
  assign w_000_534 = r534;
  assign w_000_535 = r535;
  assign w_000_536 = r536;
  assign w_000_537 = r537;
  assign w_000_538 = r538;
  assign w_000_539 = r539;
  assign w_000_540 = r540;
  assign w_000_541 = r541;
  assign w_000_542 = r542;
  assign w_000_543 = r543;
  assign w_000_544 = r544;
  assign w_000_545 = r545;
  assign w_000_546 = r546;
  assign w_000_547 = r547;
  assign w_000_548 = r548;
  assign w_000_549 = r549;
  assign w_000_550 = r550;
  assign w_000_551 = r551;
  assign w_000_552 = r552;
  assign w_000_553 = r553;
  assign w_000_554 = r554;
  assign w_000_555 = r555;
  assign w_000_556 = r556;
  assign w_000_557 = r557;
  assign w_000_558 = r558;
  assign w_000_559 = r559;
  assign w_000_560 = r560;
  assign w_000_561 = r561;
  assign w_000_562 = r562;
  assign w_000_563 = r563;
  assign w_000_564 = r564;
  assign w_000_565 = r565;
  assign w_000_566 = r566;
  assign w_000_567 = r567;
  assign w_000_568 = r568;
  assign w_000_569 = r569;
  assign w_000_570 = r570;
  assign w_000_571 = r571;
  assign w_000_572 = r572;
  assign w_000_573 = r573;
  assign w_000_574 = r574;
  assign w_000_575 = r575;
  assign w_000_576 = r576;
  assign w_000_577 = r577;
  assign w_000_578 = r578;
  assign w_000_579 = r579;
  assign w_000_580 = r580;
  assign w_000_581 = r581;
  assign w_000_582 = r582;
  assign w_000_583 = r583;
  assign w_000_584 = r584;
  assign w_000_585 = r585;
  assign w_000_586 = r586;
  assign w_000_587 = r587;
  assign w_000_588 = r588;
  assign w_000_589 = r589;
  assign w_000_590 = r590;
  assign w_000_591 = r591;
  assign w_000_592 = r592;
  assign w_000_593 = r593;
  assign w_000_594 = r594;
  assign w_000_595 = r595;
  assign w_000_596 = r596;
  assign w_000_597 = r597;
  assign w_000_598 = r598;
  assign w_000_599 = r599;
  assign w_000_600 = r600;
  assign w_000_601 = r601;
  assign w_000_602 = r602;
  assign w_000_603 = r603;
  assign w_000_604 = r604;
  assign w_000_605 = r605;
  assign w_000_606 = r606;
  assign w_000_607 = r607;
  assign w_000_608 = r608;
  assign w_000_609 = r609;
  assign w_000_610 = r610;
  assign w_000_611 = r611;
  assign w_000_612 = r612;
  assign w_000_613 = r613;
  assign w_000_614 = r614;
  assign w_000_615 = r615;
  assign w_000_616 = r616;
  assign w_000_617 = r617;
  assign w_000_618 = r618;
  assign w_000_619 = r619;
  assign w_000_620 = r620;
  assign w_000_621 = r621;
  assign w_000_622 = r622;
  assign w_000_623 = r623;
  assign w_000_624 = r624;
  assign w_000_625 = r625;
  assign w_000_626 = r626;
  assign w_000_627 = r627;
  assign w_000_628 = r628;
  assign w_000_629 = r629;
  assign w_000_630 = r630;
  assign w_000_631 = r631;
  assign w_000_632 = r632;
  assign w_000_633 = r633;
  assign w_000_634 = r634;
  assign w_000_635 = r635;
  assign w_000_636 = r636;
  assign w_000_637 = r637;
  assign w_000_638 = r638;
  assign w_000_639 = r639;
  assign w_000_640 = r640;
  assign w_000_641 = r641;
  assign w_000_642 = r642;
  assign w_000_643 = r643;
  assign w_000_644 = r644;
  assign w_000_645 = r645;
  assign w_000_646 = r646;
  assign w_000_647 = r647;
  assign w_000_648 = r648;
  assign w_000_649 = r649;
  assign w_000_650 = r650;
  assign w_000_651 = r651;
  assign w_000_652 = r652;
  assign w_000_653 = r653;
  assign w_000_654 = r654;
  assign w_000_655 = r655;
  assign w_000_656 = r656;
  assign w_000_657 = r657;
  assign w_000_658 = r658;
  assign w_000_659 = r659;
  assign w_000_660 = r660;
  assign w_000_661 = r661;
  assign w_000_662 = r662;
  assign w_000_663 = r663;
  assign w_000_664 = r664;
  assign w_000_665 = r665;
  assign w_000_666 = r666;
  assign w_000_667 = r667;
  assign w_000_668 = r668;
  assign w_000_669 = r669;
  assign w_000_670 = r670;
  assign w_000_671 = r671;
  assign w_000_672 = r672;
  assign w_000_673 = r673;
  assign w_000_674 = r674;
  assign w_000_675 = r675;
  assign w_000_676 = r676;
  assign w_000_677 = r677;
  assign w_000_678 = r678;
  assign w_000_679 = r679;
  assign w_000_680 = r680;
  assign w_000_681 = r681;
  assign w_000_682 = r682;
  assign w_000_683 = r683;
  assign w_000_684 = r684;
  assign w_000_685 = r685;
  assign w_000_686 = r686;
  assign w_000_687 = r687;
  assign w_000_688 = r688;
  assign w_000_689 = r689;
  assign w_000_690 = r690;
  assign w_000_691 = r691;
  assign w_000_692 = r692;
  assign w_000_693 = r693;
  assign w_000_694 = r694;
  assign w_000_695 = r695;
  assign w_000_696 = r696;
  assign w_000_697 = r697;
  assign w_000_698 = r698;
  assign w_000_699 = r699;
  assign w_000_700 = r700;
  assign w_000_701 = r701;
  assign w_000_702 = r702;
  assign w_000_703 = r703;
  assign w_000_704 = r704;
  assign w_000_705 = r705;
  assign w_000_706 = r706;
  assign w_000_707 = r707;
  assign w_000_708 = r708;
  assign w_000_709 = r709;
  assign w_000_710 = r710;
  assign w_000_711 = r711;
  assign w_000_712 = r712;
  assign w_000_713 = r713;
  assign w_000_714 = r714;
  assign w_000_715 = r715;
  assign w_000_716 = r716;
  assign w_000_717 = r717;
  assign w_000_718 = r718;
  assign w_000_719 = r719;
  assign w_000_720 = r720;
  assign w_000_721 = r721;
  assign w_000_722 = r722;
  assign w_000_723 = r723;
  assign w_000_724 = r724;
  assign w_000_725 = r725;
  assign w_000_726 = r726;
  assign w_000_727 = r727;
  assign w_000_728 = r728;
  assign w_000_729 = r729;
  assign w_000_730 = r730;
  assign w_000_731 = r731;
  assign w_000_732 = r732;
  assign w_000_733 = r733;
  assign w_000_734 = r734;
  assign w_000_735 = r735;
  assign w_000_736 = r736;
  assign w_000_737 = r737;
  assign w_000_738 = r738;
  assign w_000_739 = r739;
  assign w_000_740 = r740;
  assign w_000_741 = r741;
  assign w_000_742 = r742;
  assign w_000_743 = r743;
  assign w_000_744 = r744;
  assign w_000_745 = r745;
  assign w_000_746 = r746;
  assign w_000_747 = r747;
  assign w_000_748 = r748;
  assign w_000_749 = r749;
  assign w_000_750 = r750;
  assign w_000_751 = r751;
  assign w_000_752 = r752;
  assign w_000_753 = r753;
  assign w_000_754 = r754;
  assign w_000_755 = r755;
  assign w_000_756 = r756;
  assign w_000_757 = r757;
  assign w_000_758 = r758;
  assign w_000_759 = r759;
  assign w_000_760 = r760;
  assign w_000_761 = r761;
  assign w_000_762 = r762;
  assign w_000_763 = r763;
  assign w_000_764 = r764;
  assign w_000_765 = r765;
  assign w_000_766 = r766;
  assign w_000_767 = r767;
  assign w_000_768 = r768;
  assign w_000_769 = r769;
  assign w_000_770 = r770;
  assign w_000_771 = r771;
  assign w_000_772 = r772;
  assign w_000_773 = r773;
  assign w_000_774 = r774;
  assign w_000_775 = r775;
  assign w_000_776 = r776;
  assign w_000_777 = r777;
  assign w_000_778 = r778;
  assign w_000_779 = r779;
  assign w_000_780 = r780;
  assign w_000_781 = r781;
  assign w_000_782 = r782;
  assign w_000_783 = r783;
  assign w_000_784 = r784;
  assign w_000_785 = r785;
  assign w_000_786 = r786;
  assign w_000_787 = r787;
  assign w_000_788 = r788;
  assign w_000_789 = r789;
  assign w_000_790 = r790;
  assign w_000_791 = r791;
  assign w_000_792 = r792;
  assign w_000_793 = r793;
  assign w_000_794 = r794;
  assign w_000_795 = r795;
  assign w_000_796 = r796;
  assign w_000_797 = r797;
  assign w_000_798 = r798;
  assign w_000_799 = r799;
  assign w_000_800 = r800;
  assign w_000_801 = r801;
  assign w_000_802 = r802;
  assign w_000_803 = r803;
  assign w_000_804 = r804;
  assign w_000_805 = r805;
  assign w_000_806 = r806;
  assign w_000_807 = r807;
  assign w_000_808 = r808;
  assign w_000_809 = r809;
  assign w_000_810 = r810;
  assign w_000_811 = r811;
  assign w_000_812 = r812;
  assign w_000_813 = r813;
  assign w_000_814 = r814;
  assign w_000_815 = r815;
  assign w_000_816 = r816;
  assign w_000_817 = r817;
  assign w_000_818 = r818;
  assign w_000_819 = r819;
  assign w_000_820 = r820;
  assign w_000_821 = r821;
  assign w_000_822 = r822;
  assign w_000_823 = r823;
  assign w_000_824 = r824;
  assign w_000_825 = r825;
  assign w_000_826 = r826;
  assign w_000_827 = r827;
  assign w_000_828 = r828;
  assign w_000_829 = r829;
  assign w_000_830 = r830;
  assign w_000_831 = r831;
  assign w_000_832 = r832;
  assign w_000_833 = r833;
  assign w_000_834 = r834;
  assign w_000_835 = r835;
  assign w_000_836 = r836;
  assign w_000_837 = r837;
  assign w_000_838 = r838;
  assign w_000_839 = r839;
  assign w_000_840 = r840;
  assign w_000_841 = r841;
  assign w_000_842 = r842;
  assign w_000_843 = r843;
  assign w_000_844 = r844;
  assign w_000_845 = r845;
  assign w_000_846 = r846;
  assign w_000_847 = r847;
  assign w_000_848 = r848;
  assign w_000_849 = r849;
  assign w_000_850 = r850;
  assign w_000_851 = r851;
  assign w_000_852 = r852;
  assign w_000_853 = r853;
  assign w_000_854 = r854;
  assign w_000_855 = r855;
  assign w_000_856 = r856;
  assign w_000_857 = r857;
  assign w_000_858 = r858;
  assign w_000_859 = r859;
  assign w_000_860 = r860;
  assign w_000_861 = r861;
  assign w_000_862 = r862;
  assign w_000_863 = r863;
  assign w_000_864 = r864;
  assign w_000_865 = r865;
  assign w_000_866 = r866;
  assign w_000_867 = r867;
  assign w_000_868 = r868;
  assign w_000_869 = r869;
  assign w_000_870 = r870;
  assign w_000_871 = r871;
  assign w_000_872 = r872;
  assign w_000_873 = r873;
  assign w_000_874 = r874;
  assign w_000_875 = r875;
  assign w_000_876 = r876;
  assign w_000_877 = r877;
  assign w_000_878 = r878;
  assign w_000_879 = r879;
  assign w_000_880 = r880;
  assign w_000_881 = r881;
  assign w_000_882 = r882;
  assign w_000_883 = r883;
  assign w_000_884 = r884;
  assign w_000_885 = r885;
  assign w_000_886 = r886;
  assign w_000_887 = r887;
  assign w_000_888 = r888;
  assign w_000_889 = r889;
  assign w_000_890 = r890;
  assign w_000_891 = r891;
  assign w_000_892 = r892;
  assign w_000_893 = r893;
  assign w_000_894 = r894;
  assign w_000_895 = r895;
  assign w_000_896 = r896;
  assign w_000_897 = r897;
  assign w_000_898 = r898;
  assign w_000_899 = r899;
  assign w_000_900 = r900;
  assign w_000_901 = r901;
  assign w_000_902 = r902;
  assign w_000_903 = r903;
  assign w_000_904 = r904;
  assign w_000_905 = r905;
  assign w_000_906 = r906;
  assign w_000_907 = r907;
  assign w_000_908 = r908;
  assign w_000_909 = r909;
  assign w_000_910 = r910;
  assign w_000_911 = r911;
  assign w_000_912 = r912;
  assign w_000_913 = r913;
  assign w_000_914 = r914;
  assign w_000_915 = r915;
  assign w_000_916 = r916;
  assign w_000_917 = r917;
  assign w_000_918 = r918;
  assign w_000_919 = r919;
  assign w_000_920 = r920;
  assign w_000_921 = r921;
  assign w_000_922 = r922;
  assign w_000_923 = r923;
  assign w_000_924 = r924;
  assign w_000_925 = r925;
  assign w_000_926 = r926;
  assign w_000_927 = r927;
  assign w_000_928 = r928;
  assign w_000_929 = r929;
  assign w_000_930 = r930;
  assign w_000_931 = r931;
  assign w_000_932 = r932;
  assign w_000_933 = r933;
  assign w_000_934 = r934;
  assign w_000_935 = r935;
  assign w_000_936 = r936;
  assign w_000_937 = r937;
  assign w_000_938 = r938;
  assign w_000_939 = r939;
  assign w_000_940 = r940;
  assign w_000_941 = r941;
  assign w_000_942 = r942;
  assign w_000_943 = r943;
  assign w_000_944 = r944;
  assign w_000_945 = r945;
  assign w_000_946 = r946;
  assign w_000_947 = r947;
  assign w_000_948 = r948;
  assign w_000_949 = r949;
  assign w_000_950 = r950;
  assign w_000_951 = r951;
  assign w_000_952 = r952;
  assign w_000_953 = r953;
  assign w_000_954 = r954;
  assign w_000_955 = r955;
  assign w_000_956 = r956;
  assign w_000_957 = r957;
  assign w_000_958 = r958;
  assign w_000_959 = r959;
  assign w_000_960 = r960;
  assign w_000_961 = r961;
  assign w_000_962 = r962;
  assign w_000_963 = r963;
  assign w_000_964 = r964;
  assign w_000_965 = r965;
  assign w_000_966 = r966;
  assign w_000_967 = r967;
  assign w_000_968 = r968;
  assign w_000_969 = r969;
  assign w_000_970 = r970;
  assign w_000_971 = r971;
  assign w_000_972 = r972;
  assign w_000_973 = r973;
  assign w_000_974 = r974;
  assign w_000_975 = r975;
  assign w_000_976 = r976;
  assign w_000_977 = r977;
  assign w_000_978 = r978;
  assign w_000_979 = r979;
  assign w_000_980 = r980;
  assign w_000_981 = r981;
  assign w_000_982 = r982;
  assign w_000_983 = r983;
  assign w_000_984 = r984;
  assign w_000_985 = r985;
  assign w_000_986 = r986;
  assign w_000_987 = r987;
  assign w_000_988 = r988;
  assign w_000_989 = r989;
  assign w_000_990 = r990;
  assign w_000_991 = r991;
  assign w_000_992 = r992;
  assign w_000_993 = r993;
  assign w_000_994 = r994;
  assign w_000_995 = r995;
  assign w_000_996 = r996;
  assign w_000_997 = r997;
  assign w_000_998 = r998;
  assign w_000_999 = r999;
  assign w_000_1000 = r1000;
  assign w_000_1001 = r1001;
  assign w_000_1002 = r1002;
  assign w_000_1003 = r1003;
  assign w_000_1004 = r1004;
  assign w_000_1005 = r1005;
  assign w_000_1006 = r1006;
  assign w_000_1007 = r1007;
  assign w_000_1008 = r1008;
  assign w_000_1009 = r1009;
  assign w_000_1010 = r1010;
  assign w_000_1011 = r1011;
  assign w_000_1012 = r1012;
  assign w_000_1013 = r1013;
  assign w_000_1014 = r1014;
  assign w_000_1015 = r1015;
  assign w_000_1016 = r1016;
  assign w_000_1017 = r1017;
  assign w_000_1018 = r1018;
  assign w_000_1019 = r1019;
  assign w_000_1020 = r1020;
  assign w_000_1021 = r1021;
  assign w_000_1022 = r1022;
  assign w_000_1023 = r1023;
  assign w_000_1024 = r1024;
  assign w_000_1025 = r1025;
  assign w_000_1026 = r1026;
  assign w_000_1027 = r1027;
  assign w_000_1028 = r1028;
  assign w_000_1029 = r1029;
  assign w_000_1030 = r1030;
  assign w_000_1031 = r1031;
  assign w_000_1032 = r1032;
  assign w_000_1033 = r1033;
  assign w_000_1034 = r1034;
  assign w_000_1035 = r1035;
  assign w_000_1036 = r1036;
  assign w_000_1037 = r1037;
  assign w_000_1038 = r1038;
  assign w_000_1039 = r1039;
  assign w_000_1040 = r1040;
  assign w_000_1041 = r1041;
  assign w_000_1042 = r1042;
  assign w_000_1043 = r1043;
  assign w_000_1044 = r1044;
  assign w_000_1045 = r1045;
  assign w_000_1046 = r1046;
  assign w_000_1047 = r1047;
  assign w_000_1048 = r1048;
  assign w_000_1049 = r1049;
  assign w_000_1050 = r1050;
  assign w_000_1051 = r1051;
  assign w_000_1052 = r1052;
  assign w_000_1053 = r1053;
  assign w_000_1054 = r1054;
  assign w_000_1055 = r1055;
  assign w_000_1056 = r1056;
  assign w_000_1057 = r1057;
  assign w_000_1058 = r1058;
  assign w_000_1059 = r1059;
  assign w_000_1060 = r1060;
  assign w_000_1061 = r1061;
  assign w_000_1062 = r1062;
  assign w_000_1063 = r1063;
  assign w_000_1064 = r1064;
  assign w_000_1065 = r1065;
  assign w_000_1066 = r1066;
  assign w_000_1067 = r1067;
  assign w_000_1068 = r1068;
  assign w_000_1069 = r1069;
  assign w_000_1070 = r1070;
  assign w_000_1071 = r1071;
  assign w_000_1072 = r1072;
  assign w_000_1073 = r1073;
  assign w_000_1074 = r1074;
  assign w_000_1075 = r1075;
  assign w_000_1076 = r1076;
  assign w_000_1077 = r1077;
  assign w_000_1078 = r1078;
  assign w_000_1079 = r1079;
  assign w_000_1080 = r1080;
  assign w_000_1081 = r1081;
  assign w_000_1082 = r1082;
  assign w_000_1083 = r1083;
  assign w_000_1084 = r1084;
  assign w_000_1085 = r1085;
  assign w_000_1086 = r1086;
  assign w_000_1087 = r1087;
  assign w_000_1088 = r1088;
  assign w_000_1089 = r1089;
  assign w_000_1090 = r1090;
  assign w_000_1091 = r1091;
  assign w_000_1092 = r1092;
  assign w_000_1093 = r1093;
  assign w_000_1094 = r1094;
  assign w_000_1095 = r1095;
  assign w_000_1096 = r1096;
  assign w_000_1097 = r1097;
  assign w_000_1098 = r1098;
  assign w_000_1099 = r1099;
  assign w_000_1100 = r1100;
  assign w_000_1101 = r1101;
  assign w_000_1102 = r1102;
  assign w_000_1103 = r1103;
  assign w_000_1104 = r1104;
  assign w_000_1105 = r1105;
  assign w_000_1106 = r1106;
  assign w_000_1107 = r1107;
  assign w_000_1108 = r1108;
  assign w_000_1109 = r1109;
  assign w_000_1110 = r1110;
  assign w_000_1111 = r1111;
  assign w_000_1112 = r1112;
  assign w_000_1113 = r1113;
  assign w_000_1114 = r1114;
  assign w_000_1115 = r1115;
  assign w_000_1116 = r1116;
  assign w_000_1117 = r1117;
  assign w_000_1118 = r1118;
  assign w_000_1119 = r1119;
  assign w_000_1120 = r1120;
  assign w_000_1121 = r1121;
  assign w_000_1122 = r1122;
  assign w_000_1123 = r1123;
  assign w_000_1124 = r1124;
  assign w_000_1125 = r1125;
  assign w_000_1126 = r1126;
  assign w_000_1127 = r1127;
  assign w_000_1128 = r1128;
  assign w_000_1129 = r1129;
  assign w_000_1130 = r1130;
  assign w_000_1131 = r1131;
  assign w_000_1132 = r1132;
  assign w_000_1133 = r1133;
  assign w_000_1134 = r1134;
  assign w_000_1135 = r1135;
  assign w_000_1136 = r1136;
  assign w_000_1137 = r1137;
  assign w_000_1138 = r1138;
  assign w_000_1139 = r1139;
  assign w_000_1140 = r1140;
  assign w_000_1141 = r1141;
  assign w_000_1142 = r1142;
  assign w_000_1143 = r1143;
  assign w_000_1144 = r1144;
  assign w_000_1145 = r1145;
  assign w_000_1146 = r1146;
  assign w_000_1147 = r1147;
  assign w_000_1148 = r1148;
  assign w_000_1149 = r1149;
  assign w_000_1150 = r1150;
  assign w_000_1151 = r1151;
  assign w_000_1152 = r1152;
  assign w_000_1153 = r1153;
  assign w_000_1154 = r1154;
  assign w_000_1155 = r1155;
  assign w_000_1156 = r1156;
  assign w_000_1157 = r1157;
  assign w_000_1158 = r1158;
  assign w_000_1159 = r1159;
  assign w_000_1160 = r1160;
  assign w_000_1161 = r1161;
  assign w_000_1162 = r1162;
  assign w_000_1163 = r1163;
  assign w_000_1164 = r1164;
  assign w_000_1165 = r1165;
  assign w_000_1166 = r1166;
  assign w_000_1167 = r1167;
  assign w_000_1168 = r1168;
  assign w_000_1169 = r1169;
  assign w_000_1170 = r1170;
  assign w_000_1171 = r1171;
  assign w_000_1172 = r1172;
  assign w_000_1173 = r1173;
  assign w_000_1174 = r1174;
  assign w_000_1175 = r1175;
  assign w_000_1176 = r1176;
  assign w_000_1177 = r1177;
  assign w_000_1178 = r1178;
  assign w_000_1179 = r1179;
  assign w_000_1180 = r1180;
  assign w_000_1181 = r1181;
  assign w_000_1182 = r1182;
  assign w_000_1183 = r1183;
  assign w_000_1184 = r1184;
  assign w_000_1185 = r1185;
  assign w_000_1186 = r1186;
  assign w_000_1187 = r1187;
  assign w_000_1188 = r1188;
  assign w_000_1189 = r1189;
  assign w_000_1190 = r1190;
  assign w_000_1191 = r1191;
  assign w_000_1192 = r1192;
  assign w_000_1193 = r1193;
  assign w_000_1194 = r1194;
  assign w_000_1195 = r1195;
  assign w_000_1196 = r1196;
  assign w_000_1197 = r1197;
  assign w_000_1198 = r1198;
  assign w_000_1199 = r1199;
  assign w_000_1200 = r1200;
  assign w_000_1201 = r1201;
  assign w_000_1202 = r1202;
  assign w_000_1203 = r1203;
  assign w_000_1204 = r1204;
  assign w_000_1205 = r1205;
  assign w_000_1206 = r1206;
  assign w_000_1207 = r1207;
  assign w_000_1208 = r1208;
  assign w_000_1209 = r1209;
  assign w_000_1210 = r1210;
  assign w_000_1211 = r1211;
  assign w_000_1212 = r1212;
  assign w_000_1213 = r1213;
  assign w_000_1214 = r1214;
  assign w_000_1215 = r1215;
  assign w_000_1216 = r1216;
  assign w_000_1217 = r1217;
  assign w_000_1218 = r1218;
  assign w_000_1219 = r1219;
  assign w_000_1220 = r1220;
  assign w_000_1221 = r1221;
  assign w_000_1222 = r1222;
  assign w_000_1223 = r1223;
  assign w_000_1224 = r1224;
  assign w_000_1225 = r1225;
  assign w_000_1226 = r1226;
  assign w_000_1227 = r1227;
  assign w_000_1228 = r1228;
  assign w_000_1229 = r1229;
  assign w_000_1230 = r1230;
  assign w_000_1231 = r1231;
  assign w_000_1232 = r1232;
  assign w_000_1233 = r1233;
  assign w_000_1234 = r1234;
  assign w_000_1235 = r1235;
  assign w_000_1236 = r1236;
  assign w_000_1237 = r1237;
  assign w_000_1238 = r1238;
  assign w_000_1239 = r1239;
  assign w_000_1240 = r1240;
  assign w_000_1241 = r1241;
  assign w_000_1242 = r1242;
  assign w_000_1243 = r1243;
  assign w_000_1244 = r1244;
  assign w_000_1245 = r1245;
  assign w_000_1246 = r1246;
  assign w_000_1247 = r1247;
  assign w_000_1248 = r1248;
  assign w_000_1249 = r1249;
  assign w_000_1250 = r1250;
  assign w_000_1251 = r1251;
  assign w_000_1252 = r1252;
  assign w_000_1253 = r1253;
  assign w_000_1254 = r1254;
  assign w_000_1255 = r1255;
  assign w_000_1256 = r1256;
  assign w_000_1257 = r1257;
  assign w_000_1258 = r1258;
  assign w_000_1259 = r1259;
  assign w_000_1260 = r1260;
  assign w_000_1261 = r1261;
  assign w_000_1262 = r1262;
  assign w_000_1263 = r1263;
  assign w_000_1264 = r1264;
  assign w_000_1265 = r1265;
  assign w_000_1266 = r1266;
  assign w_000_1267 = r1267;
  assign w_000_1268 = r1268;
  assign w_000_1269 = r1269;
  assign w_000_1270 = r1270;
  assign w_000_1271 = r1271;
  assign w_000_1272 = r1272;
  assign w_000_1273 = r1273;
  assign w_000_1274 = r1274;
  assign w_000_1275 = r1275;
  assign w_000_1276 = r1276;
  assign w_000_1277 = r1277;
  assign w_000_1278 = r1278;
  assign w_000_1279 = r1279;
  assign w_000_1280 = r1280;
  assign w_000_1281 = r1281;
  assign w_000_1282 = r1282;
  assign w_000_1283 = r1283;
  assign w_000_1284 = r1284;
  assign w_000_1285 = r1285;
  assign w_000_1286 = r1286;
  assign w_000_1287 = r1287;
  assign w_000_1288 = r1288;
  assign w_000_1289 = r1289;
  assign w_000_1290 = r1290;
  assign w_000_1291 = r1291;
  assign w_000_1292 = r1292;
  assign w_000_1293 = r1293;
  assign w_000_1294 = r1294;
  assign w_000_1295 = r1295;
  assign w_000_1296 = r1296;
  assign w_000_1297 = r1297;
  assign w_000_1298 = r1298;
  assign w_000_1299 = r1299;
  assign w_000_1300 = r1300;
  assign w_000_1301 = r1301;
  assign w_000_1302 = r1302;
  assign w_000_1303 = r1303;
  assign w_000_1304 = r1304;
  assign w_000_1305 = r1305;
  assign w_000_1306 = r1306;
  assign w_000_1307 = r1307;
  assign w_000_1308 = r1308;
  assign w_000_1309 = r1309;
  assign w_000_1310 = r1310;
  assign w_000_1311 = r1311;
  assign w_000_1312 = r1312;
  assign w_000_1313 = r1313;
  assign w_000_1314 = r1314;
  assign w_000_1315 = r1315;
  assign w_000_1316 = r1316;
  assign w_000_1317 = r1317;
  assign w_000_1318 = r1318;
  assign w_000_1319 = r1319;
  assign w_000_1320 = r1320;
  assign w_000_1321 = r1321;
  assign w_000_1322 = r1322;
  assign w_000_1323 = r1323;
  assign w_000_1324 = r1324;
  assign w_000_1325 = r1325;
  assign w_000_1326 = r1326;
  assign w_000_1327 = r1327;
  assign w_000_1328 = r1328;
  assign w_000_1329 = r1329;
  assign w_000_1330 = r1330;
  assign w_000_1331 = r1331;
  assign w_000_1332 = r1332;
  assign w_000_1333 = r1333;
  assign w_000_1334 = r1334;
  assign w_000_1335 = r1335;
  assign w_000_1336 = r1336;
  assign w_000_1337 = r1337;
  assign w_000_1338 = r1338;
  assign w_000_1339 = r1339;
  assign w_000_1340 = r1340;
  assign w_000_1341 = r1341;
  assign w_000_1342 = r1342;
  assign w_000_1343 = r1343;
  assign w_000_1344 = r1344;
  assign w_000_1345 = r1345;
  assign w_000_1346 = r1346;
  assign w_000_1347 = r1347;
  assign w_000_1348 = r1348;
  assign w_000_1349 = r1349;
  assign w_000_1350 = r1350;
  assign w_000_1351 = r1351;
  assign w_000_1352 = r1352;
  assign w_000_1353 = r1353;
  assign w_000_1354 = r1354;
  assign w_000_1355 = r1355;
  assign w_000_1356 = r1356;
  assign w_000_1357 = r1357;
  assign w_000_1358 = r1358;
  assign w_000_1359 = r1359;
  assign w_000_1360 = r1360;
  assign w_000_1361 = r1361;
  assign w_000_1362 = r1362;
  assign w_000_1363 = r1363;
  assign w_000_1364 = r1364;
  assign w_000_1365 = r1365;
  assign w_000_1366 = r1366;
  assign w_000_1367 = r1367;
  assign w_000_1368 = r1368;
  assign w_000_1369 = r1369;
  assign w_000_1370 = r1370;
  assign w_000_1371 = r1371;
  assign w_000_1372 = r1372;
  assign w_000_1373 = r1373;
  assign w_000_1374 = r1374;
  assign w_000_1375 = r1375;
  assign w_000_1376 = r1376;
  assign w_000_1377 = r1377;
  assign w_000_1378 = r1378;
  assign w_000_1379 = r1379;
  assign w_000_1380 = r1380;
  assign w_000_1381 = r1381;
  assign w_000_1382 = r1382;
  assign w_000_1383 = r1383;
  assign w_000_1384 = r1384;
  assign w_000_1385 = r1385;
  assign w_000_1386 = r1386;
  assign w_000_1387 = r1387;
  assign w_000_1388 = r1388;
  assign w_000_1389 = r1389;
  assign w_000_1390 = r1390;
  assign w_000_1391 = r1391;
  assign w_000_1392 = r1392;
  assign w_000_1393 = r1393;
  assign w_000_1394 = r1394;
  assign w_000_1395 = r1395;
  assign w_000_1396 = r1396;
  assign w_000_1397 = r1397;
  assign w_000_1398 = r1398;
  assign w_000_1399 = r1399;
  assign w_000_1400 = r1400;
  assign w_000_1401 = r1401;
  assign w_000_1402 = r1402;
  assign w_000_1403 = r1403;
  assign w_000_1404 = r1404;
  assign w_000_1405 = r1405;
  assign w_000_1406 = r1406;
  assign w_000_1407 = r1407;
  assign w_000_1408 = r1408;
  assign w_000_1409 = r1409;
  assign w_000_1410 = r1410;
  assign w_000_1411 = r1411;
  assign w_000_1412 = r1412;
  assign w_000_1413 = r1413;
  assign w_000_1414 = r1414;
  assign w_000_1415 = r1415;
  assign w_000_1416 = r1416;
  assign w_000_1417 = r1417;
  assign w_000_1418 = r1418;
  assign w_000_1419 = r1419;
  assign w_000_1420 = r1420;
  assign w_000_1421 = r1421;
  assign w_000_1422 = r1422;
  assign w_000_1423 = r1423;
  assign w_000_1424 = r1424;
  assign w_000_1425 = r1425;
  assign w_000_1426 = r1426;
  assign w_000_1427 = r1427;
  assign w_000_1428 = r1428;
  assign w_000_1429 = r1429;
  assign w_000_1430 = r1430;
  assign w_000_1431 = r1431;
  assign w_000_1432 = r1432;
  assign w_000_1433 = r1433;
  assign w_000_1434 = r1434;
  assign w_000_1435 = r1435;
  assign w_000_1436 = r1436;
  assign w_000_1437 = r1437;
  assign w_000_1438 = r1438;
  assign w_000_1439 = r1439;
  assign w_000_1440 = r1440;
  assign w_000_1441 = r1441;
  assign w_000_1442 = r1442;
  assign w_000_1443 = r1443;
  assign w_000_1444 = r1444;
  assign w_000_1445 = r1445;
  assign w_000_1446 = r1446;
  assign w_000_1447 = r1447;
  assign w_000_1448 = r1448;
  assign w_000_1449 = r1449;
  assign w_000_1450 = r1450;
  assign w_000_1451 = r1451;
  assign w_000_1452 = r1452;
  assign w_000_1453 = r1453;
  assign w_000_1454 = r1454;
  assign w_000_1455 = r1455;
  assign w_000_1456 = r1456;
  assign w_000_1457 = r1457;
  assign w_000_1458 = r1458;
  assign w_000_1459 = r1459;
  assign w_000_1460 = r1460;
  assign w_000_1461 = r1461;
  assign w_000_1462 = r1462;
  assign w_000_1463 = r1463;
  assign w_000_1464 = r1464;
  assign w_000_1465 = r1465;
  assign w_000_1466 = r1466;
  assign w_000_1467 = r1467;
  assign w_000_1468 = r1468;
  assign w_000_1469 = r1469;
  assign w_000_1470 = r1470;
  assign w_000_1471 = r1471;
  assign w_000_1472 = r1472;
  assign w_000_1473 = r1473;
  assign w_000_1474 = r1474;
  assign w_000_1475 = r1475;
  assign w_000_1476 = r1476;
  assign w_000_1477 = r1477;
  assign w_000_1478 = r1478;
  assign w_000_1479 = r1479;
  assign w_000_1480 = r1480;
  assign w_000_1481 = r1481;
  assign w_000_1482 = r1482;
  assign w_000_1483 = r1483;
  assign w_000_1484 = r1484;
  assign w_000_1485 = r1485;
  assign w_000_1486 = r1486;
  assign w_000_1487 = r1487;
  assign w_000_1488 = r1488;
  assign w_000_1489 = r1489;
  assign w_000_1490 = r1490;
  assign w_000_1491 = r1491;
  assign w_000_1492 = r1492;
  assign w_000_1493 = r1493;
  assign w_000_1494 = r1494;
  assign w_000_1495 = r1495;
  assign w_000_1496 = r1496;
  assign w_000_1497 = r1497;
  assign w_000_1498 = r1498;
  assign w_000_1499 = r1499;
  assign w_000_1500 = r1500;
  assign w_000_1501 = r1501;
  assign w_000_1502 = r1502;
  assign w_000_1503 = r1503;
  assign w_000_1504 = r1504;
  assign w_000_1505 = r1505;
  assign w_000_1506 = r1506;
  assign w_000_1507 = r1507;
  assign w_000_1508 = r1508;
  assign w_000_1509 = r1509;
  assign w_000_1510 = r1510;
  assign w_000_1511 = r1511;
  assign w_000_1512 = r1512;
  assign w_000_1513 = r1513;
  assign w_000_1514 = r1514;
  assign w_000_1515 = r1515;
  assign w_000_1516 = r1516;
  assign w_000_1517 = r1517;
  assign w_000_1518 = r1518;
  assign w_000_1519 = r1519;
  assign w_000_1520 = r1520;
  assign w_000_1521 = r1521;
  assign w_000_1522 = r1522;
  assign w_000_1523 = r1523;
  assign w_000_1524 = r1524;
  assign w_000_1525 = r1525;
  assign w_000_1526 = r1526;
  assign w_000_1527 = r1527;
  assign w_000_1528 = r1528;
  assign w_000_1529 = r1529;
  assign w_000_1530 = r1530;
  assign w_000_1531 = r1531;
  assign w_000_1532 = r1532;
  assign w_000_1533 = r1533;
  assign w_000_1534 = r1534;
  assign w_000_1535 = r1535;
  assign w_000_1536 = r1536;
  assign w_000_1537 = r1537;
  assign w_000_1538 = r1538;
  assign w_000_1539 = r1539;
  assign w_000_1540 = r1540;
  assign w_000_1541 = r1541;
  assign w_000_1542 = r1542;
  assign w_000_1543 = r1543;
  assign w_000_1544 = r1544;
  assign w_000_1545 = r1545;
  assign w_000_1546 = r1546;
  assign w_000_1547 = r1547;
  assign w_000_1548 = r1548;
  assign w_000_1549 = r1549;
  assign w_000_1550 = r1550;
  assign w_000_1551 = r1551;
  assign w_000_1552 = r1552;
  assign w_000_1553 = r1553;
  assign w_000_1554 = r1554;
  assign w_000_1555 = r1555;
  assign w_000_1556 = r1556;
  assign w_000_1557 = r1557;
  assign w_000_1558 = r1558;
  assign w_000_1559 = r1559;
  assign w_000_1560 = r1560;
  assign w_000_1561 = r1561;
  assign w_000_1562 = r1562;
  assign w_000_1563 = r1563;
  assign w_000_1564 = r1564;
  assign w_000_1565 = r1565;
  assign w_000_1566 = r1566;
  assign w_000_1567 = r1567;
  assign w_000_1568 = r1568;
  assign w_000_1569 = r1569;
  assign w_000_1570 = r1570;
  assign w_000_1571 = r1571;
  assign w_000_1572 = r1572;
  assign w_000_1573 = r1573;
  assign w_000_1574 = r1574;
  assign w_000_1575 = r1575;
  assign w_000_1576 = r1576;
  assign w_000_1577 = r1577;
  assign w_000_1578 = r1578;
  assign w_000_1579 = r1579;
  assign w_000_1580 = r1580;
  assign w_000_1581 = r1581;
  assign w_000_1582 = r1582;
  assign w_000_1583 = r1583;
  assign w_000_1584 = r1584;
  assign w_000_1585 = r1585;
  assign w_000_1586 = r1586;
  assign w_000_1587 = r1587;
  assign w_000_1588 = r1588;
  assign w_000_1589 = r1589;
  assign w_000_1590 = r1590;
  assign w_000_1591 = r1591;
  assign w_000_1592 = r1592;
  assign w_000_1593 = r1593;
  assign w_000_1594 = r1594;
  assign w_000_1595 = r1595;
  assign w_000_1596 = r1596;
  assign w_000_1597 = r1597;
  assign w_000_1598 = r1598;
  assign w_000_1599 = r1599;
  assign w_000_1600 = r1600;
  assign w_000_1601 = r1601;
  assign w_000_1602 = r1602;
  assign w_000_1603 = r1603;
  assign w_000_1604 = r1604;
  assign w_000_1605 = r1605;
  assign w_000_1606 = r1606;
  assign w_000_1607 = r1607;
  assign w_000_1608 = r1608;
  assign w_000_1609 = r1609;
  assign w_000_1610 = r1610;
  assign w_000_1611 = r1611;
  assign w_000_1612 = r1612;
  assign w_000_1613 = r1613;
  assign w_000_1614 = r1614;
  assign w_000_1615 = r1615;
  assign w_000_1616 = r1616;
  assign w_000_1617 = r1617;
  assign w_000_1618 = r1618;
  assign w_000_1619 = r1619;
  assign w_000_1620 = r1620;
  assign w_000_1621 = r1621;
  assign w_000_1622 = r1622;
  assign w_000_1623 = r1623;
  assign w_000_1624 = r1624;
  assign w_000_1625 = r1625;
  assign w_000_1626 = r1626;
  assign w_000_1627 = r1627;
  assign w_000_1628 = r1628;
  assign w_000_1629 = r1629;
  assign w_000_1630 = r1630;
  assign w_000_1631 = r1631;
  assign w_000_1632 = r1632;
  assign w_000_1633 = r1633;
  assign w_000_1634 = r1634;
  assign w_000_1635 = r1635;
  assign w_000_1636 = r1636;
  assign w_000_1637 = r1637;
  assign w_000_1638 = r1638;
  assign w_000_1639 = r1639;
  assign w_000_1640 = r1640;
  assign w_000_1641 = r1641;
  assign w_000_1642 = r1642;
  assign w_000_1643 = r1643;
  assign w_000_1644 = r1644;
  assign w_000_1645 = r1645;
  assign w_000_1646 = r1646;
  assign w_000_1647 = r1647;
  assign w_000_1648 = r1648;
  assign w_000_1649 = r1649;
  assign w_000_1650 = r1650;
  assign w_000_1651 = r1651;
  assign w_000_1652 = r1652;
  assign w_000_1653 = r1653;
  assign w_000_1654 = r1654;
  assign w_000_1655 = r1655;
  assign w_000_1656 = r1656;
  assign w_000_1657 = r1657;
  assign w_000_1658 = r1658;
  assign w_000_1659 = r1659;
  assign w_000_1660 = r1660;
  assign w_000_1661 = r1661;
  assign w_000_1662 = r1662;
  assign w_000_1663 = r1663;
  assign w_000_1664 = r1664;
  assign w_000_1665 = r1665;
  assign w_000_1666 = r1666;
  assign w_000_1667 = r1667;
  assign w_000_1668 = r1668;
  assign w_000_1669 = r1669;
  assign w_000_1670 = r1670;
  assign w_000_1671 = r1671;
  assign w_000_1672 = r1672;
  assign w_000_1673 = r1673;
  assign w_000_1674 = r1674;
  assign w_000_1675 = r1675;
  assign w_000_1676 = r1676;
  assign w_000_1677 = r1677;
  assign w_000_1678 = r1678;
  assign w_000_1679 = r1679;
  assign w_000_1680 = r1680;
  assign w_000_1681 = r1681;
  assign w_000_1682 = r1682;
  assign w_000_1683 = r1683;
  assign w_000_1684 = r1684;
  assign w_000_1685 = r1685;
  assign w_000_1686 = r1686;
  assign w_000_1687 = r1687;
  assign w_000_1688 = r1688;
  assign w_000_1689 = r1689;
  assign w_000_1690 = r1690;
  assign w_000_1691 = r1691;
  assign w_000_1692 = r1692;
  assign w_000_1693 = r1693;
  assign w_000_1694 = r1694;
  assign w_000_1695 = r1695;
  assign w_000_1696 = r1696;
  assign w_000_1697 = r1697;
  assign w_000_1698 = r1698;
  assign w_000_1699 = r1699;
  assign w_000_1700 = r1700;
  assign w_000_1701 = r1701;
  assign w_000_1702 = r1702;
  assign w_000_1703 = r1703;
  assign w_000_1704 = r1704;
  assign w_000_1705 = r1705;
  assign w_000_1706 = r1706;
  assign w_000_1707 = r1707;
  assign w_000_1708 = r1708;
  assign w_000_1709 = r1709;
  assign w_000_1710 = r1710;
  assign w_000_1711 = r1711;
  assign w_000_1712 = r1712;
  assign w_000_1713 = r1713;
  assign w_000_1714 = r1714;
  assign w_000_1715 = r1715;
  assign w_000_1716 = r1716;
  assign w_000_1717 = r1717;
  assign w_000_1718 = r1718;
  assign w_000_1719 = r1719;
  assign w_000_1720 = r1720;
  assign w_000_1721 = r1721;
  assign w_000_1722 = r1722;
  assign w_000_1723 = r1723;
  assign w_000_1724 = r1724;
  assign w_000_1725 = r1725;
  assign w_000_1726 = r1726;
  assign w_000_1727 = r1727;
  assign w_000_1728 = r1728;
  assign w_000_1729 = r1729;
  assign w_000_1730 = r1730;
  assign w_000_1731 = r1731;
  assign w_000_1732 = r1732;
  assign w_000_1733 = r1733;
  assign w_000_1734 = r1734;
  assign w_000_1735 = r1735;
  assign w_000_1736 = r1736;
  assign w_000_1737 = r1737;
  assign w_000_1738 = r1738;
  assign w_000_1739 = r1739;
  assign w_000_1740 = r1740;
  assign w_000_1741 = r1741;
  assign w_000_1742 = r1742;
  assign w_000_1743 = r1743;
  assign w_000_1744 = r1744;
  assign w_000_1745 = r1745;
  assign w_000_1746 = r1746;
  assign w_000_1747 = r1747;
  assign w_000_1748 = r1748;
  assign w_000_1749 = r1749;
  assign w_000_1750 = r1750;
  assign w_000_1751 = r1751;
  assign w_000_1752 = r1752;
  assign w_000_1753 = r1753;
  assign w_000_1754 = r1754;
  assign w_000_1755 = r1755;
  assign w_000_1756 = r1756;
  assign w_000_1757 = r1757;
  assign w_000_1758 = r1758;
  assign w_000_1759 = r1759;
  assign w_000_1760 = r1760;
  assign w_000_1761 = r1761;
  assign w_000_1762 = r1762;
  assign w_000_1763 = r1763;
  assign w_000_1764 = r1764;
  assign w_000_1765 = r1765;
  assign w_000_1766 = r1766;
  assign w_000_1767 = r1767;
  assign w_000_1768 = r1768;
  assign w_000_1769 = r1769;
  assign w_000_1770 = r1770;
  assign w_000_1771 = r1771;
  assign w_000_1772 = r1772;
  assign w_000_1773 = r1773;
  assign w_000_1774 = r1774;
  assign w_000_1775 = r1775;
  assign w_000_1776 = r1776;
  assign w_000_1777 = r1777;
  assign w_000_1778 = r1778;
  assign w_000_1779 = r1779;
  assign w_000_1780 = r1780;
  assign w_000_1781 = r1781;
  assign w_000_1782 = r1782;
  assign w_000_1783 = r1783;
  assign w_000_1784 = r1784;
  assign w_000_1785 = r1785;
  assign w_000_1786 = r1786;
  assign w_000_1787 = r1787;
  assign w_000_1788 = r1788;
  assign w_000_1789 = r1789;
  assign w_000_1790 = r1790;
  assign w_000_1791 = r1791;
  assign w_000_1792 = r1792;
  assign w_000_1793 = r1793;
  assign w_000_1794 = r1794;
  assign w_000_1795 = r1795;
  assign w_000_1796 = r1796;
  assign w_000_1797 = r1797;
  assign w_000_1798 = r1798;
  assign w_000_1799 = r1799;
  assign w_000_1800 = r1800;
  assign w_000_1801 = r1801;
  assign w_000_1802 = r1802;
  assign w_000_1803 = r1803;
  assign w_000_1804 = r1804;
  assign w_000_1805 = r1805;
  assign w_000_1806 = r1806;
  assign w_000_1807 = r1807;
  assign w_000_1808 = r1808;
  assign w_000_1809 = r1809;
  assign w_000_1810 = r1810;
  assign w_000_1811 = r1811;
  assign w_000_1812 = r1812;
  assign w_000_1813 = r1813;
  assign w_000_1814 = r1814;
  assign w_000_1815 = r1815;
  assign w_000_1816 = r1816;
  assign w_000_1817 = r1817;
  assign w_000_1818 = r1818;
  assign w_000_1819 = r1819;
  assign w_000_1820 = r1820;
  assign w_000_1821 = r1821;
  assign w_000_1822 = r1822;
  assign w_000_1823 = r1823;
  assign w_000_1824 = r1824;
  assign w_000_1825 = r1825;
  assign w_000_1826 = r1826;
  assign w_000_1827 = r1827;
  assign w_000_1828 = r1828;
  assign w_000_1829 = r1829;
  assign w_000_1830 = r1830;
  assign w_000_1831 = r1831;
  assign w_000_1832 = r1832;
  assign w_000_1833 = r1833;
  assign w_000_1834 = r1834;
  assign w_000_1835 = r1835;
  assign w_000_1836 = r1836;
  assign w_000_1837 = r1837;
  assign w_000_1838 = r1838;
  assign w_000_1839 = r1839;
  assign w_000_1840 = r1840;
  assign w_000_1841 = r1841;
  assign w_000_1842 = r1842;
  assign w_000_1843 = r1843;
  assign w_000_1844 = r1844;
  assign w_000_1845 = r1845;
  assign w_000_1846 = r1846;
  assign w_000_1847 = r1847;
  assign w_000_1848 = r1848;
  assign w_000_1849 = r1849;
  assign w_000_1850 = r1850;
  assign w_000_1851 = r1851;
  assign w_000_1852 = r1852;
  assign w_000_1853 = r1853;
  assign w_000_1854 = r1854;
  assign w_000_1855 = r1855;
  assign w_000_1856 = r1856;
  assign w_000_1857 = r1857;
  assign w_000_1858 = r1858;
  assign w_000_1859 = r1859;
  assign w_000_1860 = r1860;
  assign w_000_1861 = r1861;
  assign w_000_1862 = r1862;
  assign w_000_1863 = r1863;
  assign w_000_1864 = r1864;
  assign w_000_1865 = r1865;
  assign w_000_1866 = r1866;
  assign w_000_1867 = r1867;
  assign w_000_1868 = r1868;
  assign w_000_1869 = r1869;
  assign w_000_1870 = r1870;
  assign w_000_1871 = r1871;
  assign w_000_1872 = r1872;
  assign w_000_1873 = r1873;
  assign w_000_1874 = r1874;
  assign w_000_1875 = r1875;
  assign w_000_1876 = r1876;
  assign w_000_1877 = r1877;
  assign w_000_1878 = r1878;
  assign w_000_1879 = r1879;
  assign w_000_1880 = r1880;
  assign w_000_1881 = r1881;
  assign w_000_1882 = r1882;
  assign w_000_1883 = r1883;
  assign w_000_1884 = r1884;
  assign w_000_1885 = r1885;
  assign w_000_1886 = r1886;
  assign w_000_1887 = r1887;
  assign w_000_1888 = r1888;
  assign w_000_1889 = r1889;
  assign w_000_1890 = r1890;
  assign w_000_1891 = r1891;
  assign w_000_1892 = r1892;
  assign w_000_1893 = r1893;
  assign w_000_1894 = r1894;
  assign w_000_1895 = r1895;
  assign w_000_1896 = r1896;
  assign w_000_1897 = r1897;
  assign w_000_1898 = r1898;
  assign w_000_1899 = r1899;
  assign w_000_1900 = r1900;
  assign w_000_1901 = r1901;
  assign w_000_1902 = r1902;
  assign w_000_1903 = r1903;
  assign w_000_1904 = r1904;
  assign w_000_1905 = r1905;
  assign w_000_1906 = r1906;
  assign w_000_1907 = r1907;
  assign w_000_1908 = r1908;
  assign w_000_1909 = r1909;
  assign w_000_1910 = r1910;
  assign w_000_1911 = r1911;
  assign w_000_1912 = r1912;
  assign w_000_1913 = r1913;
  assign w_000_1914 = r1914;
  assign w_000_1915 = r1915;
  assign w_000_1916 = r1916;
  assign w_000_1917 = r1917;
  assign w_000_1918 = r1918;
  assign w_000_1919 = r1919;
  assign w_000_1920 = r1920;
  assign w_000_1921 = r1921;
  assign w_000_1922 = r1922;
  assign w_000_1923 = r1923;
  assign w_000_1924 = r1924;
  assign w_000_1925 = r1925;
  assign w_000_1926 = r1926;
  assign w_000_1927 = r1927;
  assign w_000_1928 = r1928;
  assign w_000_1929 = r1929;
  assign w_000_1930 = r1930;
  assign w_000_1931 = r1931;
  assign w_000_1932 = r1932;
  assign w_000_1933 = r1933;
  assign w_000_1934 = r1934;
  assign w_000_1935 = r1935;
  assign w_000_1936 = r1936;
  assign w_000_1937 = r1937;
  assign w_000_1938 = r1938;
  assign w_000_1939 = r1939;
  assign w_000_1940 = r1940;
  assign w_000_1941 = r1941;
  assign w_000_1942 = r1942;
  assign w_000_1943 = r1943;
  assign w_000_1944 = r1944;
  assign w_000_1945 = r1945;
  assign w_000_1946 = r1946;
  assign w_000_1947 = r1947;
  assign w_000_1948 = r1948;
  assign w_000_1949 = r1949;
  assign w_000_1950 = r1950;
  assign w_000_1951 = r1951;
  assign w_000_1952 = r1952;
  assign w_000_1953 = r1953;
  assign w_000_1954 = r1954;
  assign w_000_1955 = r1955;
  assign w_000_1956 = r1956;
  assign w_000_1957 = r1957;
  assign w_000_1958 = r1958;
  assign w_000_1959 = r1959;
  assign w_000_1960 = r1960;
  assign w_000_1961 = r1961;
  assign w_000_1962 = r1962;
  assign w_000_1963 = r1963;
  assign w_000_1964 = r1964;
  assign w_000_1965 = r1965;
  assign w_000_1966 = r1966;
  assign w_000_1967 = r1967;
  assign w_000_1968 = r1968;
  assign w_000_1969 = r1969;
  assign w_000_1970 = r1970;
  assign w_000_1971 = r1971;
  assign w_000_1972 = r1972;
  assign w_000_1973 = r1973;
  assign w_000_1974 = r1974;
  assign w_000_1975 = r1975;
  assign w_000_1976 = r1976;
  assign w_000_1977 = r1977;
  assign w_000_1978 = r1978;
  assign w_000_1979 = r1979;
  assign w_000_1980 = r1980;
  assign w_000_1981 = r1981;
  assign w_000_1982 = r1982;
  assign w_000_1983 = r1983;
  assign w_000_1984 = r1984;
  assign w_000_1985 = r1985;
  assign w_000_1986 = r1986;
  assign w_000_1987 = r1987;
  assign w_000_1988 = r1988;
  assign w_000_1989 = r1989;
  assign w_000_1990 = r1990;
  assign w_000_1991 = r1991;
  assign w_000_1992 = r1992;
  assign w_000_1993 = r1993;
  assign w_000_1994 = r1994;
  assign w_000_1995 = r1995;
  assign w_000_1996 = r1996;
  assign w_000_1997 = r1997;

  initial begin 
    r0 = 1'b0; 
    r1 = 1'b0; 
    r2 = 1'b0; 
    r3 = 1'b0; 
    r4 = 1'b0; 
    r5 = 1'b0; 
    r6 = 1'b0; 
    r7 = 1'b0; 
    r8 = 1'b0; 
    r9 = 1'b0; 
    r10 = 1'b0; 
    r11 = 1'b0; 
    r12 = 1'b0; 
    r13 = 1'b0; 
    r14 = 1'b0; 
    r15 = 1'b0; 
    r16 = 1'b0; 
    r17 = 1'b0; 
    r18 = 1'b0; 
    r19 = 1'b0; 
    r20 = 1'b0; 
    r21 = 1'b0; 
    r22 = 1'b0; 
    r23 = 1'b0; 
    r24 = 1'b0; 
    r25 = 1'b0; 
    r26 = 1'b0; 
    r27 = 1'b0; 
    r28 = 1'b0; 
    r29 = 1'b0; 
    r30 = 1'b0; 
    r31 = 1'b0; 
    r32 = 1'b0; 
    r33 = 1'b0; 
    r34 = 1'b0; 
    r35 = 1'b0; 
    r36 = 1'b0; 
    r37 = 1'b0; 
    r38 = 1'b0; 
    r39 = 1'b0; 
    r40 = 1'b0; 
    r41 = 1'b0; 
    r42 = 1'b0; 
    r43 = 1'b0; 
    r44 = 1'b0; 
    r45 = 1'b0; 
    r46 = 1'b0; 
    r47 = 1'b0; 
    r48 = 1'b0; 
    r49 = 1'b0; 
    r50 = 1'b0; 
    r51 = 1'b0; 
    r52 = 1'b0; 
    r53 = 1'b0; 
    r54 = 1'b0; 
    r55 = 1'b0; 
    r56 = 1'b0; 
    r57 = 1'b0; 
    r58 = 1'b0; 
    r59 = 1'b0; 
    r60 = 1'b0; 
    r61 = 1'b0; 
    r62 = 1'b0; 
    r63 = 1'b0; 
    r64 = 1'b0; 
    r65 = 1'b0; 
    r66 = 1'b0; 
    r67 = 1'b0; 
    r68 = 1'b0; 
    r69 = 1'b0; 
    r70 = 1'b0; 
    r71 = 1'b0; 
    r72 = 1'b0; 
    r73 = 1'b0; 
    r74 = 1'b0; 
    r75 = 1'b0; 
    r76 = 1'b0; 
    r77 = 1'b0; 
    r78 = 1'b0; 
    r79 = 1'b0; 
    r80 = 1'b0; 
    r81 = 1'b0; 
    r82 = 1'b0; 
    r83 = 1'b0; 
    r84 = 1'b0; 
    r85 = 1'b0; 
    r86 = 1'b0; 
    r87 = 1'b0; 
    r88 = 1'b0; 
    r89 = 1'b0; 
    r90 = 1'b0; 
    r91 = 1'b0; 
    r92 = 1'b0; 
    r93 = 1'b0; 
    r94 = 1'b0; 
    r95 = 1'b0; 
    r96 = 1'b0; 
    r97 = 1'b0; 
    r98 = 1'b0; 
    r99 = 1'b0; 
    r100 = 1'b0; 
    r101 = 1'b0; 
    r102 = 1'b0; 
    r103 = 1'b0; 
    r104 = 1'b0; 
    r105 = 1'b0; 
    r106 = 1'b0; 
    r107 = 1'b0; 
    r108 = 1'b0; 
    r109 = 1'b0; 
    r110 = 1'b0; 
    r111 = 1'b0; 
    r112 = 1'b0; 
    r113 = 1'b0; 
    r114 = 1'b0; 
    r115 = 1'b0; 
    r116 = 1'b0; 
    r117 = 1'b0; 
    r118 = 1'b0; 
    r119 = 1'b0; 
    r120 = 1'b0; 
    r121 = 1'b0; 
    r122 = 1'b0; 
    r123 = 1'b0; 
    r124 = 1'b0; 
    r125 = 1'b0; 
    r126 = 1'b0; 
    r127 = 1'b0; 
    r128 = 1'b0; 
    r129 = 1'b0; 
    r130 = 1'b0; 
    r131 = 1'b0; 
    r132 = 1'b0; 
    r133 = 1'b0; 
    r134 = 1'b0; 
    r135 = 1'b0; 
    r136 = 1'b0; 
    r137 = 1'b0; 
    r138 = 1'b0; 
    r139 = 1'b0; 
    r140 = 1'b0; 
    r141 = 1'b0; 
    r142 = 1'b0; 
    r143 = 1'b0; 
    r144 = 1'b0; 
    r145 = 1'b0; 
    r146 = 1'b0; 
    r147 = 1'b0; 
    r148 = 1'b0; 
    r149 = 1'b0; 
    r150 = 1'b0; 
    r151 = 1'b0; 
    r152 = 1'b0; 
    r153 = 1'b0; 
    r154 = 1'b0; 
    r155 = 1'b0; 
    r156 = 1'b0; 
    r157 = 1'b0; 
    r158 = 1'b0; 
    r159 = 1'b0; 
    r160 = 1'b0; 
    r161 = 1'b0; 
    r162 = 1'b0; 
    r163 = 1'b0; 
    r164 = 1'b0; 
    r165 = 1'b0; 
    r166 = 1'b0; 
    r167 = 1'b0; 
    r168 = 1'b0; 
    r169 = 1'b0; 
    r170 = 1'b0; 
    r171 = 1'b0; 
    r172 = 1'b0; 
    r173 = 1'b0; 
    r174 = 1'b0; 
    r175 = 1'b0; 
    r176 = 1'b0; 
    r177 = 1'b0; 
    r178 = 1'b0; 
    r179 = 1'b0; 
    r180 = 1'b0; 
    r181 = 1'b0; 
    r182 = 1'b0; 
    r183 = 1'b0; 
    r184 = 1'b0; 
    r185 = 1'b0; 
    r186 = 1'b0; 
    r187 = 1'b0; 
    r188 = 1'b0; 
    r189 = 1'b0; 
    r190 = 1'b0; 
    r191 = 1'b0; 
    r192 = 1'b0; 
    r193 = 1'b0; 
    r194 = 1'b0; 
    r195 = 1'b0; 
    r196 = 1'b0; 
    r197 = 1'b0; 
    r198 = 1'b0; 
    r199 = 1'b0; 
    r200 = 1'b0; 
    r201 = 1'b0; 
    r202 = 1'b0; 
    r203 = 1'b0; 
    r204 = 1'b0; 
    r205 = 1'b0; 
    r206 = 1'b0; 
    r207 = 1'b0; 
    r208 = 1'b0; 
    r209 = 1'b0; 
    r210 = 1'b0; 
    r211 = 1'b0; 
    r212 = 1'b0; 
    r213 = 1'b0; 
    r214 = 1'b0; 
    r215 = 1'b0; 
    r216 = 1'b0; 
    r217 = 1'b0; 
    r218 = 1'b0; 
    r219 = 1'b0; 
    r220 = 1'b0; 
    r221 = 1'b0; 
    r222 = 1'b0; 
    r223 = 1'b0; 
    r224 = 1'b0; 
    r225 = 1'b0; 
    r226 = 1'b0; 
    r227 = 1'b0; 
    r228 = 1'b0; 
    r229 = 1'b0; 
    r230 = 1'b0; 
    r231 = 1'b0; 
    r232 = 1'b0; 
    r233 = 1'b0; 
    r234 = 1'b0; 
    r235 = 1'b0; 
    r236 = 1'b0; 
    r237 = 1'b0; 
    r238 = 1'b0; 
    r239 = 1'b0; 
    r240 = 1'b0; 
    r241 = 1'b0; 
    r242 = 1'b0; 
    r243 = 1'b0; 
    r244 = 1'b0; 
    r245 = 1'b0; 
    r246 = 1'b0; 
    r247 = 1'b0; 
    r248 = 1'b0; 
    r249 = 1'b0; 
    r250 = 1'b0; 
    r251 = 1'b0; 
    r252 = 1'b0; 
    r253 = 1'b0; 
    r254 = 1'b0; 
    r255 = 1'b0; 
    r256 = 1'b0; 
    r257 = 1'b0; 
    r258 = 1'b0; 
    r259 = 1'b0; 
    r260 = 1'b0; 
    r261 = 1'b0; 
    r262 = 1'b0; 
    r263 = 1'b0; 
    r264 = 1'b0; 
    r265 = 1'b0; 
    r266 = 1'b0; 
    r267 = 1'b0; 
    r268 = 1'b0; 
    r269 = 1'b0; 
    r270 = 1'b0; 
    r271 = 1'b0; 
    r272 = 1'b0; 
    r273 = 1'b0; 
    r274 = 1'b0; 
    r275 = 1'b0; 
    r276 = 1'b0; 
    r277 = 1'b0; 
    r278 = 1'b0; 
    r279 = 1'b0; 
    r280 = 1'b0; 
    r281 = 1'b0; 
    r282 = 1'b0; 
    r283 = 1'b0; 
    r284 = 1'b0; 
    r285 = 1'b0; 
    r286 = 1'b0; 
    r287 = 1'b0; 
    r288 = 1'b0; 
    r289 = 1'b0; 
    r290 = 1'b0; 
    r291 = 1'b0; 
    r292 = 1'b0; 
    r293 = 1'b0; 
    r294 = 1'b0; 
    r295 = 1'b0; 
    r296 = 1'b0; 
    r297 = 1'b0; 
    r298 = 1'b0; 
    r299 = 1'b0; 
    r300 = 1'b0; 
    r301 = 1'b0; 
    r302 = 1'b0; 
    r303 = 1'b0; 
    r304 = 1'b0; 
    r305 = 1'b0; 
    r306 = 1'b0; 
    r307 = 1'b0; 
    r308 = 1'b0; 
    r309 = 1'b0; 
    r310 = 1'b0; 
    r311 = 1'b0; 
    r312 = 1'b0; 
    r313 = 1'b0; 
    r314 = 1'b0; 
    r315 = 1'b0; 
    r316 = 1'b0; 
    r317 = 1'b0; 
    r318 = 1'b0; 
    r319 = 1'b0; 
    r320 = 1'b0; 
    r321 = 1'b0; 
    r322 = 1'b0; 
    r323 = 1'b0; 
    r324 = 1'b0; 
    r325 = 1'b0; 
    r326 = 1'b0; 
    r327 = 1'b0; 
    r328 = 1'b0; 
    r329 = 1'b0; 
    r330 = 1'b0; 
    r331 = 1'b0; 
    r332 = 1'b0; 
    r333 = 1'b0; 
    r334 = 1'b0; 
    r335 = 1'b0; 
    r336 = 1'b0; 
    r337 = 1'b0; 
    r338 = 1'b0; 
    r339 = 1'b0; 
    r340 = 1'b0; 
    r341 = 1'b0; 
    r342 = 1'b0; 
    r343 = 1'b0; 
    r344 = 1'b0; 
    r345 = 1'b0; 
    r346 = 1'b0; 
    r347 = 1'b0; 
    r348 = 1'b0; 
    r349 = 1'b0; 
    r350 = 1'b0; 
    r351 = 1'b0; 
    r352 = 1'b0; 
    r353 = 1'b0; 
    r354 = 1'b0; 
    r355 = 1'b0; 
    r356 = 1'b0; 
    r357 = 1'b0; 
    r358 = 1'b0; 
    r359 = 1'b0; 
    r360 = 1'b0; 
    r361 = 1'b0; 
    r362 = 1'b0; 
    r363 = 1'b0; 
    r364 = 1'b0; 
    r365 = 1'b0; 
    r366 = 1'b0; 
    r367 = 1'b0; 
    r368 = 1'b0; 
    r369 = 1'b0; 
    r370 = 1'b0; 
    r371 = 1'b0; 
    r372 = 1'b0; 
    r373 = 1'b0; 
    r374 = 1'b0; 
    r375 = 1'b0; 
    r376 = 1'b0; 
    r377 = 1'b0; 
    r378 = 1'b0; 
    r379 = 1'b0; 
    r380 = 1'b0; 
    r381 = 1'b0; 
    r382 = 1'b0; 
    r383 = 1'b0; 
    r384 = 1'b0; 
    r385 = 1'b0; 
    r386 = 1'b0; 
    r387 = 1'b0; 
    r388 = 1'b0; 
    r389 = 1'b0; 
    r390 = 1'b0; 
    r391 = 1'b0; 
    r392 = 1'b0; 
    r393 = 1'b0; 
    r394 = 1'b0; 
    r395 = 1'b0; 
    r396 = 1'b0; 
    r397 = 1'b0; 
    r398 = 1'b0; 
    r399 = 1'b0; 
    r400 = 1'b0; 
    r401 = 1'b0; 
    r402 = 1'b0; 
    r403 = 1'b0; 
    r404 = 1'b0; 
    r405 = 1'b0; 
    r406 = 1'b0; 
    r407 = 1'b0; 
    r408 = 1'b0; 
    r409 = 1'b0; 
    r410 = 1'b0; 
    r411 = 1'b0; 
    r412 = 1'b0; 
    r413 = 1'b0; 
    r414 = 1'b0; 
    r415 = 1'b0; 
    r416 = 1'b0; 
    r417 = 1'b0; 
    r418 = 1'b0; 
    r419 = 1'b0; 
    r420 = 1'b0; 
    r421 = 1'b0; 
    r422 = 1'b0; 
    r423 = 1'b0; 
    r424 = 1'b0; 
    r425 = 1'b0; 
    r426 = 1'b0; 
    r427 = 1'b0; 
    r428 = 1'b0; 
    r429 = 1'b0; 
    r430 = 1'b0; 
    r431 = 1'b0; 
    r432 = 1'b0; 
    r433 = 1'b0; 
    r434 = 1'b0; 
    r435 = 1'b0; 
    r436 = 1'b0; 
    r437 = 1'b0; 
    r438 = 1'b0; 
    r439 = 1'b0; 
    r440 = 1'b0; 
    r441 = 1'b0; 
    r442 = 1'b0; 
    r443 = 1'b0; 
    r444 = 1'b0; 
    r445 = 1'b0; 
    r446 = 1'b0; 
    r447 = 1'b0; 
    r448 = 1'b0; 
    r449 = 1'b0; 
    r450 = 1'b0; 
    r451 = 1'b0; 
    r452 = 1'b0; 
    r453 = 1'b0; 
    r454 = 1'b0; 
    r455 = 1'b0; 
    r456 = 1'b0; 
    r457 = 1'b0; 
    r458 = 1'b0; 
    r459 = 1'b0; 
    r460 = 1'b0; 
    r461 = 1'b0; 
    r462 = 1'b0; 
    r463 = 1'b0; 
    r464 = 1'b0; 
    r465 = 1'b0; 
    r466 = 1'b0; 
    r467 = 1'b0; 
    r468 = 1'b0; 
    r469 = 1'b0; 
    r470 = 1'b0; 
    r471 = 1'b0; 
    r472 = 1'b0; 
    r473 = 1'b0; 
    r474 = 1'b0; 
    r475 = 1'b0; 
    r476 = 1'b0; 
    r477 = 1'b0; 
    r478 = 1'b0; 
    r479 = 1'b0; 
    r480 = 1'b0; 
    r481 = 1'b0; 
    r482 = 1'b0; 
    r483 = 1'b0; 
    r484 = 1'b0; 
    r485 = 1'b0; 
    r486 = 1'b0; 
    r487 = 1'b0; 
    r488 = 1'b0; 
    r489 = 1'b0; 
    r490 = 1'b0; 
    r491 = 1'b0; 
    r492 = 1'b0; 
    r493 = 1'b0; 
    r494 = 1'b0; 
    r495 = 1'b0; 
    r496 = 1'b0; 
    r497 = 1'b0; 
    r498 = 1'b0; 
    r499 = 1'b0; 
    r500 = 1'b0; 
    r501 = 1'b0; 
    r502 = 1'b0; 
    r503 = 1'b0; 
    r504 = 1'b0; 
    r505 = 1'b0; 
    r506 = 1'b0; 
    r507 = 1'b0; 
    r508 = 1'b0; 
    r509 = 1'b0; 
    r510 = 1'b0; 
    r511 = 1'b0; 
    r512 = 1'b0; 
    r513 = 1'b0; 
    r514 = 1'b0; 
    r515 = 1'b0; 
    r516 = 1'b0; 
    r517 = 1'b0; 
    r518 = 1'b0; 
    r519 = 1'b0; 
    r520 = 1'b0; 
    r521 = 1'b0; 
    r522 = 1'b0; 
    r523 = 1'b0; 
    r524 = 1'b0; 
    r525 = 1'b0; 
    r526 = 1'b0; 
    r527 = 1'b0; 
    r528 = 1'b0; 
    r529 = 1'b0; 
    r530 = 1'b0; 
    r531 = 1'b0; 
    r532 = 1'b0; 
    r533 = 1'b0; 
    r534 = 1'b0; 
    r535 = 1'b0; 
    r536 = 1'b0; 
    r537 = 1'b0; 
    r538 = 1'b0; 
    r539 = 1'b0; 
    r540 = 1'b0; 
    r541 = 1'b0; 
    r542 = 1'b0; 
    r543 = 1'b0; 
    r544 = 1'b0; 
    r545 = 1'b0; 
    r546 = 1'b0; 
    r547 = 1'b0; 
    r548 = 1'b0; 
    r549 = 1'b0; 
    r550 = 1'b0; 
    r551 = 1'b0; 
    r552 = 1'b0; 
    r553 = 1'b0; 
    r554 = 1'b0; 
    r555 = 1'b0; 
    r556 = 1'b0; 
    r557 = 1'b0; 
    r558 = 1'b0; 
    r559 = 1'b0; 
    r560 = 1'b0; 
    r561 = 1'b0; 
    r562 = 1'b0; 
    r563 = 1'b0; 
    r564 = 1'b0; 
    r565 = 1'b0; 
    r566 = 1'b0; 
    r567 = 1'b0; 
    r568 = 1'b0; 
    r569 = 1'b0; 
    r570 = 1'b0; 
    r571 = 1'b0; 
    r572 = 1'b0; 
    r573 = 1'b0; 
    r574 = 1'b0; 
    r575 = 1'b0; 
    r576 = 1'b0; 
    r577 = 1'b0; 
    r578 = 1'b0; 
    r579 = 1'b0; 
    r580 = 1'b0; 
    r581 = 1'b0; 
    r582 = 1'b0; 
    r583 = 1'b0; 
    r584 = 1'b0; 
    r585 = 1'b0; 
    r586 = 1'b0; 
    r587 = 1'b0; 
    r588 = 1'b0; 
    r589 = 1'b0; 
    r590 = 1'b0; 
    r591 = 1'b0; 
    r592 = 1'b0; 
    r593 = 1'b0; 
    r594 = 1'b0; 
    r595 = 1'b0; 
    r596 = 1'b0; 
    r597 = 1'b0; 
    r598 = 1'b0; 
    r599 = 1'b0; 
    r600 = 1'b0; 
    r601 = 1'b0; 
    r602 = 1'b0; 
    r603 = 1'b0; 
    r604 = 1'b0; 
    r605 = 1'b0; 
    r606 = 1'b0; 
    r607 = 1'b0; 
    r608 = 1'b0; 
    r609 = 1'b0; 
    r610 = 1'b0; 
    r611 = 1'b0; 
    r612 = 1'b0; 
    r613 = 1'b0; 
    r614 = 1'b0; 
    r615 = 1'b0; 
    r616 = 1'b0; 
    r617 = 1'b0; 
    r618 = 1'b0; 
    r619 = 1'b0; 
    r620 = 1'b0; 
    r621 = 1'b0; 
    r622 = 1'b0; 
    r623 = 1'b0; 
    r624 = 1'b0; 
    r625 = 1'b0; 
    r626 = 1'b0; 
    r627 = 1'b0; 
    r628 = 1'b0; 
    r629 = 1'b0; 
    r630 = 1'b0; 
    r631 = 1'b0; 
    r632 = 1'b0; 
    r633 = 1'b0; 
    r634 = 1'b0; 
    r635 = 1'b0; 
    r636 = 1'b0; 
    r637 = 1'b0; 
    r638 = 1'b0; 
    r639 = 1'b0; 
    r640 = 1'b0; 
    r641 = 1'b0; 
    r642 = 1'b0; 
    r643 = 1'b0; 
    r644 = 1'b0; 
    r645 = 1'b0; 
    r646 = 1'b0; 
    r647 = 1'b0; 
    r648 = 1'b0; 
    r649 = 1'b0; 
    r650 = 1'b0; 
    r651 = 1'b0; 
    r652 = 1'b0; 
    r653 = 1'b0; 
    r654 = 1'b0; 
    r655 = 1'b0; 
    r656 = 1'b0; 
    r657 = 1'b0; 
    r658 = 1'b0; 
    r659 = 1'b0; 
    r660 = 1'b0; 
    r661 = 1'b0; 
    r662 = 1'b0; 
    r663 = 1'b0; 
    r664 = 1'b0; 
    r665 = 1'b0; 
    r666 = 1'b0; 
    r667 = 1'b0; 
    r668 = 1'b0; 
    r669 = 1'b0; 
    r670 = 1'b0; 
    r671 = 1'b0; 
    r672 = 1'b0; 
    r673 = 1'b0; 
    r674 = 1'b0; 
    r675 = 1'b0; 
    r676 = 1'b0; 
    r677 = 1'b0; 
    r678 = 1'b0; 
    r679 = 1'b0; 
    r680 = 1'b0; 
    r681 = 1'b0; 
    r682 = 1'b0; 
    r683 = 1'b0; 
    r684 = 1'b0; 
    r685 = 1'b0; 
    r686 = 1'b0; 
    r687 = 1'b0; 
    r688 = 1'b0; 
    r689 = 1'b0; 
    r690 = 1'b0; 
    r691 = 1'b0; 
    r692 = 1'b0; 
    r693 = 1'b0; 
    r694 = 1'b0; 
    r695 = 1'b0; 
    r696 = 1'b0; 
    r697 = 1'b0; 
    r698 = 1'b0; 
    r699 = 1'b0; 
    r700 = 1'b0; 
    r701 = 1'b0; 
    r702 = 1'b0; 
    r703 = 1'b0; 
    r704 = 1'b0; 
    r705 = 1'b0; 
    r706 = 1'b0; 
    r707 = 1'b0; 
    r708 = 1'b0; 
    r709 = 1'b0; 
    r710 = 1'b0; 
    r711 = 1'b0; 
    r712 = 1'b0; 
    r713 = 1'b0; 
    r714 = 1'b0; 
    r715 = 1'b0; 
    r716 = 1'b0; 
    r717 = 1'b0; 
    r718 = 1'b0; 
    r719 = 1'b0; 
    r720 = 1'b0; 
    r721 = 1'b0; 
    r722 = 1'b0; 
    r723 = 1'b0; 
    r724 = 1'b0; 
    r725 = 1'b0; 
    r726 = 1'b0; 
    r727 = 1'b0; 
    r728 = 1'b0; 
    r729 = 1'b0; 
    r730 = 1'b0; 
    r731 = 1'b0; 
    r732 = 1'b0; 
    r733 = 1'b0; 
    r734 = 1'b0; 
    r735 = 1'b0; 
    r736 = 1'b0; 
    r737 = 1'b0; 
    r738 = 1'b0; 
    r739 = 1'b0; 
    r740 = 1'b0; 
    r741 = 1'b0; 
    r742 = 1'b0; 
    r743 = 1'b0; 
    r744 = 1'b0; 
    r745 = 1'b0; 
    r746 = 1'b0; 
    r747 = 1'b0; 
    r748 = 1'b0; 
    r749 = 1'b0; 
    r750 = 1'b0; 
    r751 = 1'b0; 
    r752 = 1'b0; 
    r753 = 1'b0; 
    r754 = 1'b0; 
    r755 = 1'b0; 
    r756 = 1'b0; 
    r757 = 1'b0; 
    r758 = 1'b0; 
    r759 = 1'b0; 
    r760 = 1'b0; 
    r761 = 1'b0; 
    r762 = 1'b0; 
    r763 = 1'b0; 
    r764 = 1'b0; 
    r765 = 1'b0; 
    r766 = 1'b0; 
    r767 = 1'b0; 
    r768 = 1'b0; 
    r769 = 1'b0; 
    r770 = 1'b0; 
    r771 = 1'b0; 
    r772 = 1'b0; 
    r773 = 1'b0; 
    r774 = 1'b0; 
    r775 = 1'b0; 
    r776 = 1'b0; 
    r777 = 1'b0; 
    r778 = 1'b0; 
    r779 = 1'b0; 
    r780 = 1'b0; 
    r781 = 1'b0; 
    r782 = 1'b0; 
    r783 = 1'b0; 
    r784 = 1'b0; 
    r785 = 1'b0; 
    r786 = 1'b0; 
    r787 = 1'b0; 
    r788 = 1'b0; 
    r789 = 1'b0; 
    r790 = 1'b0; 
    r791 = 1'b0; 
    r792 = 1'b0; 
    r793 = 1'b0; 
    r794 = 1'b0; 
    r795 = 1'b0; 
    r796 = 1'b0; 
    r797 = 1'b0; 
    r798 = 1'b0; 
    r799 = 1'b0; 
    r800 = 1'b0; 
    r801 = 1'b0; 
    r802 = 1'b0; 
    r803 = 1'b0; 
    r804 = 1'b0; 
    r805 = 1'b0; 
    r806 = 1'b0; 
    r807 = 1'b0; 
    r808 = 1'b0; 
    r809 = 1'b0; 
    r810 = 1'b0; 
    r811 = 1'b0; 
    r812 = 1'b0; 
    r813 = 1'b0; 
    r814 = 1'b0; 
    r815 = 1'b0; 
    r816 = 1'b0; 
    r817 = 1'b0; 
    r818 = 1'b0; 
    r819 = 1'b0; 
    r820 = 1'b0; 
    r821 = 1'b0; 
    r822 = 1'b0; 
    r823 = 1'b0; 
    r824 = 1'b0; 
    r825 = 1'b0; 
    r826 = 1'b0; 
    r827 = 1'b0; 
    r828 = 1'b0; 
    r829 = 1'b0; 
    r830 = 1'b0; 
    r831 = 1'b0; 
    r832 = 1'b0; 
    r833 = 1'b0; 
    r834 = 1'b0; 
    r835 = 1'b0; 
    r836 = 1'b0; 
    r837 = 1'b0; 
    r838 = 1'b0; 
    r839 = 1'b0; 
    r840 = 1'b0; 
    r841 = 1'b0; 
    r842 = 1'b0; 
    r843 = 1'b0; 
    r844 = 1'b0; 
    r845 = 1'b0; 
    r846 = 1'b0; 
    r847 = 1'b0; 
    r848 = 1'b0; 
    r849 = 1'b0; 
    r850 = 1'b0; 
    r851 = 1'b0; 
    r852 = 1'b0; 
    r853 = 1'b0; 
    r854 = 1'b0; 
    r855 = 1'b0; 
    r856 = 1'b0; 
    r857 = 1'b0; 
    r858 = 1'b0; 
    r859 = 1'b0; 
    r860 = 1'b0; 
    r861 = 1'b0; 
    r862 = 1'b0; 
    r863 = 1'b0; 
    r864 = 1'b0; 
    r865 = 1'b0; 
    r866 = 1'b0; 
    r867 = 1'b0; 
    r868 = 1'b0; 
    r869 = 1'b0; 
    r870 = 1'b0; 
    r871 = 1'b0; 
    r872 = 1'b0; 
    r873 = 1'b0; 
    r874 = 1'b0; 
    r875 = 1'b0; 
    r876 = 1'b0; 
    r877 = 1'b0; 
    r878 = 1'b0; 
    r879 = 1'b0; 
    r880 = 1'b0; 
    r881 = 1'b0; 
    r882 = 1'b0; 
    r883 = 1'b0; 
    r884 = 1'b0; 
    r885 = 1'b0; 
    r886 = 1'b0; 
    r887 = 1'b0; 
    r888 = 1'b0; 
    r889 = 1'b0; 
    r890 = 1'b0; 
    r891 = 1'b0; 
    r892 = 1'b0; 
    r893 = 1'b0; 
    r894 = 1'b0; 
    r895 = 1'b0; 
    r896 = 1'b0; 
    r897 = 1'b0; 
    r898 = 1'b0; 
    r899 = 1'b0; 
    r900 = 1'b0; 
    r901 = 1'b0; 
    r902 = 1'b0; 
    r903 = 1'b0; 
    r904 = 1'b0; 
    r905 = 1'b0; 
    r906 = 1'b0; 
    r907 = 1'b0; 
    r908 = 1'b0; 
    r909 = 1'b0; 
    r910 = 1'b0; 
    r911 = 1'b0; 
    r912 = 1'b0; 
    r913 = 1'b0; 
    r914 = 1'b0; 
    r915 = 1'b0; 
    r916 = 1'b0; 
    r917 = 1'b0; 
    r918 = 1'b0; 
    r919 = 1'b0; 
    r920 = 1'b0; 
    r921 = 1'b0; 
    r922 = 1'b0; 
    r923 = 1'b0; 
    r924 = 1'b0; 
    r925 = 1'b0; 
    r926 = 1'b0; 
    r927 = 1'b0; 
    r928 = 1'b0; 
    r929 = 1'b0; 
    r930 = 1'b0; 
    r931 = 1'b0; 
    r932 = 1'b0; 
    r933 = 1'b0; 
    r934 = 1'b0; 
    r935 = 1'b0; 
    r936 = 1'b0; 
    r937 = 1'b0; 
    r938 = 1'b0; 
    r939 = 1'b0; 
    r940 = 1'b0; 
    r941 = 1'b0; 
    r942 = 1'b0; 
    r943 = 1'b0; 
    r944 = 1'b0; 
    r945 = 1'b0; 
    r946 = 1'b0; 
    r947 = 1'b0; 
    r948 = 1'b0; 
    r949 = 1'b0; 
    r950 = 1'b0; 
    r951 = 1'b0; 
    r952 = 1'b0; 
    r953 = 1'b0; 
    r954 = 1'b0; 
    r955 = 1'b0; 
    r956 = 1'b0; 
    r957 = 1'b0; 
    r958 = 1'b0; 
    r959 = 1'b0; 
    r960 = 1'b0; 
    r961 = 1'b0; 
    r962 = 1'b0; 
    r963 = 1'b0; 
    r964 = 1'b0; 
    r965 = 1'b0; 
    r966 = 1'b0; 
    r967 = 1'b0; 
    r968 = 1'b0; 
    r969 = 1'b0; 
    r970 = 1'b0; 
    r971 = 1'b0; 
    r972 = 1'b0; 
    r973 = 1'b0; 
    r974 = 1'b0; 
    r975 = 1'b0; 
    r976 = 1'b0; 
    r977 = 1'b0; 
    r978 = 1'b0; 
    r979 = 1'b0; 
    r980 = 1'b0; 
    r981 = 1'b0; 
    r982 = 1'b0; 
    r983 = 1'b0; 
    r984 = 1'b0; 
    r985 = 1'b0; 
    r986 = 1'b0; 
    r987 = 1'b0; 
    r988 = 1'b0; 
    r989 = 1'b0; 
    r990 = 1'b0; 
    r991 = 1'b0; 
    r992 = 1'b0; 
    r993 = 1'b0; 
    r994 = 1'b0; 
    r995 = 1'b0; 
    r996 = 1'b0; 
    r997 = 1'b0; 
    r998 = 1'b0; 
    r999 = 1'b0; 
    r1000 = 1'b0; 
    r1001 = 1'b0; 
    r1002 = 1'b0; 
    r1003 = 1'b0; 
    r1004 = 1'b0; 
    r1005 = 1'b0; 
    r1006 = 1'b0; 
    r1007 = 1'b0; 
    r1008 = 1'b0; 
    r1009 = 1'b0; 
    r1010 = 1'b0; 
    r1011 = 1'b0; 
    r1012 = 1'b0; 
    r1013 = 1'b0; 
    r1014 = 1'b0; 
    r1015 = 1'b0; 
    r1016 = 1'b0; 
    r1017 = 1'b0; 
    r1018 = 1'b0; 
    r1019 = 1'b0; 
    r1020 = 1'b0; 
    r1021 = 1'b0; 
    r1022 = 1'b0; 
    r1023 = 1'b0; 
    r1024 = 1'b0; 
    r1025 = 1'b0; 
    r1026 = 1'b0; 
    r1027 = 1'b0; 
    r1028 = 1'b0; 
    r1029 = 1'b0; 
    r1030 = 1'b0; 
    r1031 = 1'b0; 
    r1032 = 1'b0; 
    r1033 = 1'b0; 
    r1034 = 1'b0; 
    r1035 = 1'b0; 
    r1036 = 1'b0; 
    r1037 = 1'b0; 
    r1038 = 1'b0; 
    r1039 = 1'b0; 
    r1040 = 1'b0; 
    r1041 = 1'b0; 
    r1042 = 1'b0; 
    r1043 = 1'b0; 
    r1044 = 1'b0; 
    r1045 = 1'b0; 
    r1046 = 1'b0; 
    r1047 = 1'b0; 
    r1048 = 1'b0; 
    r1049 = 1'b0; 
    r1050 = 1'b0; 
    r1051 = 1'b0; 
    r1052 = 1'b0; 
    r1053 = 1'b0; 
    r1054 = 1'b0; 
    r1055 = 1'b0; 
    r1056 = 1'b0; 
    r1057 = 1'b0; 
    r1058 = 1'b0; 
    r1059 = 1'b0; 
    r1060 = 1'b0; 
    r1061 = 1'b0; 
    r1062 = 1'b0; 
    r1063 = 1'b0; 
    r1064 = 1'b0; 
    r1065 = 1'b0; 
    r1066 = 1'b0; 
    r1067 = 1'b0; 
    r1068 = 1'b0; 
    r1069 = 1'b0; 
    r1070 = 1'b0; 
    r1071 = 1'b0; 
    r1072 = 1'b0; 
    r1073 = 1'b0; 
    r1074 = 1'b0; 
    r1075 = 1'b0; 
    r1076 = 1'b0; 
    r1077 = 1'b0; 
    r1078 = 1'b0; 
    r1079 = 1'b0; 
    r1080 = 1'b0; 
    r1081 = 1'b0; 
    r1082 = 1'b0; 
    r1083 = 1'b0; 
    r1084 = 1'b0; 
    r1085 = 1'b0; 
    r1086 = 1'b0; 
    r1087 = 1'b0; 
    r1088 = 1'b0; 
    r1089 = 1'b0; 
    r1090 = 1'b0; 
    r1091 = 1'b0; 
    r1092 = 1'b0; 
    r1093 = 1'b0; 
    r1094 = 1'b0; 
    r1095 = 1'b0; 
    r1096 = 1'b0; 
    r1097 = 1'b0; 
    r1098 = 1'b0; 
    r1099 = 1'b0; 
    r1100 = 1'b0; 
    r1101 = 1'b0; 
    r1102 = 1'b0; 
    r1103 = 1'b0; 
    r1104 = 1'b0; 
    r1105 = 1'b0; 
    r1106 = 1'b0; 
    r1107 = 1'b0; 
    r1108 = 1'b0; 
    r1109 = 1'b0; 
    r1110 = 1'b0; 
    r1111 = 1'b0; 
    r1112 = 1'b0; 
    r1113 = 1'b0; 
    r1114 = 1'b0; 
    r1115 = 1'b0; 
    r1116 = 1'b0; 
    r1117 = 1'b0; 
    r1118 = 1'b0; 
    r1119 = 1'b0; 
    r1120 = 1'b0; 
    r1121 = 1'b0; 
    r1122 = 1'b0; 
    r1123 = 1'b0; 
    r1124 = 1'b0; 
    r1125 = 1'b0; 
    r1126 = 1'b0; 
    r1127 = 1'b0; 
    r1128 = 1'b0; 
    r1129 = 1'b0; 
    r1130 = 1'b0; 
    r1131 = 1'b0; 
    r1132 = 1'b0; 
    r1133 = 1'b0; 
    r1134 = 1'b0; 
    r1135 = 1'b0; 
    r1136 = 1'b0; 
    r1137 = 1'b0; 
    r1138 = 1'b0; 
    r1139 = 1'b0; 
    r1140 = 1'b0; 
    r1141 = 1'b0; 
    r1142 = 1'b0; 
    r1143 = 1'b0; 
    r1144 = 1'b0; 
    r1145 = 1'b0; 
    r1146 = 1'b0; 
    r1147 = 1'b0; 
    r1148 = 1'b0; 
    r1149 = 1'b0; 
    r1150 = 1'b0; 
    r1151 = 1'b0; 
    r1152 = 1'b0; 
    r1153 = 1'b0; 
    r1154 = 1'b0; 
    r1155 = 1'b0; 
    r1156 = 1'b0; 
    r1157 = 1'b0; 
    r1158 = 1'b0; 
    r1159 = 1'b0; 
    r1160 = 1'b0; 
    r1161 = 1'b0; 
    r1162 = 1'b0; 
    r1163 = 1'b0; 
    r1164 = 1'b0; 
    r1165 = 1'b0; 
    r1166 = 1'b0; 
    r1167 = 1'b0; 
    r1168 = 1'b0; 
    r1169 = 1'b0; 
    r1170 = 1'b0; 
    r1171 = 1'b0; 
    r1172 = 1'b0; 
    r1173 = 1'b0; 
    r1174 = 1'b0; 
    r1175 = 1'b0; 
    r1176 = 1'b0; 
    r1177 = 1'b0; 
    r1178 = 1'b0; 
    r1179 = 1'b0; 
    r1180 = 1'b0; 
    r1181 = 1'b0; 
    r1182 = 1'b0; 
    r1183 = 1'b0; 
    r1184 = 1'b0; 
    r1185 = 1'b0; 
    r1186 = 1'b0; 
    r1187 = 1'b0; 
    r1188 = 1'b0; 
    r1189 = 1'b0; 
    r1190 = 1'b0; 
    r1191 = 1'b0; 
    r1192 = 1'b0; 
    r1193 = 1'b0; 
    r1194 = 1'b0; 
    r1195 = 1'b0; 
    r1196 = 1'b0; 
    r1197 = 1'b0; 
    r1198 = 1'b0; 
    r1199 = 1'b0; 
    r1200 = 1'b0; 
    r1201 = 1'b0; 
    r1202 = 1'b0; 
    r1203 = 1'b0; 
    r1204 = 1'b0; 
    r1205 = 1'b0; 
    r1206 = 1'b0; 
    r1207 = 1'b0; 
    r1208 = 1'b0; 
    r1209 = 1'b0; 
    r1210 = 1'b0; 
    r1211 = 1'b0; 
    r1212 = 1'b0; 
    r1213 = 1'b0; 
    r1214 = 1'b0; 
    r1215 = 1'b0; 
    r1216 = 1'b0; 
    r1217 = 1'b0; 
    r1218 = 1'b0; 
    r1219 = 1'b0; 
    r1220 = 1'b0; 
    r1221 = 1'b0; 
    r1222 = 1'b0; 
    r1223 = 1'b0; 
    r1224 = 1'b0; 
    r1225 = 1'b0; 
    r1226 = 1'b0; 
    r1227 = 1'b0; 
    r1228 = 1'b0; 
    r1229 = 1'b0; 
    r1230 = 1'b0; 
    r1231 = 1'b0; 
    r1232 = 1'b0; 
    r1233 = 1'b0; 
    r1234 = 1'b0; 
    r1235 = 1'b0; 
    r1236 = 1'b0; 
    r1237 = 1'b0; 
    r1238 = 1'b0; 
    r1239 = 1'b0; 
    r1240 = 1'b0; 
    r1241 = 1'b0; 
    r1242 = 1'b0; 
    r1243 = 1'b0; 
    r1244 = 1'b0; 
    r1245 = 1'b0; 
    r1246 = 1'b0; 
    r1247 = 1'b0; 
    r1248 = 1'b0; 
    r1249 = 1'b0; 
    r1250 = 1'b0; 
    r1251 = 1'b0; 
    r1252 = 1'b0; 
    r1253 = 1'b0; 
    r1254 = 1'b0; 
    r1255 = 1'b0; 
    r1256 = 1'b0; 
    r1257 = 1'b0; 
    r1258 = 1'b0; 
    r1259 = 1'b0; 
    r1260 = 1'b0; 
    r1261 = 1'b0; 
    r1262 = 1'b0; 
    r1263 = 1'b0; 
    r1264 = 1'b0; 
    r1265 = 1'b0; 
    r1266 = 1'b0; 
    r1267 = 1'b0; 
    r1268 = 1'b0; 
    r1269 = 1'b0; 
    r1270 = 1'b0; 
    r1271 = 1'b0; 
    r1272 = 1'b0; 
    r1273 = 1'b0; 
    r1274 = 1'b0; 
    r1275 = 1'b0; 
    r1276 = 1'b0; 
    r1277 = 1'b0; 
    r1278 = 1'b0; 
    r1279 = 1'b0; 
    r1280 = 1'b0; 
    r1281 = 1'b0; 
    r1282 = 1'b0; 
    r1283 = 1'b0; 
    r1284 = 1'b0; 
    r1285 = 1'b0; 
    r1286 = 1'b0; 
    r1287 = 1'b0; 
    r1288 = 1'b0; 
    r1289 = 1'b0; 
    r1290 = 1'b0; 
    r1291 = 1'b0; 
    r1292 = 1'b0; 
    r1293 = 1'b0; 
    r1294 = 1'b0; 
    r1295 = 1'b0; 
    r1296 = 1'b0; 
    r1297 = 1'b0; 
    r1298 = 1'b0; 
    r1299 = 1'b0; 
    r1300 = 1'b0; 
    r1301 = 1'b0; 
    r1302 = 1'b0; 
    r1303 = 1'b0; 
    r1304 = 1'b0; 
    r1305 = 1'b0; 
    r1306 = 1'b0; 
    r1307 = 1'b0; 
    r1308 = 1'b0; 
    r1309 = 1'b0; 
    r1310 = 1'b0; 
    r1311 = 1'b0; 
    r1312 = 1'b0; 
    r1313 = 1'b0; 
    r1314 = 1'b0; 
    r1315 = 1'b0; 
    r1316 = 1'b0; 
    r1317 = 1'b0; 
    r1318 = 1'b0; 
    r1319 = 1'b0; 
    r1320 = 1'b0; 
    r1321 = 1'b0; 
    r1322 = 1'b0; 
    r1323 = 1'b0; 
    r1324 = 1'b0; 
    r1325 = 1'b0; 
    r1326 = 1'b0; 
    r1327 = 1'b0; 
    r1328 = 1'b0; 
    r1329 = 1'b0; 
    r1330 = 1'b0; 
    r1331 = 1'b0; 
    r1332 = 1'b0; 
    r1333 = 1'b0; 
    r1334 = 1'b0; 
    r1335 = 1'b0; 
    r1336 = 1'b0; 
    r1337 = 1'b0; 
    r1338 = 1'b0; 
    r1339 = 1'b0; 
    r1340 = 1'b0; 
    r1341 = 1'b0; 
    r1342 = 1'b0; 
    r1343 = 1'b0; 
    r1344 = 1'b0; 
    r1345 = 1'b0; 
    r1346 = 1'b0; 
    r1347 = 1'b0; 
    r1348 = 1'b0; 
    r1349 = 1'b0; 
    r1350 = 1'b0; 
    r1351 = 1'b0; 
    r1352 = 1'b0; 
    r1353 = 1'b0; 
    r1354 = 1'b0; 
    r1355 = 1'b0; 
    r1356 = 1'b0; 
    r1357 = 1'b0; 
    r1358 = 1'b0; 
    r1359 = 1'b0; 
    r1360 = 1'b0; 
    r1361 = 1'b0; 
    r1362 = 1'b0; 
    r1363 = 1'b0; 
    r1364 = 1'b0; 
    r1365 = 1'b0; 
    r1366 = 1'b0; 
    r1367 = 1'b0; 
    r1368 = 1'b0; 
    r1369 = 1'b0; 
    r1370 = 1'b0; 
    r1371 = 1'b0; 
    r1372 = 1'b0; 
    r1373 = 1'b0; 
    r1374 = 1'b0; 
    r1375 = 1'b0; 
    r1376 = 1'b0; 
    r1377 = 1'b0; 
    r1378 = 1'b0; 
    r1379 = 1'b0; 
    r1380 = 1'b0; 
    r1381 = 1'b0; 
    r1382 = 1'b0; 
    r1383 = 1'b0; 
    r1384 = 1'b0; 
    r1385 = 1'b0; 
    r1386 = 1'b0; 
    r1387 = 1'b0; 
    r1388 = 1'b0; 
    r1389 = 1'b0; 
    r1390 = 1'b0; 
    r1391 = 1'b0; 
    r1392 = 1'b0; 
    r1393 = 1'b0; 
    r1394 = 1'b0; 
    r1395 = 1'b0; 
    r1396 = 1'b0; 
    r1397 = 1'b0; 
    r1398 = 1'b0; 
    r1399 = 1'b0; 
    r1400 = 1'b0; 
    r1401 = 1'b0; 
    r1402 = 1'b0; 
    r1403 = 1'b0; 
    r1404 = 1'b0; 
    r1405 = 1'b0; 
    r1406 = 1'b0; 
    r1407 = 1'b0; 
    r1408 = 1'b0; 
    r1409 = 1'b0; 
    r1410 = 1'b0; 
    r1411 = 1'b0; 
    r1412 = 1'b0; 
    r1413 = 1'b0; 
    r1414 = 1'b0; 
    r1415 = 1'b0; 
    r1416 = 1'b0; 
    r1417 = 1'b0; 
    r1418 = 1'b0; 
    r1419 = 1'b0; 
    r1420 = 1'b0; 
    r1421 = 1'b0; 
    r1422 = 1'b0; 
    r1423 = 1'b0; 
    r1424 = 1'b0; 
    r1425 = 1'b0; 
    r1426 = 1'b0; 
    r1427 = 1'b0; 
    r1428 = 1'b0; 
    r1429 = 1'b0; 
    r1430 = 1'b0; 
    r1431 = 1'b0; 
    r1432 = 1'b0; 
    r1433 = 1'b0; 
    r1434 = 1'b0; 
    r1435 = 1'b0; 
    r1436 = 1'b0; 
    r1437 = 1'b0; 
    r1438 = 1'b0; 
    r1439 = 1'b0; 
    r1440 = 1'b0; 
    r1441 = 1'b0; 
    r1442 = 1'b0; 
    r1443 = 1'b0; 
    r1444 = 1'b0; 
    r1445 = 1'b0; 
    r1446 = 1'b0; 
    r1447 = 1'b0; 
    r1448 = 1'b0; 
    r1449 = 1'b0; 
    r1450 = 1'b0; 
    r1451 = 1'b0; 
    r1452 = 1'b0; 
    r1453 = 1'b0; 
    r1454 = 1'b0; 
    r1455 = 1'b0; 
    r1456 = 1'b0; 
    r1457 = 1'b0; 
    r1458 = 1'b0; 
    r1459 = 1'b0; 
    r1460 = 1'b0; 
    r1461 = 1'b0; 
    r1462 = 1'b0; 
    r1463 = 1'b0; 
    r1464 = 1'b0; 
    r1465 = 1'b0; 
    r1466 = 1'b0; 
    r1467 = 1'b0; 
    r1468 = 1'b0; 
    r1469 = 1'b0; 
    r1470 = 1'b0; 
    r1471 = 1'b0; 
    r1472 = 1'b0; 
    r1473 = 1'b0; 
    r1474 = 1'b0; 
    r1475 = 1'b0; 
    r1476 = 1'b0; 
    r1477 = 1'b0; 
    r1478 = 1'b0; 
    r1479 = 1'b0; 
    r1480 = 1'b0; 
    r1481 = 1'b0; 
    r1482 = 1'b0; 
    r1483 = 1'b0; 
    r1484 = 1'b0; 
    r1485 = 1'b0; 
    r1486 = 1'b0; 
    r1487 = 1'b0; 
    r1488 = 1'b0; 
    r1489 = 1'b0; 
    r1490 = 1'b0; 
    r1491 = 1'b0; 
    r1492 = 1'b0; 
    r1493 = 1'b0; 
    r1494 = 1'b0; 
    r1495 = 1'b0; 
    r1496 = 1'b0; 
    r1497 = 1'b0; 
    r1498 = 1'b0; 
    r1499 = 1'b0; 
    r1500 = 1'b0; 
    r1501 = 1'b0; 
    r1502 = 1'b0; 
    r1503 = 1'b0; 
    r1504 = 1'b0; 
    r1505 = 1'b0; 
    r1506 = 1'b0; 
    r1507 = 1'b0; 
    r1508 = 1'b0; 
    r1509 = 1'b0; 
    r1510 = 1'b0; 
    r1511 = 1'b0; 
    r1512 = 1'b0; 
    r1513 = 1'b0; 
    r1514 = 1'b0; 
    r1515 = 1'b0; 
    r1516 = 1'b0; 
    r1517 = 1'b0; 
    r1518 = 1'b0; 
    r1519 = 1'b0; 
    r1520 = 1'b0; 
    r1521 = 1'b0; 
    r1522 = 1'b0; 
    r1523 = 1'b0; 
    r1524 = 1'b0; 
    r1525 = 1'b0; 
    r1526 = 1'b0; 
    r1527 = 1'b0; 
    r1528 = 1'b0; 
    r1529 = 1'b0; 
    r1530 = 1'b0; 
    r1531 = 1'b0; 
    r1532 = 1'b0; 
    r1533 = 1'b0; 
    r1534 = 1'b0; 
    r1535 = 1'b0; 
    r1536 = 1'b0; 
    r1537 = 1'b0; 
    r1538 = 1'b0; 
    r1539 = 1'b0; 
    r1540 = 1'b0; 
    r1541 = 1'b0; 
    r1542 = 1'b0; 
    r1543 = 1'b0; 
    r1544 = 1'b0; 
    r1545 = 1'b0; 
    r1546 = 1'b0; 
    r1547 = 1'b0; 
    r1548 = 1'b0; 
    r1549 = 1'b0; 
    r1550 = 1'b0; 
    r1551 = 1'b0; 
    r1552 = 1'b0; 
    r1553 = 1'b0; 
    r1554 = 1'b0; 
    r1555 = 1'b0; 
    r1556 = 1'b0; 
    r1557 = 1'b0; 
    r1558 = 1'b0; 
    r1559 = 1'b0; 
    r1560 = 1'b0; 
    r1561 = 1'b0; 
    r1562 = 1'b0; 
    r1563 = 1'b0; 
    r1564 = 1'b0; 
    r1565 = 1'b0; 
    r1566 = 1'b0; 
    r1567 = 1'b0; 
    r1568 = 1'b0; 
    r1569 = 1'b0; 
    r1570 = 1'b0; 
    r1571 = 1'b0; 
    r1572 = 1'b0; 
    r1573 = 1'b0; 
    r1574 = 1'b0; 
    r1575 = 1'b0; 
    r1576 = 1'b0; 
    r1577 = 1'b0; 
    r1578 = 1'b0; 
    r1579 = 1'b0; 
    r1580 = 1'b0; 
    r1581 = 1'b0; 
    r1582 = 1'b0; 
    r1583 = 1'b0; 
    r1584 = 1'b0; 
    r1585 = 1'b0; 
    r1586 = 1'b0; 
    r1587 = 1'b0; 
    r1588 = 1'b0; 
    r1589 = 1'b0; 
    r1590 = 1'b0; 
    r1591 = 1'b0; 
    r1592 = 1'b0; 
    r1593 = 1'b0; 
    r1594 = 1'b0; 
    r1595 = 1'b0; 
    r1596 = 1'b0; 
    r1597 = 1'b0; 
    r1598 = 1'b0; 
    r1599 = 1'b0; 
    r1600 = 1'b0; 
    r1601 = 1'b0; 
    r1602 = 1'b0; 
    r1603 = 1'b0; 
    r1604 = 1'b0; 
    r1605 = 1'b0; 
    r1606 = 1'b0; 
    r1607 = 1'b0; 
    r1608 = 1'b0; 
    r1609 = 1'b0; 
    r1610 = 1'b0; 
    r1611 = 1'b0; 
    r1612 = 1'b0; 
    r1613 = 1'b0; 
    r1614 = 1'b0; 
    r1615 = 1'b0; 
    r1616 = 1'b0; 
    r1617 = 1'b0; 
    r1618 = 1'b0; 
    r1619 = 1'b0; 
    r1620 = 1'b0; 
    r1621 = 1'b0; 
    r1622 = 1'b0; 
    r1623 = 1'b0; 
    r1624 = 1'b0; 
    r1625 = 1'b0; 
    r1626 = 1'b0; 
    r1627 = 1'b0; 
    r1628 = 1'b0; 
    r1629 = 1'b0; 
    r1630 = 1'b0; 
    r1631 = 1'b0; 
    r1632 = 1'b0; 
    r1633 = 1'b0; 
    r1634 = 1'b0; 
    r1635 = 1'b0; 
    r1636 = 1'b0; 
    r1637 = 1'b0; 
    r1638 = 1'b0; 
    r1639 = 1'b0; 
    r1640 = 1'b0; 
    r1641 = 1'b0; 
    r1642 = 1'b0; 
    r1643 = 1'b0; 
    r1644 = 1'b0; 
    r1645 = 1'b0; 
    r1646 = 1'b0; 
    r1647 = 1'b0; 
    r1648 = 1'b0; 
    r1649 = 1'b0; 
    r1650 = 1'b0; 
    r1651 = 1'b0; 
    r1652 = 1'b0; 
    r1653 = 1'b0; 
    r1654 = 1'b0; 
    r1655 = 1'b0; 
    r1656 = 1'b0; 
    r1657 = 1'b0; 
    r1658 = 1'b0; 
    r1659 = 1'b0; 
    r1660 = 1'b0; 
    r1661 = 1'b0; 
    r1662 = 1'b0; 
    r1663 = 1'b0; 
    r1664 = 1'b0; 
    r1665 = 1'b0; 
    r1666 = 1'b0; 
    r1667 = 1'b0; 
    r1668 = 1'b0; 
    r1669 = 1'b0; 
    r1670 = 1'b0; 
    r1671 = 1'b0; 
    r1672 = 1'b0; 
    r1673 = 1'b0; 
    r1674 = 1'b0; 
    r1675 = 1'b0; 
    r1676 = 1'b0; 
    r1677 = 1'b0; 
    r1678 = 1'b0; 
    r1679 = 1'b0; 
    r1680 = 1'b0; 
    r1681 = 1'b0; 
    r1682 = 1'b0; 
    r1683 = 1'b0; 
    r1684 = 1'b0; 
    r1685 = 1'b0; 
    r1686 = 1'b0; 
    r1687 = 1'b0; 
    r1688 = 1'b0; 
    r1689 = 1'b0; 
    r1690 = 1'b0; 
    r1691 = 1'b0; 
    r1692 = 1'b0; 
    r1693 = 1'b0; 
    r1694 = 1'b0; 
    r1695 = 1'b0; 
    r1696 = 1'b0; 
    r1697 = 1'b0; 
    r1698 = 1'b0; 
    r1699 = 1'b0; 
    r1700 = 1'b0; 
    r1701 = 1'b0; 
    r1702 = 1'b0; 
    r1703 = 1'b0; 
    r1704 = 1'b0; 
    r1705 = 1'b0; 
    r1706 = 1'b0; 
    r1707 = 1'b0; 
    r1708 = 1'b0; 
    r1709 = 1'b0; 
    r1710 = 1'b0; 
    r1711 = 1'b0; 
    r1712 = 1'b0; 
    r1713 = 1'b0; 
    r1714 = 1'b0; 
    r1715 = 1'b0; 
    r1716 = 1'b0; 
    r1717 = 1'b0; 
    r1718 = 1'b0; 
    r1719 = 1'b0; 
    r1720 = 1'b0; 
    r1721 = 1'b0; 
    r1722 = 1'b0; 
    r1723 = 1'b0; 
    r1724 = 1'b0; 
    r1725 = 1'b0; 
    r1726 = 1'b0; 
    r1727 = 1'b0; 
    r1728 = 1'b0; 
    r1729 = 1'b0; 
    r1730 = 1'b0; 
    r1731 = 1'b0; 
    r1732 = 1'b0; 
    r1733 = 1'b0; 
    r1734 = 1'b0; 
    r1735 = 1'b0; 
    r1736 = 1'b0; 
    r1737 = 1'b0; 
    r1738 = 1'b0; 
    r1739 = 1'b0; 
    r1740 = 1'b0; 
    r1741 = 1'b0; 
    r1742 = 1'b0; 
    r1743 = 1'b0; 
    r1744 = 1'b0; 
    r1745 = 1'b0; 
    r1746 = 1'b0; 
    r1747 = 1'b0; 
    r1748 = 1'b0; 
    r1749 = 1'b0; 
    r1750 = 1'b0; 
    r1751 = 1'b0; 
    r1752 = 1'b0; 
    r1753 = 1'b0; 
    r1754 = 1'b0; 
    r1755 = 1'b0; 
    r1756 = 1'b0; 
    r1757 = 1'b0; 
    r1758 = 1'b0; 
    r1759 = 1'b0; 
    r1760 = 1'b0; 
    r1761 = 1'b0; 
    r1762 = 1'b0; 
    r1763 = 1'b0; 
    r1764 = 1'b0; 
    r1765 = 1'b0; 
    r1766 = 1'b0; 
    r1767 = 1'b0; 
    r1768 = 1'b0; 
    r1769 = 1'b0; 
    r1770 = 1'b0; 
    r1771 = 1'b0; 
    r1772 = 1'b0; 
    r1773 = 1'b0; 
    r1774 = 1'b0; 
    r1775 = 1'b0; 
    r1776 = 1'b0; 
    r1777 = 1'b0; 
    r1778 = 1'b0; 
    r1779 = 1'b0; 
    r1780 = 1'b0; 
    r1781 = 1'b0; 
    r1782 = 1'b0; 
    r1783 = 1'b0; 
    r1784 = 1'b0; 
    r1785 = 1'b0; 
    r1786 = 1'b0; 
    r1787 = 1'b0; 
    r1788 = 1'b0; 
    r1789 = 1'b0; 
    r1790 = 1'b0; 
    r1791 = 1'b0; 
    r1792 = 1'b0; 
    r1793 = 1'b0; 
    r1794 = 1'b0; 
    r1795 = 1'b0; 
    r1796 = 1'b0; 
    r1797 = 1'b0; 
    r1798 = 1'b0; 
    r1799 = 1'b0; 
    r1800 = 1'b0; 
    r1801 = 1'b0; 
    r1802 = 1'b0; 
    r1803 = 1'b0; 
    r1804 = 1'b0; 
    r1805 = 1'b0; 
    r1806 = 1'b0; 
    r1807 = 1'b0; 
    r1808 = 1'b0; 
    r1809 = 1'b0; 
    r1810 = 1'b0; 
    r1811 = 1'b0; 
    r1812 = 1'b0; 
    r1813 = 1'b0; 
    r1814 = 1'b0; 
    r1815 = 1'b0; 
    r1816 = 1'b0; 
    r1817 = 1'b0; 
    r1818 = 1'b0; 
    r1819 = 1'b0; 
    r1820 = 1'b0; 
    r1821 = 1'b0; 
    r1822 = 1'b0; 
    r1823 = 1'b0; 
    r1824 = 1'b0; 
    r1825 = 1'b0; 
    r1826 = 1'b0; 
    r1827 = 1'b0; 
    r1828 = 1'b0; 
    r1829 = 1'b0; 
    r1830 = 1'b0; 
    r1831 = 1'b0; 
    r1832 = 1'b0; 
    r1833 = 1'b0; 
    r1834 = 1'b0; 
    r1835 = 1'b0; 
    r1836 = 1'b0; 
    r1837 = 1'b0; 
    r1838 = 1'b0; 
    r1839 = 1'b0; 
    r1840 = 1'b0; 
    r1841 = 1'b0; 
    r1842 = 1'b0; 
    r1843 = 1'b0; 
    r1844 = 1'b0; 
    r1845 = 1'b0; 
    r1846 = 1'b0; 
    r1847 = 1'b0; 
    r1848 = 1'b0; 
    r1849 = 1'b0; 
    r1850 = 1'b0; 
    r1851 = 1'b0; 
    r1852 = 1'b0; 
    r1853 = 1'b0; 
    r1854 = 1'b0; 
    r1855 = 1'b0; 
    r1856 = 1'b0; 
    r1857 = 1'b0; 
    r1858 = 1'b0; 
    r1859 = 1'b0; 
    r1860 = 1'b0; 
    r1861 = 1'b0; 
    r1862 = 1'b0; 
    r1863 = 1'b0; 
    r1864 = 1'b0; 
    r1865 = 1'b0; 
    r1866 = 1'b0; 
    r1867 = 1'b0; 
    r1868 = 1'b0; 
    r1869 = 1'b0; 
    r1870 = 1'b0; 
    r1871 = 1'b0; 
    r1872 = 1'b0; 
    r1873 = 1'b0; 
    r1874 = 1'b0; 
    r1875 = 1'b0; 
    r1876 = 1'b0; 
    r1877 = 1'b0; 
    r1878 = 1'b0; 
    r1879 = 1'b0; 
    r1880 = 1'b0; 
    r1881 = 1'b0; 
    r1882 = 1'b0; 
    r1883 = 1'b0; 
    r1884 = 1'b0; 
    r1885 = 1'b0; 
    r1886 = 1'b0; 
    r1887 = 1'b0; 
    r1888 = 1'b0; 
    r1889 = 1'b0; 
    r1890 = 1'b0; 
    r1891 = 1'b0; 
    r1892 = 1'b0; 
    r1893 = 1'b0; 
    r1894 = 1'b0; 
    r1895 = 1'b0; 
    r1896 = 1'b0; 
    r1897 = 1'b0; 
    r1898 = 1'b0; 
    r1899 = 1'b0; 
    r1900 = 1'b0; 
    r1901 = 1'b0; 
    r1902 = 1'b0; 
    r1903 = 1'b0; 
    r1904 = 1'b0; 
    r1905 = 1'b0; 
    r1906 = 1'b0; 
    r1907 = 1'b0; 
    r1908 = 1'b0; 
    r1909 = 1'b0; 
    r1910 = 1'b0; 
    r1911 = 1'b0; 
    r1912 = 1'b0; 
    r1913 = 1'b0; 
    r1914 = 1'b0; 
    r1915 = 1'b0; 
    r1916 = 1'b0; 
    r1917 = 1'b0; 
    r1918 = 1'b0; 
    r1919 = 1'b0; 
    r1920 = 1'b0; 
    r1921 = 1'b0; 
    r1922 = 1'b0; 
    r1923 = 1'b0; 
    r1924 = 1'b0; 
    r1925 = 1'b0; 
    r1926 = 1'b0; 
    r1927 = 1'b0; 
    r1928 = 1'b0; 
    r1929 = 1'b0; 
    r1930 = 1'b0; 
    r1931 = 1'b0; 
    r1932 = 1'b0; 
    r1933 = 1'b0; 
    r1934 = 1'b0; 
    r1935 = 1'b0; 
    r1936 = 1'b0; 
    r1937 = 1'b0; 
    r1938 = 1'b0; 
    r1939 = 1'b0; 
    r1940 = 1'b0; 
    r1941 = 1'b0; 
    r1942 = 1'b0; 
    r1943 = 1'b0; 
    r1944 = 1'b0; 
    r1945 = 1'b0; 
    r1946 = 1'b0; 
    r1947 = 1'b0; 
    r1948 = 1'b0; 
    r1949 = 1'b0; 
    r1950 = 1'b0; 
    r1951 = 1'b0; 
    r1952 = 1'b0; 
    r1953 = 1'b0; 
    r1954 = 1'b0; 
    r1955 = 1'b0; 
    r1956 = 1'b0; 
    r1957 = 1'b0; 
    r1958 = 1'b0; 
    r1959 = 1'b0; 
    r1960 = 1'b0; 
    r1961 = 1'b0; 
    r1962 = 1'b0; 
    r1963 = 1'b0; 
    r1964 = 1'b0; 
    r1965 = 1'b0; 
    r1966 = 1'b0; 
    r1967 = 1'b0; 
    r1968 = 1'b0; 
    r1969 = 1'b0; 
    r1970 = 1'b0; 
    r1971 = 1'b0; 
    r1972 = 1'b0; 
    r1973 = 1'b0; 
    r1974 = 1'b0; 
    r1975 = 1'b0; 
    r1976 = 1'b0; 
    r1977 = 1'b0; 
    r1978 = 1'b0; 
    r1979 = 1'b0; 
    r1980 = 1'b0; 
    r1981 = 1'b0; 
    r1982 = 1'b0; 
    r1983 = 1'b0; 
    r1984 = 1'b0; 
    r1985 = 1'b0; 
    r1986 = 1'b0; 
    r1987 = 1'b0; 
    r1988 = 1'b0; 
    r1989 = 1'b0; 
    r1990 = 1'b0; 
    r1991 = 1'b0; 
    r1992 = 1'b0; 
    r1993 = 1'b0; 
    r1994 = 1'b0; 
    r1995 = 1'b0; 
    r1996 = 1'b0; 
    r1997 = 1'b0; 
    $monitor("%t %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b  ", $time, w_000_000, w_000_001, w_000_002, w_000_003, w_000_004, w_000_005, w_000_006, w_000_007, w_000_008, w_000_009, w_000_010, w_000_011, w_000_012, w_000_013, w_000_014, w_000_015, w_000_016, w_000_017, w_000_018, w_000_019, w_000_020, w_000_021, w_000_022, w_000_023, w_000_024, w_000_025, w_000_026, w_000_027, w_000_028, w_000_029, w_000_030, w_000_031, w_000_032, w_000_033, w_000_034, w_000_035, w_000_036, w_000_037, w_000_038, w_000_039, w_000_040, w_000_041, w_000_042, w_000_043, w_000_044, w_000_045, w_000_046, w_000_047, w_000_048, w_000_049, w_000_050, w_000_051, w_000_052, w_000_053, w_000_054, w_000_055, w_000_056, w_000_057, w_000_058, w_000_059, w_000_060, w_000_061, w_000_062, w_000_063, w_000_064, w_000_065, w_000_066, w_000_067, w_000_068, w_000_069, w_000_070, w_000_071, w_000_072, w_000_073, w_000_074, w_000_075, w_000_076, w_000_077, w_000_078, w_000_079, w_000_080, w_000_081, w_000_082, w_000_083, w_000_084, w_000_085, w_000_086, w_000_087, w_000_088, w_000_089, w_000_090, w_000_091, w_000_092, w_000_093, w_000_094, w_000_095, w_000_096, w_000_097, w_000_098, w_000_099, w_000_100, w_000_101, w_000_102, w_000_103, w_000_104, w_000_105, w_000_106, w_000_107, w_000_108, w_000_109, w_000_110, w_000_111, w_000_112, w_000_113, w_000_114, w_000_115, w_000_116, w_000_117, w_000_118, w_000_119, w_000_120, w_000_121, w_000_122, w_000_123, w_000_124, w_000_125, w_000_126, w_000_127, w_000_128, w_000_129, w_000_130, w_000_131, w_000_132, w_000_133, w_000_134, w_000_135, w_000_136, w_000_137, w_000_138, w_000_139, w_000_140, w_000_141, w_000_142, w_000_143, w_000_144, w_000_145, w_000_146, w_000_147, w_000_148, w_000_149, w_000_150, w_000_151, w_000_152, w_000_153, w_000_154, w_000_155, w_000_156, w_000_157, w_000_158, w_000_159, w_000_160, w_000_161, w_000_162, w_000_163, w_000_164, w_000_165, w_000_166, w_000_167, w_000_168, w_000_169, w_000_170, w_000_171, w_000_172, w_000_173, w_000_174, w_000_175, w_000_176, w_000_177, w_000_178, w_000_179, w_000_180, w_000_181, w_000_182, w_000_183, w_000_184, w_000_185, w_000_186, w_000_187, w_000_188, w_000_189, w_000_190, w_000_191, w_000_192, w_000_193, w_000_194, w_000_195, w_000_196, w_000_197, w_000_198, w_000_199, w_000_200, w_000_201, w_000_202, w_000_203, w_000_204, w_000_205, w_000_206, w_000_207, w_000_208, w_000_209, w_000_210, w_000_211, w_000_212, w_000_213, w_000_214, w_000_215, w_000_216, w_000_217, w_000_218, w_000_219, w_000_220, w_000_221, w_000_222, w_000_223, w_000_224, w_000_225, w_000_226, w_000_227, w_000_228, w_000_229, w_000_230, w_000_231, w_000_232, w_000_233, w_000_234, w_000_235, w_000_236, w_000_237, w_000_238, w_000_239, w_000_240, w_000_241, w_000_242, w_000_243, w_000_244, w_000_245, w_000_246, w_000_247, w_000_248, w_000_249, w_000_250, w_000_251, w_000_252, w_000_253, w_000_254, w_000_255, w_000_256, w_000_257, w_000_258, w_000_259, w_000_260, w_000_261, w_000_262, w_000_263, w_000_264, w_000_265, w_000_266, w_000_267, w_000_268, w_000_269, w_000_270, w_000_271, w_000_272, w_000_273, w_000_274, w_000_275, w_000_276, w_000_277, w_000_278, w_000_279, w_000_280, w_000_281, w_000_282, w_000_283, w_000_284, w_000_285, w_000_286, w_000_287, w_000_288, w_000_289, w_000_290, w_000_291, w_000_292, w_000_293, w_000_294, w_000_295, w_000_296, w_000_297, w_000_298, w_000_299, w_000_300, w_000_301, w_000_302, w_000_303, w_000_304, w_000_305, w_000_306, w_000_307, w_000_308, w_000_309, w_000_310, w_000_311, w_000_312, w_000_313, w_000_314, w_000_315, w_000_316, w_000_317, w_000_318, w_000_319, w_000_320, w_000_321, w_000_322, w_000_323, w_000_324, w_000_325, w_000_326, w_000_327, w_000_328, w_000_329, w_000_330, w_000_331, w_000_332, w_000_333, w_000_334, w_000_335, w_000_336, w_000_337, w_000_338, w_000_339, w_000_340, w_000_341, w_000_342, w_000_343, w_000_344, w_000_345, w_000_346, w_000_347, w_000_348, w_000_349, w_000_350, w_000_351, w_000_352, w_000_353, w_000_354, w_000_355, w_000_356, w_000_357, w_000_358, w_000_359, w_000_360, w_000_361, w_000_362, w_000_363, w_000_364, w_000_365, w_000_366, w_000_367, w_000_368, w_000_369, w_000_370, w_000_371, w_000_372, w_000_373, w_000_374, w_000_375, w_000_376, w_000_377, w_000_378, w_000_379, w_000_380, w_000_381, w_000_382, w_000_383, w_000_384, w_000_385, w_000_386, w_000_387, w_000_388, w_000_389, w_000_390, w_000_391, w_000_392, w_000_393, w_000_394, w_000_395, w_000_396, w_000_397, w_000_398, w_000_399, w_000_400, w_000_401, w_000_402, w_000_403, w_000_404, w_000_405, w_000_406, w_000_407, w_000_408, w_000_409, w_000_410, w_000_411, w_000_412, w_000_413, w_000_414, w_000_415, w_000_416, w_000_417, w_000_418, w_000_419, w_000_420, w_000_421, w_000_422, w_000_423, w_000_424, w_000_425, w_000_426, w_000_427, w_000_428, w_000_429, w_000_430, w_000_431, w_000_432, w_000_433, w_000_434, w_000_435, w_000_436, w_000_437, w_000_438, w_000_439, w_000_440, w_000_441, w_000_442, w_000_443, w_000_444, w_000_445, w_000_446, w_000_447, w_000_448, w_000_449, w_000_450, w_000_451, w_000_452, w_000_453, w_000_454, w_000_455, w_000_456, w_000_457, w_000_458, w_000_459, w_000_460, w_000_461, w_000_462, w_000_463, w_000_464, w_000_465, w_000_466, w_000_467, w_000_468, w_000_469, w_000_470, w_000_471, w_000_472, w_000_473, w_000_474, w_000_475, w_000_476, w_000_477, w_000_478, w_000_479, w_000_480, w_000_481, w_000_482, w_000_483, w_000_484, w_000_485, w_000_486, w_000_487, w_000_488, w_000_489, w_000_490, w_000_491, w_000_492, w_000_493, w_000_494, w_000_495, w_000_496, w_000_497, w_000_498, w_000_499, w_000_500, w_000_501, w_000_502, w_000_503, w_000_504, w_000_505, w_000_506, w_000_507, w_000_508, w_000_509, w_000_510, w_000_511, w_000_512, w_000_513, w_000_514, w_000_515, w_000_516, w_000_517, w_000_518, w_000_519, w_000_520, w_000_521, w_000_522, w_000_523, w_000_524, w_000_525, w_000_526, w_000_527, w_000_528, w_000_529, w_000_530, w_000_531, w_000_532, w_000_533, w_000_534, w_000_535, w_000_536, w_000_537, w_000_538, w_000_539, w_000_540, w_000_541, w_000_542, w_000_543, w_000_544, w_000_545, w_000_546, w_000_547, w_000_548, w_000_549, w_000_550, w_000_551, w_000_552, w_000_553, w_000_554, w_000_555, w_000_556, w_000_557, w_000_558, w_000_559, w_000_560, w_000_561, w_000_562, w_000_563, w_000_564, w_000_565, w_000_566, w_000_567, w_000_568, w_000_569, w_000_570, w_000_571, w_000_572, w_000_573, w_000_574, w_000_575, w_000_576, w_000_577, w_000_578, w_000_579, w_000_580, w_000_581, w_000_582, w_000_583, w_000_584, w_000_585, w_000_586, w_000_587, w_000_588, w_000_589, w_000_590, w_000_591, w_000_592, w_000_593, w_000_594, w_000_595, w_000_596, w_000_597, w_000_598, w_000_599, w_000_600, w_000_601, w_000_602, w_000_603, w_000_604, w_000_605, w_000_606, w_000_607, w_000_608, w_000_609, w_000_610, w_000_611, w_000_612, w_000_613, w_000_614, w_000_615, w_000_616, w_000_617, w_000_618, w_000_619, w_000_620, w_000_621, w_000_622, w_000_623, w_000_624, w_000_625, w_000_626, w_000_627, w_000_628, w_000_629, w_000_630, w_000_631, w_000_632, w_000_633, w_000_634, w_000_635, w_000_636, w_000_637, w_000_638, w_000_639, w_000_640, w_000_641, w_000_642, w_000_643, w_000_644, w_000_645, w_000_646, w_000_647, w_000_648, w_000_649, w_000_650, w_000_651, w_000_652, w_000_653, w_000_654, w_000_655, w_000_656, w_000_657, w_000_658, w_000_659, w_000_660, w_000_661, w_000_662, w_000_663, w_000_664, w_000_665, w_000_666, w_000_667, w_000_668, w_000_669, w_000_670, w_000_671, w_000_672, w_000_673, w_000_674, w_000_675, w_000_676, w_000_677, w_000_678, w_000_679, w_000_680, w_000_681, w_000_682, w_000_683, w_000_684, w_000_685, w_000_686, w_000_687, w_000_688, w_000_689, w_000_690, w_000_691, w_000_692, w_000_693, w_000_694, w_000_695, w_000_696, w_000_697, w_000_698, w_000_699, w_000_700, w_000_701, w_000_702, w_000_703, w_000_704, w_000_705, w_000_706, w_000_707, w_000_708, w_000_709, w_000_710, w_000_711, w_000_712, w_000_713, w_000_714, w_000_715, w_000_716, w_000_717, w_000_718, w_000_719, w_000_720, w_000_721, w_000_722, w_000_723, w_000_724, w_000_725, w_000_726, w_000_727, w_000_728, w_000_729, w_000_730, w_000_731, w_000_732, w_000_733, w_000_734, w_000_735, w_000_736, w_000_737, w_000_738, w_000_739, w_000_740, w_000_741, w_000_742, w_000_743, w_000_744, w_000_745, w_000_746, w_000_747, w_000_748, w_000_749, w_000_750, w_000_751, w_000_752, w_000_753, w_000_754, w_000_755, w_000_756, w_000_757, w_000_758, w_000_759, w_000_760, w_000_761, w_000_762, w_000_763, w_000_764, w_000_765, w_000_766, w_000_767, w_000_768, w_000_769, w_000_770, w_000_771, w_000_772, w_000_773, w_000_774, w_000_775, w_000_776, w_000_777, w_000_778, w_000_779, w_000_780, w_000_781, w_000_782, w_000_783, w_000_784, w_000_785, w_000_786, w_000_787, w_000_788, w_000_789, w_000_790, w_000_791, w_000_792, w_000_793, w_000_794, w_000_795, w_000_796, w_000_797, w_000_798, w_000_799, w_000_800, w_000_801, w_000_802, w_000_803, w_000_804, w_000_805, w_000_806, w_000_807, w_000_808, w_000_809, w_000_810, w_000_811, w_000_812, w_000_813, w_000_814, w_000_815, w_000_816, w_000_817, w_000_818, w_000_819, w_000_820, w_000_821, w_000_822, w_000_823, w_000_824, w_000_825, w_000_826, w_000_827, w_000_828, w_000_829, w_000_830, w_000_831, w_000_832, w_000_833, w_000_834, w_000_835, w_000_836, w_000_837, w_000_838, w_000_839, w_000_840, w_000_841, w_000_842, w_000_843, w_000_844, w_000_845, w_000_846, w_000_847, w_000_848, w_000_849, w_000_850, w_000_851, w_000_852, w_000_853, w_000_854, w_000_855, w_000_856, w_000_857, w_000_858, w_000_859, w_000_860, w_000_861, w_000_862, w_000_863, w_000_864, w_000_865, w_000_866, w_000_867, w_000_868, w_000_869, w_000_870, w_000_871, w_000_872, w_000_873, w_000_874, w_000_875, w_000_876, w_000_877, w_000_878, w_000_879, w_000_880, w_000_881, w_000_882, w_000_883, w_000_884, w_000_885, w_000_886, w_000_887, w_000_888, w_000_889, w_000_890, w_000_891, w_000_892, w_000_893, w_000_894, w_000_895, w_000_896, w_000_897, w_000_898, w_000_899, w_000_900, w_000_901, w_000_902, w_000_903, w_000_904, w_000_905, w_000_906, w_000_907, w_000_908, w_000_909, w_000_910, w_000_911, w_000_912, w_000_913, w_000_914, w_000_915, w_000_916, w_000_917, w_000_918, w_000_919, w_000_920, w_000_921, w_000_922, w_000_923, w_000_924, w_000_925, w_000_926, w_000_927, w_000_928, w_000_929, w_000_930, w_000_931, w_000_932, w_000_933, w_000_934, w_000_935, w_000_936, w_000_937, w_000_938, w_000_939, w_000_940, w_000_941, w_000_942, w_000_943, w_000_944, w_000_945, w_000_946, w_000_947, w_000_948, w_000_949, w_000_950, w_000_951, w_000_952, w_000_953, w_000_954, w_000_955, w_000_956, w_000_957, w_000_958, w_000_959, w_000_960, w_000_961, w_000_962, w_000_963, w_000_964, w_000_965, w_000_966, w_000_967, w_000_968, w_000_969, w_000_970, w_000_971, w_000_972, w_000_973, w_000_974, w_000_975, w_000_976, w_000_977, w_000_978, w_000_979, w_000_980, w_000_981, w_000_982, w_000_983, w_000_984, w_000_985, w_000_986, w_000_987, w_000_988, w_000_989, w_000_990, w_000_991, w_000_992, w_000_993, w_000_994, w_000_995, w_000_996, w_000_997, w_000_998, w_000_999, w_000_1000, w_000_1001, w_000_1002, w_000_1003, w_000_1004, w_000_1005, w_000_1006, w_000_1007, w_000_1008, w_000_1009, w_000_1010, w_000_1011, w_000_1012, w_000_1013, w_000_1014, w_000_1015, w_000_1016, w_000_1017, w_000_1018, w_000_1019, w_000_1020, w_000_1021, w_000_1022, w_000_1023, w_000_1024, w_000_1025, w_000_1026, w_000_1027, w_000_1028, w_000_1029, w_000_1030, w_000_1031, w_000_1032, w_000_1033, w_000_1034, w_000_1035, w_000_1036, w_000_1037, w_000_1038, w_000_1039, w_000_1040, w_000_1041, w_000_1042, w_000_1043, w_000_1044, w_000_1045, w_000_1046, w_000_1047, w_000_1048, w_000_1049, w_000_1050, w_000_1051, w_000_1052, w_000_1053, w_000_1054, w_000_1055, w_000_1056, w_000_1057, w_000_1058, w_000_1059, w_000_1060, w_000_1061, w_000_1062, w_000_1063, w_000_1064, w_000_1065, w_000_1066, w_000_1067, w_000_1068, w_000_1069, w_000_1070, w_000_1071, w_000_1072, w_000_1073, w_000_1074, w_000_1075, w_000_1076, w_000_1077, w_000_1078, w_000_1079, w_000_1080, w_000_1081, w_000_1082, w_000_1083, w_000_1084, w_000_1085, w_000_1086, w_000_1087, w_000_1088, w_000_1089, w_000_1090, w_000_1091, w_000_1092, w_000_1093, w_000_1094, w_000_1095, w_000_1096, w_000_1097, w_000_1098, w_000_1099, w_000_1100, w_000_1101, w_000_1102, w_000_1103, w_000_1104, w_000_1105, w_000_1106, w_000_1107, w_000_1108, w_000_1109, w_000_1110, w_000_1111, w_000_1112, w_000_1113, w_000_1114, w_000_1115, w_000_1116, w_000_1117, w_000_1118, w_000_1119, w_000_1120, w_000_1121, w_000_1122, w_000_1123, w_000_1124, w_000_1125, w_000_1126, w_000_1127, w_000_1128, w_000_1129, w_000_1130, w_000_1131, w_000_1132, w_000_1133, w_000_1134, w_000_1135, w_000_1136, w_000_1137, w_000_1138, w_000_1139, w_000_1140, w_000_1141, w_000_1142, w_000_1143, w_000_1144, w_000_1145, w_000_1146, w_000_1147, w_000_1148, w_000_1149, w_000_1150, w_000_1151, w_000_1152, w_000_1153, w_000_1154, w_000_1155, w_000_1156, w_000_1157, w_000_1158, w_000_1159, w_000_1160, w_000_1161, w_000_1162, w_000_1163, w_000_1164, w_000_1165, w_000_1166, w_000_1167, w_000_1168, w_000_1169, w_000_1170, w_000_1171, w_000_1172, w_000_1173, w_000_1174, w_000_1175, w_000_1176, w_000_1177, w_000_1178, w_000_1179, w_000_1180, w_000_1181, w_000_1182, w_000_1183, w_000_1184, w_000_1185, w_000_1186, w_000_1187, w_000_1188, w_000_1189, w_000_1190, w_000_1191, w_000_1192, w_000_1193, w_000_1194, w_000_1195, w_000_1196, w_000_1197, w_000_1198, w_000_1199, w_000_1200, w_000_1201, w_000_1202, w_000_1203, w_000_1204, w_000_1205, w_000_1206, w_000_1207, w_000_1208, w_000_1209, w_000_1210, w_000_1211, w_000_1212, w_000_1213, w_000_1214, w_000_1215, w_000_1216, w_000_1217, w_000_1218, w_000_1219, w_000_1220, w_000_1221, w_000_1222, w_000_1223, w_000_1224, w_000_1225, w_000_1226, w_000_1227, w_000_1228, w_000_1229, w_000_1230, w_000_1231, w_000_1232, w_000_1233, w_000_1234, w_000_1235, w_000_1236, w_000_1237, w_000_1238, w_000_1239, w_000_1240, w_000_1241, w_000_1242, w_000_1243, w_000_1244, w_000_1245, w_000_1246, w_000_1247, w_000_1248, w_000_1249, w_000_1250, w_000_1251, w_000_1252, w_000_1253, w_000_1254, w_000_1255, w_000_1256, w_000_1257, w_000_1258, w_000_1259, w_000_1260, w_000_1261, w_000_1262, w_000_1263, w_000_1264, w_000_1265, w_000_1266, w_000_1267, w_000_1268, w_000_1269, w_000_1270, w_000_1271, w_000_1272, w_000_1273, w_000_1274, w_000_1275, w_000_1276, w_000_1277, w_000_1278, w_000_1279, w_000_1280, w_000_1281, w_000_1282, w_000_1283, w_000_1284, w_000_1285, w_000_1286, w_000_1287, w_000_1288, w_000_1289, w_000_1290, w_000_1291, w_000_1292, w_000_1293, w_000_1294, w_000_1295, w_000_1296, w_000_1297, w_000_1298, w_000_1299, w_000_1300, w_000_1301, w_000_1302, w_000_1303, w_000_1304, w_000_1305, w_000_1306, w_000_1307, w_000_1308, w_000_1309, w_000_1310, w_000_1311, w_000_1312, w_000_1313, w_000_1314, w_000_1315, w_000_1316, w_000_1317, w_000_1318, w_000_1319, w_000_1320, w_000_1321, w_000_1322, w_000_1323, w_000_1324, w_000_1325, w_000_1326, w_000_1327, w_000_1328, w_000_1329, w_000_1330, w_000_1331, w_000_1332, w_000_1333, w_000_1334, w_000_1335, w_000_1336, w_000_1337, w_000_1338, w_000_1339, w_000_1340, w_000_1341, w_000_1342, w_000_1343, w_000_1344, w_000_1345, w_000_1346, w_000_1347, w_000_1348, w_000_1349, w_000_1350, w_000_1351, w_000_1352, w_000_1353, w_000_1354, w_000_1355, w_000_1356, w_000_1357, w_000_1358, w_000_1359, w_000_1360, w_000_1361, w_000_1362, w_000_1363, w_000_1364, w_000_1365, w_000_1366, w_000_1367, w_000_1368, w_000_1369, w_000_1370, w_000_1371, w_000_1372, w_000_1373, w_000_1374, w_000_1375, w_000_1376, w_000_1377, w_000_1378, w_000_1379, w_000_1380, w_000_1381, w_000_1382, w_000_1383, w_000_1384, w_000_1385, w_000_1386, w_000_1387, w_000_1388, w_000_1389, w_000_1390, w_000_1391, w_000_1392, w_000_1393, w_000_1394, w_000_1395, w_000_1396, w_000_1397, w_000_1398, w_000_1399, w_000_1400, w_000_1401, w_000_1402, w_000_1403, w_000_1404, w_000_1405, w_000_1406, w_000_1407, w_000_1408, w_000_1409, w_000_1410, w_000_1411, w_000_1412, w_000_1413, w_000_1414, w_000_1415, w_000_1416, w_000_1417, w_000_1418, w_000_1419, w_000_1420, w_000_1421, w_000_1422, w_000_1423, w_000_1424, w_000_1425, w_000_1426, w_000_1427, w_000_1428, w_000_1429, w_000_1430, w_000_1431, w_000_1432, w_000_1433, w_000_1434, w_000_1435, w_000_1436, w_000_1437, w_000_1438, w_000_1439, w_000_1440, w_000_1441, w_000_1442, w_000_1443, w_000_1444, w_000_1445, w_000_1446, w_000_1447, w_000_1448, w_000_1449, w_000_1450, w_000_1451, w_000_1452, w_000_1453, w_000_1454, w_000_1455, w_000_1456, w_000_1457, w_000_1458, w_000_1459, w_000_1460, w_000_1461, w_000_1462, w_000_1463, w_000_1464, w_000_1465, w_000_1466, w_000_1467, w_000_1468, w_000_1469, w_000_1470, w_000_1471, w_000_1472, w_000_1473, w_000_1474, w_000_1475, w_000_1476, w_000_1477, w_000_1478, w_000_1479, w_000_1480, w_000_1481, w_000_1482, w_000_1483, w_000_1484, w_000_1485, w_000_1486, w_000_1487, w_000_1488, w_000_1489, w_000_1490, w_000_1491, w_000_1492, w_000_1493, w_000_1494, w_000_1495, w_000_1496, w_000_1497, w_000_1498, w_000_1499, w_000_1500, w_000_1501, w_000_1502, w_000_1503, w_000_1504, w_000_1505, w_000_1506, w_000_1507, w_000_1508, w_000_1509, w_000_1510, w_000_1511, w_000_1512, w_000_1513, w_000_1514, w_000_1515, w_000_1516, w_000_1517, w_000_1518, w_000_1519, w_000_1520, w_000_1521, w_000_1522, w_000_1523, w_000_1524, w_000_1525, w_000_1526, w_000_1527, w_000_1528, w_000_1529, w_000_1530, w_000_1531, w_000_1532, w_000_1533, w_000_1534, w_000_1535, w_000_1536, w_000_1537, w_000_1538, w_000_1539, w_000_1540, w_000_1541, w_000_1542, w_000_1543, w_000_1544, w_000_1545, w_000_1546, w_000_1547, w_000_1548, w_000_1549, w_000_1550, w_000_1551, w_000_1552, w_000_1553, w_000_1554, w_000_1555, w_000_1556, w_000_1557, w_000_1558, w_000_1559, w_000_1560, w_000_1561, w_000_1562, w_000_1563, w_000_1564, w_000_1565, w_000_1566, w_000_1567, w_000_1568, w_000_1569, w_000_1570, w_000_1571, w_000_1572, w_000_1573, w_000_1574, w_000_1575, w_000_1576, w_000_1577, w_000_1578, w_000_1579, w_000_1580, w_000_1581, w_000_1582, w_000_1583, w_000_1584, w_000_1585, w_000_1586, w_000_1587, w_000_1588, w_000_1589, w_000_1590, w_000_1591, w_000_1592, w_000_1593, w_000_1594, w_000_1595, w_000_1596, w_000_1597, w_000_1598, w_000_1599, w_000_1600, w_000_1601, w_000_1602, w_000_1603, w_000_1604, w_000_1605, w_000_1606, w_000_1607, w_000_1608, w_000_1609, w_000_1610, w_000_1611, w_000_1612, w_000_1613, w_000_1614, w_000_1615, w_000_1616, w_000_1617, w_000_1618, w_000_1619, w_000_1620, w_000_1621, w_000_1622, w_000_1623, w_000_1624, w_000_1625, w_000_1626, w_000_1627, w_000_1628, w_000_1629, w_000_1630, w_000_1631, w_000_1632, w_000_1633, w_000_1634, w_000_1635, w_000_1636, w_000_1637, w_000_1638, w_000_1639, w_000_1640, w_000_1641, w_000_1642, w_000_1643, w_000_1644, w_000_1645, w_000_1646, w_000_1647, w_000_1648, w_000_1649, w_000_1650, w_000_1651, w_000_1652, w_000_1653, w_000_1654, w_000_1655, w_000_1656, w_000_1657, w_000_1658, w_000_1659, w_000_1660, w_000_1661, w_000_1662, w_000_1663, w_000_1664, w_000_1665, w_000_1666, w_000_1667, w_000_1668, w_000_1669, w_000_1670, w_000_1671, w_000_1672, w_000_1673, w_000_1674, w_000_1675, w_000_1676, w_000_1677, w_000_1678, w_000_1679, w_000_1680, w_000_1681, w_000_1682, w_000_1683, w_000_1684, w_000_1685, w_000_1686, w_000_1687, w_000_1688, w_000_1689, w_000_1690, w_000_1691, w_000_1692, w_000_1693, w_000_1694, w_000_1695, w_000_1696, w_000_1697, w_000_1698, w_000_1699, w_000_1700, w_000_1701, w_000_1702, w_000_1703, w_000_1704, w_000_1705, w_000_1706, w_000_1707, w_000_1708, w_000_1709, w_000_1710, w_000_1711, w_000_1712, w_000_1713, w_000_1714, w_000_1715, w_000_1716, w_000_1717, w_000_1718, w_000_1719, w_000_1720, w_000_1721, w_000_1722, w_000_1723, w_000_1724, w_000_1725, w_000_1726, w_000_1727, w_000_1728, w_000_1729, w_000_1730, w_000_1731, w_000_1732, w_000_1733, w_000_1734, w_000_1735, w_000_1736, w_000_1737, w_000_1738, w_000_1739, w_000_1740, w_000_1741, w_000_1742, w_000_1743, w_000_1744, w_000_1745, w_000_1746, w_000_1747, w_000_1748, w_000_1749, w_000_1750, w_000_1751, w_000_1752, w_000_1753, w_000_1754, w_000_1755, w_000_1756, w_000_1757, w_000_1758, w_000_1759, w_000_1760, w_000_1761, w_000_1762, w_000_1763, w_000_1764, w_000_1765, w_000_1766, w_000_1767, w_000_1768, w_000_1769, w_000_1770, w_000_1771, w_000_1772, w_000_1773, w_000_1774, w_000_1775, w_000_1776, w_000_1777, w_000_1778, w_000_1779, w_000_1780, w_000_1781, w_000_1782, w_000_1783, w_000_1784, w_000_1785, w_000_1786, w_000_1787, w_000_1788, w_000_1789, w_000_1790, w_000_1791, w_000_1792, w_000_1793, w_000_1794, w_000_1795, w_000_1796, w_000_1797, w_000_1798, w_000_1799, w_000_1800, w_000_1801, w_000_1802, w_000_1803, w_000_1804, w_000_1805, w_000_1806, w_000_1807, w_000_1808, w_000_1809, w_000_1810, w_000_1811, w_000_1812, w_000_1813, w_000_1814, w_000_1815, w_000_1816, w_000_1817, w_000_1818, w_000_1819, w_000_1820, w_000_1821, w_000_1822, w_000_1823, w_000_1824, w_000_1825, w_000_1826, w_000_1827, w_000_1828, w_000_1829, w_000_1830, w_000_1831, w_000_1832, w_000_1833, w_000_1834, w_000_1835, w_000_1836, w_000_1837, w_000_1838, w_000_1839, w_000_1840, w_000_1841, w_000_1842, w_000_1843, w_000_1844, w_000_1845, w_000_1846, w_000_1847, w_000_1848, w_000_1849, w_000_1850, w_000_1851, w_000_1852, w_000_1853, w_000_1854, w_000_1855, w_000_1856, w_000_1857, w_000_1858, w_000_1859, w_000_1860, w_000_1861, w_000_1862, w_000_1863, w_000_1864, w_000_1865, w_000_1866, w_000_1867, w_000_1868, w_000_1869, w_000_1870, w_000_1871, w_000_1872, w_000_1873, w_000_1874, w_000_1875, w_000_1876, w_000_1877, w_000_1878, w_000_1879, w_000_1880, w_000_1881, w_000_1882, w_000_1883, w_000_1884, w_000_1885, w_000_1886, w_000_1887, w_000_1888, w_000_1889, w_000_1890, w_000_1891, w_000_1892, w_000_1893, w_000_1894, w_000_1895, w_000_1896, w_000_1897, w_000_1898, w_000_1899, w_000_1900, w_000_1901, w_000_1902, w_000_1903, w_000_1904, w_000_1905, w_000_1906, w_000_1907, w_000_1908, w_000_1909, w_000_1910, w_000_1911, w_000_1912, w_000_1913, w_000_1914, w_000_1915, w_000_1916, w_000_1917, w_000_1918, w_000_1919, w_000_1920, w_000_1921, w_000_1922, w_000_1923, w_000_1924, w_000_1925, w_000_1926, w_000_1927, w_000_1928, w_000_1929, w_000_1930, w_000_1931, w_000_1932, w_000_1933, w_000_1934, w_000_1935, w_000_1936, w_000_1937, w_000_1938, w_000_1939, w_000_1940, w_000_1941, w_000_1942, w_000_1943, w_000_1944, w_000_1945, w_000_1946, w_000_1947, w_000_1948, w_000_1949, w_000_1950, w_000_1951, w_000_1952, w_000_1953, w_000_1954, w_000_1955, w_000_1956, w_000_1957, w_000_1958, w_000_1959, w_000_1960, w_000_1961, w_000_1962, w_000_1963, w_000_1964, w_000_1965, w_000_1966, w_000_1967, w_000_1968, w_000_1969, w_000_1970, w_000_1971, w_000_1972, w_000_1973, w_000_1974, w_000_1975, w_000_1976, w_000_1977, w_000_1978, w_000_1979, w_000_1980, w_000_1981, w_000_1982, w_000_1983, w_000_1984, w_000_1985, w_000_1986, w_000_1987, w_000_1988, w_000_1989, w_000_1990, w_000_1991, w_000_1992, w_000_1993, w_000_1994, w_000_1995, w_000_1996, w_000_1997, w_2000_000, w_2000_001, w_2000_002, w_2000_003, w_2000_004, w_2000_005, w_2000_006, w_2000_007, w_2000_008, w_2000_009, w_2000_010, w_2000_011, w_2000_012, w_2000_013, w_2000_014, w_2000_015, w_2000_016, w_2000_017, w_2000_018, w_2000_019, w_2000_020, w_2000_021, w_2000_022, w_2000_023, w_2000_024, w_2000_025, w_2000_026, w_2000_027, w_2000_028, w_2000_029, w_2000_030, w_2000_031, w_2000_032, w_2000_033, w_2000_034, w_2000_035, w_2000_036, w_2000_037, w_2000_038, w_2000_039, w_2000_040, w_2000_041, w_2000_042, w_2000_043, w_2000_044, w_2000_045, w_2000_046, w_2000_047, w_2000_048, w_2000_049, w_2000_050, w_2000_051, w_2000_052, w_2000_053, w_2000_054, w_2000_055, w_2000_056, w_2000_057, w_2000_058, w_2000_059, w_2000_060, w_2000_061, w_2000_062, w_2000_063, w_2000_064, w_2000_065, w_2000_066, w_2000_067, w_2000_068, w_2000_069, w_2000_070, w_2000_071, w_2000_072, w_2000_073, w_2000_074, w_2000_075, w_2000_076, w_2000_077, w_2000_078, w_2000_079, w_2000_080, w_2000_081, w_2000_082, w_2000_083, w_2000_084, w_2000_085, w_2000_086, w_2000_087, w_2000_088, w_2000_089, w_2000_090, w_2000_091, w_2000_092, w_2000_093, w_2000_094, w_2000_095, w_2000_096, w_2000_097, w_2000_098, w_2000_099, w_2000_100, w_2000_101, w_2000_102, w_2000_103, w_2000_104, w_2000_105, w_2000_106, w_2000_107, w_2000_108, w_2000_109, w_2000_110);
    #100;
    $finish;
  end
  always #1 r0 = ~r0;
  always #2 r1 = ~r1;
  always #4 r2 = ~r2;
  always #8 r3 = ~r3;
  always #16 r4 = ~r4;
  always #32 r5 = ~r5;
  always #64 r6 = ~r6;
  always #128 r7 = ~r7;
  always #256 r8 = ~r8;
  always #512 r9 = ~r9;
  always #1024 r10 = ~r10;
  always #2048 r11 = ~r11;
  always #4096 r12 = ~r12;
  always #8192 r13 = ~r13;
  always #16384 r14 = ~r14;
  always #32768 r15 = ~r15;
  always #65536 r16 = ~r16;
  always #131072 r17 = ~r17;
  always #262144 r18 = ~r18;
  always #524288 r19 = ~r19;
  always #1048576 r20 = ~r20;
  always #2097152 r21 = ~r21;
  always #4194304 r22 = ~r22;
  always #8388608 r23 = ~r23;
  always #16777216 r24 = ~r24;
  always #33554432 r25 = ~r25;
  always #67108864 r26 = ~r26;
  always #134217728 r27 = ~r27;
  always #268435456 r28 = ~r28;
  always #536870912 r29 = ~r29;
  always #1073741824 r30 = ~r30;
  always #2147483648 r31 = ~r31;
  always #4294967296 r32 = ~r32;
  always #8589934592 r33 = ~r33;
  always #17179869184 r34 = ~r34;
  always #34359738368 r35 = ~r35;
  always #68719476736 r36 = ~r36;
  always #137438953472 r37 = ~r37;
  always #274877906944 r38 = ~r38;
  always #549755813888 r39 = ~r39;
  always #1099511627776 r40 = ~r40;
  always #2199023255552 r41 = ~r41;
  always #4398046511104 r42 = ~r42;
  always #8796093022208 r43 = ~r43;
  always #17592186044416 r44 = ~r44;
  always #35184372088832 r45 = ~r45;
  always #70368744177664 r46 = ~r46;
  always #140737488355328 r47 = ~r47;
  always #281474976710656 r48 = ~r48;
  always #562949953421312 r49 = ~r49;
  always #1125899906842624 r50 = ~r50;
  always #2251799813685248 r51 = ~r51;
  always #4503599627370496 r52 = ~r52;
  always #9007199254740992 r53 = ~r53;
  always #18014398509481984 r54 = ~r54;
  always #36028797018963968 r55 = ~r55;
  always #72057594037927936 r56 = ~r56;
  always #144115188075855872 r57 = ~r57;
  always #288230376151711744 r58 = ~r58;
  always #576460752303423488 r59 = ~r59;
  always #1152921504606846976 r60 = ~r60;
  always #2305843009213693952 r61 = ~r61;
  always #4611686018427387904 r62 = ~r62;
  always #9223372036854775808 r63 = ~r63;
  always #1 r64 = ~r64;
  always #2 r65 = ~r65;
  always #4 r66 = ~r66;
  always #8 r67 = ~r67;
  always #16 r68 = ~r68;
  always #32 r69 = ~r69;
  always #64 r70 = ~r70;
  always #128 r71 = ~r71;
  always #256 r72 = ~r72;
  always #512 r73 = ~r73;
  always #1024 r74 = ~r74;
  always #2048 r75 = ~r75;
  always #4096 r76 = ~r76;
  always #8192 r77 = ~r77;
  always #16384 r78 = ~r78;
  always #32768 r79 = ~r79;
  always #65536 r80 = ~r80;
  always #131072 r81 = ~r81;
  always #262144 r82 = ~r82;
  always #524288 r83 = ~r83;
  always #1048576 r84 = ~r84;
  always #2097152 r85 = ~r85;
  always #4194304 r86 = ~r86;
  always #8388608 r87 = ~r87;
  always #16777216 r88 = ~r88;
  always #33554432 r89 = ~r89;
  always #67108864 r90 = ~r90;
  always #134217728 r91 = ~r91;
  always #268435456 r92 = ~r92;
  always #536870912 r93 = ~r93;
  always #1073741824 r94 = ~r94;
  always #2147483648 r95 = ~r95;
  always #4294967296 r96 = ~r96;
  always #8589934592 r97 = ~r97;
  always #17179869184 r98 = ~r98;
  always #34359738368 r99 = ~r99;
  always #68719476736 r100 = ~r100;
  always #137438953472 r101 = ~r101;
  always #274877906944 r102 = ~r102;
  always #549755813888 r103 = ~r103;
  always #1099511627776 r104 = ~r104;
  always #2199023255552 r105 = ~r105;
  always #4398046511104 r106 = ~r106;
  always #8796093022208 r107 = ~r107;
  always #17592186044416 r108 = ~r108;
  always #35184372088832 r109 = ~r109;
  always #70368744177664 r110 = ~r110;
  always #140737488355328 r111 = ~r111;
  always #281474976710656 r112 = ~r112;
  always #562949953421312 r113 = ~r113;
  always #1125899906842624 r114 = ~r114;
  always #2251799813685248 r115 = ~r115;
  always #4503599627370496 r116 = ~r116;
  always #9007199254740992 r117 = ~r117;
  always #18014398509481984 r118 = ~r118;
  always #36028797018963968 r119 = ~r119;
  always #72057594037927936 r120 = ~r120;
  always #144115188075855872 r121 = ~r121;
  always #288230376151711744 r122 = ~r122;
  always #576460752303423488 r123 = ~r123;
  always #1152921504606846976 r124 = ~r124;
  always #2305843009213693952 r125 = ~r125;
  always #4611686018427387904 r126 = ~r126;
  always #9223372036854775808 r127 = ~r127;
  always #1 r128 = ~r128;
  always #2 r129 = ~r129;
  always #4 r130 = ~r130;
  always #8 r131 = ~r131;
  always #16 r132 = ~r132;
  always #32 r133 = ~r133;
  always #64 r134 = ~r134;
  always #128 r135 = ~r135;
  always #256 r136 = ~r136;
  always #512 r137 = ~r137;
  always #1024 r138 = ~r138;
  always #2048 r139 = ~r139;
  always #4096 r140 = ~r140;
  always #8192 r141 = ~r141;
  always #16384 r142 = ~r142;
  always #32768 r143 = ~r143;
  always #65536 r144 = ~r144;
  always #131072 r145 = ~r145;
  always #262144 r146 = ~r146;
  always #524288 r147 = ~r147;
  always #1048576 r148 = ~r148;
  always #2097152 r149 = ~r149;
  always #4194304 r150 = ~r150;
  always #8388608 r151 = ~r151;
  always #16777216 r152 = ~r152;
  always #33554432 r153 = ~r153;
  always #67108864 r154 = ~r154;
  always #134217728 r155 = ~r155;
  always #268435456 r156 = ~r156;
  always #536870912 r157 = ~r157;
  always #1073741824 r158 = ~r158;
  always #2147483648 r159 = ~r159;
  always #4294967296 r160 = ~r160;
  always #8589934592 r161 = ~r161;
  always #17179869184 r162 = ~r162;
  always #34359738368 r163 = ~r163;
  always #68719476736 r164 = ~r164;
  always #137438953472 r165 = ~r165;
  always #274877906944 r166 = ~r166;
  always #549755813888 r167 = ~r167;
  always #1099511627776 r168 = ~r168;
  always #2199023255552 r169 = ~r169;
  always #4398046511104 r170 = ~r170;
  always #8796093022208 r171 = ~r171;
  always #17592186044416 r172 = ~r172;
  always #35184372088832 r173 = ~r173;
  always #70368744177664 r174 = ~r174;
  always #140737488355328 r175 = ~r175;
  always #281474976710656 r176 = ~r176;
  always #562949953421312 r177 = ~r177;
  always #1125899906842624 r178 = ~r178;
  always #2251799813685248 r179 = ~r179;
  always #4503599627370496 r180 = ~r180;
  always #9007199254740992 r181 = ~r181;
  always #18014398509481984 r182 = ~r182;
  always #36028797018963968 r183 = ~r183;
  always #72057594037927936 r184 = ~r184;
  always #144115188075855872 r185 = ~r185;
  always #288230376151711744 r186 = ~r186;
  always #576460752303423488 r187 = ~r187;
  always #1152921504606846976 r188 = ~r188;
  always #2305843009213693952 r189 = ~r189;
  always #4611686018427387904 r190 = ~r190;
  always #9223372036854775808 r191 = ~r191;
  always #1 r192 = ~r192;
  always #2 r193 = ~r193;
  always #4 r194 = ~r194;
  always #8 r195 = ~r195;
  always #16 r196 = ~r196;
  always #32 r197 = ~r197;
  always #64 r198 = ~r198;
  always #128 r199 = ~r199;
  always #256 r200 = ~r200;
  always #512 r201 = ~r201;
  always #1024 r202 = ~r202;
  always #2048 r203 = ~r203;
  always #4096 r204 = ~r204;
  always #8192 r205 = ~r205;
  always #16384 r206 = ~r206;
  always #32768 r207 = ~r207;
  always #65536 r208 = ~r208;
  always #131072 r209 = ~r209;
  always #262144 r210 = ~r210;
  always #524288 r211 = ~r211;
  always #1048576 r212 = ~r212;
  always #2097152 r213 = ~r213;
  always #4194304 r214 = ~r214;
  always #8388608 r215 = ~r215;
  always #16777216 r216 = ~r216;
  always #33554432 r217 = ~r217;
  always #67108864 r218 = ~r218;
  always #134217728 r219 = ~r219;
  always #268435456 r220 = ~r220;
  always #536870912 r221 = ~r221;
  always #1073741824 r222 = ~r222;
  always #2147483648 r223 = ~r223;
  always #4294967296 r224 = ~r224;
  always #8589934592 r225 = ~r225;
  always #17179869184 r226 = ~r226;
  always #34359738368 r227 = ~r227;
  always #68719476736 r228 = ~r228;
  always #137438953472 r229 = ~r229;
  always #274877906944 r230 = ~r230;
  always #549755813888 r231 = ~r231;
  always #1099511627776 r232 = ~r232;
  always #2199023255552 r233 = ~r233;
  always #4398046511104 r234 = ~r234;
  always #8796093022208 r235 = ~r235;
  always #17592186044416 r236 = ~r236;
  always #35184372088832 r237 = ~r237;
  always #70368744177664 r238 = ~r238;
  always #140737488355328 r239 = ~r239;
  always #281474976710656 r240 = ~r240;
  always #562949953421312 r241 = ~r241;
  always #1125899906842624 r242 = ~r242;
  always #2251799813685248 r243 = ~r243;
  always #4503599627370496 r244 = ~r244;
  always #9007199254740992 r245 = ~r245;
  always #18014398509481984 r246 = ~r246;
  always #36028797018963968 r247 = ~r247;
  always #72057594037927936 r248 = ~r248;
  always #144115188075855872 r249 = ~r249;
  always #288230376151711744 r250 = ~r250;
  always #576460752303423488 r251 = ~r251;
  always #1152921504606846976 r252 = ~r252;
  always #2305843009213693952 r253 = ~r253;
  always #4611686018427387904 r254 = ~r254;
  always #9223372036854775808 r255 = ~r255;
  always #1 r256 = ~r256;
  always #2 r257 = ~r257;
  always #4 r258 = ~r258;
  always #8 r259 = ~r259;
  always #16 r260 = ~r260;
  always #32 r261 = ~r261;
  always #64 r262 = ~r262;
  always #128 r263 = ~r263;
  always #256 r264 = ~r264;
  always #512 r265 = ~r265;
  always #1024 r266 = ~r266;
  always #2048 r267 = ~r267;
  always #4096 r268 = ~r268;
  always #8192 r269 = ~r269;
  always #16384 r270 = ~r270;
  always #32768 r271 = ~r271;
  always #65536 r272 = ~r272;
  always #131072 r273 = ~r273;
  always #262144 r274 = ~r274;
  always #524288 r275 = ~r275;
  always #1048576 r276 = ~r276;
  always #2097152 r277 = ~r277;
  always #4194304 r278 = ~r278;
  always #8388608 r279 = ~r279;
  always #16777216 r280 = ~r280;
  always #33554432 r281 = ~r281;
  always #67108864 r282 = ~r282;
  always #134217728 r283 = ~r283;
  always #268435456 r284 = ~r284;
  always #536870912 r285 = ~r285;
  always #1073741824 r286 = ~r286;
  always #2147483648 r287 = ~r287;
  always #4294967296 r288 = ~r288;
  always #8589934592 r289 = ~r289;
  always #17179869184 r290 = ~r290;
  always #34359738368 r291 = ~r291;
  always #68719476736 r292 = ~r292;
  always #137438953472 r293 = ~r293;
  always #274877906944 r294 = ~r294;
  always #549755813888 r295 = ~r295;
  always #1099511627776 r296 = ~r296;
  always #2199023255552 r297 = ~r297;
  always #4398046511104 r298 = ~r298;
  always #8796093022208 r299 = ~r299;
  always #17592186044416 r300 = ~r300;
  always #35184372088832 r301 = ~r301;
  always #70368744177664 r302 = ~r302;
  always #140737488355328 r303 = ~r303;
  always #281474976710656 r304 = ~r304;
  always #562949953421312 r305 = ~r305;
  always #1125899906842624 r306 = ~r306;
  always #2251799813685248 r307 = ~r307;
  always #4503599627370496 r308 = ~r308;
  always #9007199254740992 r309 = ~r309;
  always #18014398509481984 r310 = ~r310;
  always #36028797018963968 r311 = ~r311;
  always #72057594037927936 r312 = ~r312;
  always #144115188075855872 r313 = ~r313;
  always #288230376151711744 r314 = ~r314;
  always #576460752303423488 r315 = ~r315;
  always #1152921504606846976 r316 = ~r316;
  always #2305843009213693952 r317 = ~r317;
  always #4611686018427387904 r318 = ~r318;
  always #9223372036854775808 r319 = ~r319;
  always #1 r320 = ~r320;
  always #2 r321 = ~r321;
  always #4 r322 = ~r322;
  always #8 r323 = ~r323;
  always #16 r324 = ~r324;
  always #32 r325 = ~r325;
  always #64 r326 = ~r326;
  always #128 r327 = ~r327;
  always #256 r328 = ~r328;
  always #512 r329 = ~r329;
  always #1024 r330 = ~r330;
  always #2048 r331 = ~r331;
  always #4096 r332 = ~r332;
  always #8192 r333 = ~r333;
  always #16384 r334 = ~r334;
  always #32768 r335 = ~r335;
  always #65536 r336 = ~r336;
  always #131072 r337 = ~r337;
  always #262144 r338 = ~r338;
  always #524288 r339 = ~r339;
  always #1048576 r340 = ~r340;
  always #2097152 r341 = ~r341;
  always #4194304 r342 = ~r342;
  always #8388608 r343 = ~r343;
  always #16777216 r344 = ~r344;
  always #33554432 r345 = ~r345;
  always #67108864 r346 = ~r346;
  always #134217728 r347 = ~r347;
  always #268435456 r348 = ~r348;
  always #536870912 r349 = ~r349;
  always #1073741824 r350 = ~r350;
  always #2147483648 r351 = ~r351;
  always #4294967296 r352 = ~r352;
  always #8589934592 r353 = ~r353;
  always #17179869184 r354 = ~r354;
  always #34359738368 r355 = ~r355;
  always #68719476736 r356 = ~r356;
  always #137438953472 r357 = ~r357;
  always #274877906944 r358 = ~r358;
  always #549755813888 r359 = ~r359;
  always #1099511627776 r360 = ~r360;
  always #2199023255552 r361 = ~r361;
  always #4398046511104 r362 = ~r362;
  always #8796093022208 r363 = ~r363;
  always #17592186044416 r364 = ~r364;
  always #35184372088832 r365 = ~r365;
  always #70368744177664 r366 = ~r366;
  always #140737488355328 r367 = ~r367;
  always #281474976710656 r368 = ~r368;
  always #562949953421312 r369 = ~r369;
  always #1125899906842624 r370 = ~r370;
  always #2251799813685248 r371 = ~r371;
  always #4503599627370496 r372 = ~r372;
  always #9007199254740992 r373 = ~r373;
  always #18014398509481984 r374 = ~r374;
  always #36028797018963968 r375 = ~r375;
  always #72057594037927936 r376 = ~r376;
  always #144115188075855872 r377 = ~r377;
  always #288230376151711744 r378 = ~r378;
  always #576460752303423488 r379 = ~r379;
  always #1152921504606846976 r380 = ~r380;
  always #2305843009213693952 r381 = ~r381;
  always #4611686018427387904 r382 = ~r382;
  always #9223372036854775808 r383 = ~r383;
  always #1 r384 = ~r384;
  always #2 r385 = ~r385;
  always #4 r386 = ~r386;
  always #8 r387 = ~r387;
  always #16 r388 = ~r388;
  always #32 r389 = ~r389;
  always #64 r390 = ~r390;
  always #128 r391 = ~r391;
  always #256 r392 = ~r392;
  always #512 r393 = ~r393;
  always #1024 r394 = ~r394;
  always #2048 r395 = ~r395;
  always #4096 r396 = ~r396;
  always #8192 r397 = ~r397;
  always #16384 r398 = ~r398;
  always #32768 r399 = ~r399;
  always #65536 r400 = ~r400;
  always #131072 r401 = ~r401;
  always #262144 r402 = ~r402;
  always #524288 r403 = ~r403;
  always #1048576 r404 = ~r404;
  always #2097152 r405 = ~r405;
  always #4194304 r406 = ~r406;
  always #8388608 r407 = ~r407;
  always #16777216 r408 = ~r408;
  always #33554432 r409 = ~r409;
  always #67108864 r410 = ~r410;
  always #134217728 r411 = ~r411;
  always #268435456 r412 = ~r412;
  always #536870912 r413 = ~r413;
  always #1073741824 r414 = ~r414;
  always #2147483648 r415 = ~r415;
  always #4294967296 r416 = ~r416;
  always #8589934592 r417 = ~r417;
  always #17179869184 r418 = ~r418;
  always #34359738368 r419 = ~r419;
  always #68719476736 r420 = ~r420;
  always #137438953472 r421 = ~r421;
  always #274877906944 r422 = ~r422;
  always #549755813888 r423 = ~r423;
  always #1099511627776 r424 = ~r424;
  always #2199023255552 r425 = ~r425;
  always #4398046511104 r426 = ~r426;
  always #8796093022208 r427 = ~r427;
  always #17592186044416 r428 = ~r428;
  always #35184372088832 r429 = ~r429;
  always #70368744177664 r430 = ~r430;
  always #140737488355328 r431 = ~r431;
  always #281474976710656 r432 = ~r432;
  always #562949953421312 r433 = ~r433;
  always #1125899906842624 r434 = ~r434;
  always #2251799813685248 r435 = ~r435;
  always #4503599627370496 r436 = ~r436;
  always #9007199254740992 r437 = ~r437;
  always #18014398509481984 r438 = ~r438;
  always #36028797018963968 r439 = ~r439;
  always #72057594037927936 r440 = ~r440;
  always #144115188075855872 r441 = ~r441;
  always #288230376151711744 r442 = ~r442;
  always #576460752303423488 r443 = ~r443;
  always #1152921504606846976 r444 = ~r444;
  always #2305843009213693952 r445 = ~r445;
  always #4611686018427387904 r446 = ~r446;
  always #9223372036854775808 r447 = ~r447;
  always #1 r448 = ~r448;
  always #2 r449 = ~r449;
  always #4 r450 = ~r450;
  always #8 r451 = ~r451;
  always #16 r452 = ~r452;
  always #32 r453 = ~r453;
  always #64 r454 = ~r454;
  always #128 r455 = ~r455;
  always #256 r456 = ~r456;
  always #512 r457 = ~r457;
  always #1024 r458 = ~r458;
  always #2048 r459 = ~r459;
  always #4096 r460 = ~r460;
  always #8192 r461 = ~r461;
  always #16384 r462 = ~r462;
  always #32768 r463 = ~r463;
  always #65536 r464 = ~r464;
  always #131072 r465 = ~r465;
  always #262144 r466 = ~r466;
  always #524288 r467 = ~r467;
  always #1048576 r468 = ~r468;
  always #2097152 r469 = ~r469;
  always #4194304 r470 = ~r470;
  always #8388608 r471 = ~r471;
  always #16777216 r472 = ~r472;
  always #33554432 r473 = ~r473;
  always #67108864 r474 = ~r474;
  always #134217728 r475 = ~r475;
  always #268435456 r476 = ~r476;
  always #536870912 r477 = ~r477;
  always #1073741824 r478 = ~r478;
  always #2147483648 r479 = ~r479;
  always #4294967296 r480 = ~r480;
  always #8589934592 r481 = ~r481;
  always #17179869184 r482 = ~r482;
  always #34359738368 r483 = ~r483;
  always #68719476736 r484 = ~r484;
  always #137438953472 r485 = ~r485;
  always #274877906944 r486 = ~r486;
  always #549755813888 r487 = ~r487;
  always #1099511627776 r488 = ~r488;
  always #2199023255552 r489 = ~r489;
  always #4398046511104 r490 = ~r490;
  always #8796093022208 r491 = ~r491;
  always #17592186044416 r492 = ~r492;
  always #35184372088832 r493 = ~r493;
  always #70368744177664 r494 = ~r494;
  always #140737488355328 r495 = ~r495;
  always #281474976710656 r496 = ~r496;
  always #562949953421312 r497 = ~r497;
  always #1125899906842624 r498 = ~r498;
  always #2251799813685248 r499 = ~r499;
  always #4503599627370496 r500 = ~r500;
  always #9007199254740992 r501 = ~r501;
  always #18014398509481984 r502 = ~r502;
  always #36028797018963968 r503 = ~r503;
  always #72057594037927936 r504 = ~r504;
  always #144115188075855872 r505 = ~r505;
  always #288230376151711744 r506 = ~r506;
  always #576460752303423488 r507 = ~r507;
  always #1152921504606846976 r508 = ~r508;
  always #2305843009213693952 r509 = ~r509;
  always #4611686018427387904 r510 = ~r510;
  always #9223372036854775808 r511 = ~r511;
  always #1 r512 = ~r512;
  always #2 r513 = ~r513;
  always #4 r514 = ~r514;
  always #8 r515 = ~r515;
  always #16 r516 = ~r516;
  always #32 r517 = ~r517;
  always #64 r518 = ~r518;
  always #128 r519 = ~r519;
  always #256 r520 = ~r520;
  always #512 r521 = ~r521;
  always #1024 r522 = ~r522;
  always #2048 r523 = ~r523;
  always #4096 r524 = ~r524;
  always #8192 r525 = ~r525;
  always #16384 r526 = ~r526;
  always #32768 r527 = ~r527;
  always #65536 r528 = ~r528;
  always #131072 r529 = ~r529;
  always #262144 r530 = ~r530;
  always #524288 r531 = ~r531;
  always #1048576 r532 = ~r532;
  always #2097152 r533 = ~r533;
  always #4194304 r534 = ~r534;
  always #8388608 r535 = ~r535;
  always #16777216 r536 = ~r536;
  always #33554432 r537 = ~r537;
  always #67108864 r538 = ~r538;
  always #134217728 r539 = ~r539;
  always #268435456 r540 = ~r540;
  always #536870912 r541 = ~r541;
  always #1073741824 r542 = ~r542;
  always #2147483648 r543 = ~r543;
  always #4294967296 r544 = ~r544;
  always #8589934592 r545 = ~r545;
  always #17179869184 r546 = ~r546;
  always #34359738368 r547 = ~r547;
  always #68719476736 r548 = ~r548;
  always #137438953472 r549 = ~r549;
  always #274877906944 r550 = ~r550;
  always #549755813888 r551 = ~r551;
  always #1099511627776 r552 = ~r552;
  always #2199023255552 r553 = ~r553;
  always #4398046511104 r554 = ~r554;
  always #8796093022208 r555 = ~r555;
  always #17592186044416 r556 = ~r556;
  always #35184372088832 r557 = ~r557;
  always #70368744177664 r558 = ~r558;
  always #140737488355328 r559 = ~r559;
  always #281474976710656 r560 = ~r560;
  always #562949953421312 r561 = ~r561;
  always #1125899906842624 r562 = ~r562;
  always #2251799813685248 r563 = ~r563;
  always #4503599627370496 r564 = ~r564;
  always #9007199254740992 r565 = ~r565;
  always #18014398509481984 r566 = ~r566;
  always #36028797018963968 r567 = ~r567;
  always #72057594037927936 r568 = ~r568;
  always #144115188075855872 r569 = ~r569;
  always #288230376151711744 r570 = ~r570;
  always #576460752303423488 r571 = ~r571;
  always #1152921504606846976 r572 = ~r572;
  always #2305843009213693952 r573 = ~r573;
  always #4611686018427387904 r574 = ~r574;
  always #9223372036854775808 r575 = ~r575;
  always #1 r576 = ~r576;
  always #2 r577 = ~r577;
  always #4 r578 = ~r578;
  always #8 r579 = ~r579;
  always #16 r580 = ~r580;
  always #32 r581 = ~r581;
  always #64 r582 = ~r582;
  always #128 r583 = ~r583;
  always #256 r584 = ~r584;
  always #512 r585 = ~r585;
  always #1024 r586 = ~r586;
  always #2048 r587 = ~r587;
  always #4096 r588 = ~r588;
  always #8192 r589 = ~r589;
  always #16384 r590 = ~r590;
  always #32768 r591 = ~r591;
  always #65536 r592 = ~r592;
  always #131072 r593 = ~r593;
  always #262144 r594 = ~r594;
  always #524288 r595 = ~r595;
  always #1048576 r596 = ~r596;
  always #2097152 r597 = ~r597;
  always #4194304 r598 = ~r598;
  always #8388608 r599 = ~r599;
  always #16777216 r600 = ~r600;
  always #33554432 r601 = ~r601;
  always #67108864 r602 = ~r602;
  always #134217728 r603 = ~r603;
  always #268435456 r604 = ~r604;
  always #536870912 r605 = ~r605;
  always #1073741824 r606 = ~r606;
  always #2147483648 r607 = ~r607;
  always #4294967296 r608 = ~r608;
  always #8589934592 r609 = ~r609;
  always #17179869184 r610 = ~r610;
  always #34359738368 r611 = ~r611;
  always #68719476736 r612 = ~r612;
  always #137438953472 r613 = ~r613;
  always #274877906944 r614 = ~r614;
  always #549755813888 r615 = ~r615;
  always #1099511627776 r616 = ~r616;
  always #2199023255552 r617 = ~r617;
  always #4398046511104 r618 = ~r618;
  always #8796093022208 r619 = ~r619;
  always #17592186044416 r620 = ~r620;
  always #35184372088832 r621 = ~r621;
  always #70368744177664 r622 = ~r622;
  always #140737488355328 r623 = ~r623;
  always #281474976710656 r624 = ~r624;
  always #562949953421312 r625 = ~r625;
  always #1125899906842624 r626 = ~r626;
  always #2251799813685248 r627 = ~r627;
  always #4503599627370496 r628 = ~r628;
  always #9007199254740992 r629 = ~r629;
  always #18014398509481984 r630 = ~r630;
  always #36028797018963968 r631 = ~r631;
  always #72057594037927936 r632 = ~r632;
  always #144115188075855872 r633 = ~r633;
  always #288230376151711744 r634 = ~r634;
  always #576460752303423488 r635 = ~r635;
  always #1152921504606846976 r636 = ~r636;
  always #2305843009213693952 r637 = ~r637;
  always #4611686018427387904 r638 = ~r638;
  always #9223372036854775808 r639 = ~r639;
  always #1 r640 = ~r640;
  always #2 r641 = ~r641;
  always #4 r642 = ~r642;
  always #8 r643 = ~r643;
  always #16 r644 = ~r644;
  always #32 r645 = ~r645;
  always #64 r646 = ~r646;
  always #128 r647 = ~r647;
  always #256 r648 = ~r648;
  always #512 r649 = ~r649;
  always #1024 r650 = ~r650;
  always #2048 r651 = ~r651;
  always #4096 r652 = ~r652;
  always #8192 r653 = ~r653;
  always #16384 r654 = ~r654;
  always #32768 r655 = ~r655;
  always #65536 r656 = ~r656;
  always #131072 r657 = ~r657;
  always #262144 r658 = ~r658;
  always #524288 r659 = ~r659;
  always #1048576 r660 = ~r660;
  always #2097152 r661 = ~r661;
  always #4194304 r662 = ~r662;
  always #8388608 r663 = ~r663;
  always #16777216 r664 = ~r664;
  always #33554432 r665 = ~r665;
  always #67108864 r666 = ~r666;
  always #134217728 r667 = ~r667;
  always #268435456 r668 = ~r668;
  always #536870912 r669 = ~r669;
  always #1073741824 r670 = ~r670;
  always #2147483648 r671 = ~r671;
  always #4294967296 r672 = ~r672;
  always #8589934592 r673 = ~r673;
  always #17179869184 r674 = ~r674;
  always #34359738368 r675 = ~r675;
  always #68719476736 r676 = ~r676;
  always #137438953472 r677 = ~r677;
  always #274877906944 r678 = ~r678;
  always #549755813888 r679 = ~r679;
  always #1099511627776 r680 = ~r680;
  always #2199023255552 r681 = ~r681;
  always #4398046511104 r682 = ~r682;
  always #8796093022208 r683 = ~r683;
  always #17592186044416 r684 = ~r684;
  always #35184372088832 r685 = ~r685;
  always #70368744177664 r686 = ~r686;
  always #140737488355328 r687 = ~r687;
  always #281474976710656 r688 = ~r688;
  always #562949953421312 r689 = ~r689;
  always #1125899906842624 r690 = ~r690;
  always #2251799813685248 r691 = ~r691;
  always #4503599627370496 r692 = ~r692;
  always #9007199254740992 r693 = ~r693;
  always #18014398509481984 r694 = ~r694;
  always #36028797018963968 r695 = ~r695;
  always #72057594037927936 r696 = ~r696;
  always #144115188075855872 r697 = ~r697;
  always #288230376151711744 r698 = ~r698;
  always #576460752303423488 r699 = ~r699;
  always #1152921504606846976 r700 = ~r700;
  always #2305843009213693952 r701 = ~r701;
  always #4611686018427387904 r702 = ~r702;
  always #9223372036854775808 r703 = ~r703;
  always #1 r704 = ~r704;
  always #2 r705 = ~r705;
  always #4 r706 = ~r706;
  always #8 r707 = ~r707;
  always #16 r708 = ~r708;
  always #32 r709 = ~r709;
  always #64 r710 = ~r710;
  always #128 r711 = ~r711;
  always #256 r712 = ~r712;
  always #512 r713 = ~r713;
  always #1024 r714 = ~r714;
  always #2048 r715 = ~r715;
  always #4096 r716 = ~r716;
  always #8192 r717 = ~r717;
  always #16384 r718 = ~r718;
  always #32768 r719 = ~r719;
  always #65536 r720 = ~r720;
  always #131072 r721 = ~r721;
  always #262144 r722 = ~r722;
  always #524288 r723 = ~r723;
  always #1048576 r724 = ~r724;
  always #2097152 r725 = ~r725;
  always #4194304 r726 = ~r726;
  always #8388608 r727 = ~r727;
  always #16777216 r728 = ~r728;
  always #33554432 r729 = ~r729;
  always #67108864 r730 = ~r730;
  always #134217728 r731 = ~r731;
  always #268435456 r732 = ~r732;
  always #536870912 r733 = ~r733;
  always #1073741824 r734 = ~r734;
  always #2147483648 r735 = ~r735;
  always #4294967296 r736 = ~r736;
  always #8589934592 r737 = ~r737;
  always #17179869184 r738 = ~r738;
  always #34359738368 r739 = ~r739;
  always #68719476736 r740 = ~r740;
  always #137438953472 r741 = ~r741;
  always #274877906944 r742 = ~r742;
  always #549755813888 r743 = ~r743;
  always #1099511627776 r744 = ~r744;
  always #2199023255552 r745 = ~r745;
  always #4398046511104 r746 = ~r746;
  always #8796093022208 r747 = ~r747;
  always #17592186044416 r748 = ~r748;
  always #35184372088832 r749 = ~r749;
  always #70368744177664 r750 = ~r750;
  always #140737488355328 r751 = ~r751;
  always #281474976710656 r752 = ~r752;
  always #562949953421312 r753 = ~r753;
  always #1125899906842624 r754 = ~r754;
  always #2251799813685248 r755 = ~r755;
  always #4503599627370496 r756 = ~r756;
  always #9007199254740992 r757 = ~r757;
  always #18014398509481984 r758 = ~r758;
  always #36028797018963968 r759 = ~r759;
  always #72057594037927936 r760 = ~r760;
  always #144115188075855872 r761 = ~r761;
  always #288230376151711744 r762 = ~r762;
  always #576460752303423488 r763 = ~r763;
  always #1152921504606846976 r764 = ~r764;
  always #2305843009213693952 r765 = ~r765;
  always #4611686018427387904 r766 = ~r766;
  always #9223372036854775808 r767 = ~r767;
  always #1 r768 = ~r768;
  always #2 r769 = ~r769;
  always #4 r770 = ~r770;
  always #8 r771 = ~r771;
  always #16 r772 = ~r772;
  always #32 r773 = ~r773;
  always #64 r774 = ~r774;
  always #128 r775 = ~r775;
  always #256 r776 = ~r776;
  always #512 r777 = ~r777;
  always #1024 r778 = ~r778;
  always #2048 r779 = ~r779;
  always #4096 r780 = ~r780;
  always #8192 r781 = ~r781;
  always #16384 r782 = ~r782;
  always #32768 r783 = ~r783;
  always #65536 r784 = ~r784;
  always #131072 r785 = ~r785;
  always #262144 r786 = ~r786;
  always #524288 r787 = ~r787;
  always #1048576 r788 = ~r788;
  always #2097152 r789 = ~r789;
  always #4194304 r790 = ~r790;
  always #8388608 r791 = ~r791;
  always #16777216 r792 = ~r792;
  always #33554432 r793 = ~r793;
  always #67108864 r794 = ~r794;
  always #134217728 r795 = ~r795;
  always #268435456 r796 = ~r796;
  always #536870912 r797 = ~r797;
  always #1073741824 r798 = ~r798;
  always #2147483648 r799 = ~r799;
  always #4294967296 r800 = ~r800;
  always #8589934592 r801 = ~r801;
  always #17179869184 r802 = ~r802;
  always #34359738368 r803 = ~r803;
  always #68719476736 r804 = ~r804;
  always #137438953472 r805 = ~r805;
  always #274877906944 r806 = ~r806;
  always #549755813888 r807 = ~r807;
  always #1099511627776 r808 = ~r808;
  always #2199023255552 r809 = ~r809;
  always #4398046511104 r810 = ~r810;
  always #8796093022208 r811 = ~r811;
  always #17592186044416 r812 = ~r812;
  always #35184372088832 r813 = ~r813;
  always #70368744177664 r814 = ~r814;
  always #140737488355328 r815 = ~r815;
  always #281474976710656 r816 = ~r816;
  always #562949953421312 r817 = ~r817;
  always #1125899906842624 r818 = ~r818;
  always #2251799813685248 r819 = ~r819;
  always #4503599627370496 r820 = ~r820;
  always #9007199254740992 r821 = ~r821;
  always #18014398509481984 r822 = ~r822;
  always #36028797018963968 r823 = ~r823;
  always #72057594037927936 r824 = ~r824;
  always #144115188075855872 r825 = ~r825;
  always #288230376151711744 r826 = ~r826;
  always #576460752303423488 r827 = ~r827;
  always #1152921504606846976 r828 = ~r828;
  always #2305843009213693952 r829 = ~r829;
  always #4611686018427387904 r830 = ~r830;
  always #9223372036854775808 r831 = ~r831;
  always #1 r832 = ~r832;
  always #2 r833 = ~r833;
  always #4 r834 = ~r834;
  always #8 r835 = ~r835;
  always #16 r836 = ~r836;
  always #32 r837 = ~r837;
  always #64 r838 = ~r838;
  always #128 r839 = ~r839;
  always #256 r840 = ~r840;
  always #512 r841 = ~r841;
  always #1024 r842 = ~r842;
  always #2048 r843 = ~r843;
  always #4096 r844 = ~r844;
  always #8192 r845 = ~r845;
  always #16384 r846 = ~r846;
  always #32768 r847 = ~r847;
  always #65536 r848 = ~r848;
  always #131072 r849 = ~r849;
  always #262144 r850 = ~r850;
  always #524288 r851 = ~r851;
  always #1048576 r852 = ~r852;
  always #2097152 r853 = ~r853;
  always #4194304 r854 = ~r854;
  always #8388608 r855 = ~r855;
  always #16777216 r856 = ~r856;
  always #33554432 r857 = ~r857;
  always #67108864 r858 = ~r858;
  always #134217728 r859 = ~r859;
  always #268435456 r860 = ~r860;
  always #536870912 r861 = ~r861;
  always #1073741824 r862 = ~r862;
  always #2147483648 r863 = ~r863;
  always #4294967296 r864 = ~r864;
  always #8589934592 r865 = ~r865;
  always #17179869184 r866 = ~r866;
  always #34359738368 r867 = ~r867;
  always #68719476736 r868 = ~r868;
  always #137438953472 r869 = ~r869;
  always #274877906944 r870 = ~r870;
  always #549755813888 r871 = ~r871;
  always #1099511627776 r872 = ~r872;
  always #2199023255552 r873 = ~r873;
  always #4398046511104 r874 = ~r874;
  always #8796093022208 r875 = ~r875;
  always #17592186044416 r876 = ~r876;
  always #35184372088832 r877 = ~r877;
  always #70368744177664 r878 = ~r878;
  always #140737488355328 r879 = ~r879;
  always #281474976710656 r880 = ~r880;
  always #562949953421312 r881 = ~r881;
  always #1125899906842624 r882 = ~r882;
  always #2251799813685248 r883 = ~r883;
  always #4503599627370496 r884 = ~r884;
  always #9007199254740992 r885 = ~r885;
  always #18014398509481984 r886 = ~r886;
  always #36028797018963968 r887 = ~r887;
  always #72057594037927936 r888 = ~r888;
  always #144115188075855872 r889 = ~r889;
  always #288230376151711744 r890 = ~r890;
  always #576460752303423488 r891 = ~r891;
  always #1152921504606846976 r892 = ~r892;
  always #2305843009213693952 r893 = ~r893;
  always #4611686018427387904 r894 = ~r894;
  always #9223372036854775808 r895 = ~r895;
  always #1 r896 = ~r896;
  always #2 r897 = ~r897;
  always #4 r898 = ~r898;
  always #8 r899 = ~r899;
  always #16 r900 = ~r900;
  always #32 r901 = ~r901;
  always #64 r902 = ~r902;
  always #128 r903 = ~r903;
  always #256 r904 = ~r904;
  always #512 r905 = ~r905;
  always #1024 r906 = ~r906;
  always #2048 r907 = ~r907;
  always #4096 r908 = ~r908;
  always #8192 r909 = ~r909;
  always #16384 r910 = ~r910;
  always #32768 r911 = ~r911;
  always #65536 r912 = ~r912;
  always #131072 r913 = ~r913;
  always #262144 r914 = ~r914;
  always #524288 r915 = ~r915;
  always #1048576 r916 = ~r916;
  always #2097152 r917 = ~r917;
  always #4194304 r918 = ~r918;
  always #8388608 r919 = ~r919;
  always #16777216 r920 = ~r920;
  always #33554432 r921 = ~r921;
  always #67108864 r922 = ~r922;
  always #134217728 r923 = ~r923;
  always #268435456 r924 = ~r924;
  always #536870912 r925 = ~r925;
  always #1073741824 r926 = ~r926;
  always #2147483648 r927 = ~r927;
  always #4294967296 r928 = ~r928;
  always #8589934592 r929 = ~r929;
  always #17179869184 r930 = ~r930;
  always #34359738368 r931 = ~r931;
  always #68719476736 r932 = ~r932;
  always #137438953472 r933 = ~r933;
  always #274877906944 r934 = ~r934;
  always #549755813888 r935 = ~r935;
  always #1099511627776 r936 = ~r936;
  always #2199023255552 r937 = ~r937;
  always #4398046511104 r938 = ~r938;
  always #8796093022208 r939 = ~r939;
  always #17592186044416 r940 = ~r940;
  always #35184372088832 r941 = ~r941;
  always #70368744177664 r942 = ~r942;
  always #140737488355328 r943 = ~r943;
  always #281474976710656 r944 = ~r944;
  always #562949953421312 r945 = ~r945;
  always #1125899906842624 r946 = ~r946;
  always #2251799813685248 r947 = ~r947;
  always #4503599627370496 r948 = ~r948;
  always #9007199254740992 r949 = ~r949;
  always #18014398509481984 r950 = ~r950;
  always #36028797018963968 r951 = ~r951;
  always #72057594037927936 r952 = ~r952;
  always #144115188075855872 r953 = ~r953;
  always #288230376151711744 r954 = ~r954;
  always #576460752303423488 r955 = ~r955;
  always #1152921504606846976 r956 = ~r956;
  always #2305843009213693952 r957 = ~r957;
  always #4611686018427387904 r958 = ~r958;
  always #9223372036854775808 r959 = ~r959;
  always #1 r960 = ~r960;
  always #2 r961 = ~r961;
  always #4 r962 = ~r962;
  always #8 r963 = ~r963;
  always #16 r964 = ~r964;
  always #32 r965 = ~r965;
  always #64 r966 = ~r966;
  always #128 r967 = ~r967;
  always #256 r968 = ~r968;
  always #512 r969 = ~r969;
  always #1024 r970 = ~r970;
  always #2048 r971 = ~r971;
  always #4096 r972 = ~r972;
  always #8192 r973 = ~r973;
  always #16384 r974 = ~r974;
  always #32768 r975 = ~r975;
  always #65536 r976 = ~r976;
  always #131072 r977 = ~r977;
  always #262144 r978 = ~r978;
  always #524288 r979 = ~r979;
  always #1048576 r980 = ~r980;
  always #2097152 r981 = ~r981;
  always #4194304 r982 = ~r982;
  always #8388608 r983 = ~r983;
  always #16777216 r984 = ~r984;
  always #33554432 r985 = ~r985;
  always #67108864 r986 = ~r986;
  always #134217728 r987 = ~r987;
  always #268435456 r988 = ~r988;
  always #536870912 r989 = ~r989;
  always #1073741824 r990 = ~r990;
  always #2147483648 r991 = ~r991;
  always #4294967296 r992 = ~r992;
  always #8589934592 r993 = ~r993;
  always #17179869184 r994 = ~r994;
  always #34359738368 r995 = ~r995;
  always #68719476736 r996 = ~r996;
  always #137438953472 r997 = ~r997;
  always #274877906944 r998 = ~r998;
  always #549755813888 r999 = ~r999;
  always #1099511627776 r1000 = ~r1000;
  always #2199023255552 r1001 = ~r1001;
  always #4398046511104 r1002 = ~r1002;
  always #8796093022208 r1003 = ~r1003;
  always #17592186044416 r1004 = ~r1004;
  always #35184372088832 r1005 = ~r1005;
  always #70368744177664 r1006 = ~r1006;
  always #140737488355328 r1007 = ~r1007;
  always #281474976710656 r1008 = ~r1008;
  always #562949953421312 r1009 = ~r1009;
  always #1125899906842624 r1010 = ~r1010;
  always #2251799813685248 r1011 = ~r1011;
  always #4503599627370496 r1012 = ~r1012;
  always #9007199254740992 r1013 = ~r1013;
  always #18014398509481984 r1014 = ~r1014;
  always #36028797018963968 r1015 = ~r1015;
  always #72057594037927936 r1016 = ~r1016;
  always #144115188075855872 r1017 = ~r1017;
  always #288230376151711744 r1018 = ~r1018;
  always #576460752303423488 r1019 = ~r1019;
  always #1152921504606846976 r1020 = ~r1020;
  always #2305843009213693952 r1021 = ~r1021;
  always #4611686018427387904 r1022 = ~r1022;
  always #9223372036854775808 r1023 = ~r1023;
  always #1 r1024 = ~r1024;
  always #2 r1025 = ~r1025;
  always #4 r1026 = ~r1026;
  always #8 r1027 = ~r1027;
  always #16 r1028 = ~r1028;
  always #32 r1029 = ~r1029;
  always #64 r1030 = ~r1030;
  always #128 r1031 = ~r1031;
  always #256 r1032 = ~r1032;
  always #512 r1033 = ~r1033;
  always #1024 r1034 = ~r1034;
  always #2048 r1035 = ~r1035;
  always #4096 r1036 = ~r1036;
  always #8192 r1037 = ~r1037;
  always #16384 r1038 = ~r1038;
  always #32768 r1039 = ~r1039;
  always #65536 r1040 = ~r1040;
  always #131072 r1041 = ~r1041;
  always #262144 r1042 = ~r1042;
  always #524288 r1043 = ~r1043;
  always #1048576 r1044 = ~r1044;
  always #2097152 r1045 = ~r1045;
  always #4194304 r1046 = ~r1046;
  always #8388608 r1047 = ~r1047;
  always #16777216 r1048 = ~r1048;
  always #33554432 r1049 = ~r1049;
  always #67108864 r1050 = ~r1050;
  always #134217728 r1051 = ~r1051;
  always #268435456 r1052 = ~r1052;
  always #536870912 r1053 = ~r1053;
  always #1073741824 r1054 = ~r1054;
  always #2147483648 r1055 = ~r1055;
  always #4294967296 r1056 = ~r1056;
  always #8589934592 r1057 = ~r1057;
  always #17179869184 r1058 = ~r1058;
  always #34359738368 r1059 = ~r1059;
  always #68719476736 r1060 = ~r1060;
  always #137438953472 r1061 = ~r1061;
  always #274877906944 r1062 = ~r1062;
  always #549755813888 r1063 = ~r1063;
  always #1099511627776 r1064 = ~r1064;
  always #2199023255552 r1065 = ~r1065;
  always #4398046511104 r1066 = ~r1066;
  always #8796093022208 r1067 = ~r1067;
  always #17592186044416 r1068 = ~r1068;
  always #35184372088832 r1069 = ~r1069;
  always #70368744177664 r1070 = ~r1070;
  always #140737488355328 r1071 = ~r1071;
  always #281474976710656 r1072 = ~r1072;
  always #562949953421312 r1073 = ~r1073;
  always #1125899906842624 r1074 = ~r1074;
  always #2251799813685248 r1075 = ~r1075;
  always #4503599627370496 r1076 = ~r1076;
  always #9007199254740992 r1077 = ~r1077;
  always #18014398509481984 r1078 = ~r1078;
  always #36028797018963968 r1079 = ~r1079;
  always #72057594037927936 r1080 = ~r1080;
  always #144115188075855872 r1081 = ~r1081;
  always #288230376151711744 r1082 = ~r1082;
  always #576460752303423488 r1083 = ~r1083;
  always #1152921504606846976 r1084 = ~r1084;
  always #2305843009213693952 r1085 = ~r1085;
  always #4611686018427387904 r1086 = ~r1086;
  always #9223372036854775808 r1087 = ~r1087;
  always #1 r1088 = ~r1088;
  always #2 r1089 = ~r1089;
  always #4 r1090 = ~r1090;
  always #8 r1091 = ~r1091;
  always #16 r1092 = ~r1092;
  always #32 r1093 = ~r1093;
  always #64 r1094 = ~r1094;
  always #128 r1095 = ~r1095;
  always #256 r1096 = ~r1096;
  always #512 r1097 = ~r1097;
  always #1024 r1098 = ~r1098;
  always #2048 r1099 = ~r1099;
  always #4096 r1100 = ~r1100;
  always #8192 r1101 = ~r1101;
  always #16384 r1102 = ~r1102;
  always #32768 r1103 = ~r1103;
  always #65536 r1104 = ~r1104;
  always #131072 r1105 = ~r1105;
  always #262144 r1106 = ~r1106;
  always #524288 r1107 = ~r1107;
  always #1048576 r1108 = ~r1108;
  always #2097152 r1109 = ~r1109;
  always #4194304 r1110 = ~r1110;
  always #8388608 r1111 = ~r1111;
  always #16777216 r1112 = ~r1112;
  always #33554432 r1113 = ~r1113;
  always #67108864 r1114 = ~r1114;
  always #134217728 r1115 = ~r1115;
  always #268435456 r1116 = ~r1116;
  always #536870912 r1117 = ~r1117;
  always #1073741824 r1118 = ~r1118;
  always #2147483648 r1119 = ~r1119;
  always #4294967296 r1120 = ~r1120;
  always #8589934592 r1121 = ~r1121;
  always #17179869184 r1122 = ~r1122;
  always #34359738368 r1123 = ~r1123;
  always #68719476736 r1124 = ~r1124;
  always #137438953472 r1125 = ~r1125;
  always #274877906944 r1126 = ~r1126;
  always #549755813888 r1127 = ~r1127;
  always #1099511627776 r1128 = ~r1128;
  always #2199023255552 r1129 = ~r1129;
  always #4398046511104 r1130 = ~r1130;
  always #8796093022208 r1131 = ~r1131;
  always #17592186044416 r1132 = ~r1132;
  always #35184372088832 r1133 = ~r1133;
  always #70368744177664 r1134 = ~r1134;
  always #140737488355328 r1135 = ~r1135;
  always #281474976710656 r1136 = ~r1136;
  always #562949953421312 r1137 = ~r1137;
  always #1125899906842624 r1138 = ~r1138;
  always #2251799813685248 r1139 = ~r1139;
  always #4503599627370496 r1140 = ~r1140;
  always #9007199254740992 r1141 = ~r1141;
  always #18014398509481984 r1142 = ~r1142;
  always #36028797018963968 r1143 = ~r1143;
  always #72057594037927936 r1144 = ~r1144;
  always #144115188075855872 r1145 = ~r1145;
  always #288230376151711744 r1146 = ~r1146;
  always #576460752303423488 r1147 = ~r1147;
  always #1152921504606846976 r1148 = ~r1148;
  always #2305843009213693952 r1149 = ~r1149;
  always #4611686018427387904 r1150 = ~r1150;
  always #9223372036854775808 r1151 = ~r1151;
  always #1 r1152 = ~r1152;
  always #2 r1153 = ~r1153;
  always #4 r1154 = ~r1154;
  always #8 r1155 = ~r1155;
  always #16 r1156 = ~r1156;
  always #32 r1157 = ~r1157;
  always #64 r1158 = ~r1158;
  always #128 r1159 = ~r1159;
  always #256 r1160 = ~r1160;
  always #512 r1161 = ~r1161;
  always #1024 r1162 = ~r1162;
  always #2048 r1163 = ~r1163;
  always #4096 r1164 = ~r1164;
  always #8192 r1165 = ~r1165;
  always #16384 r1166 = ~r1166;
  always #32768 r1167 = ~r1167;
  always #65536 r1168 = ~r1168;
  always #131072 r1169 = ~r1169;
  always #262144 r1170 = ~r1170;
  always #524288 r1171 = ~r1171;
  always #1048576 r1172 = ~r1172;
  always #2097152 r1173 = ~r1173;
  always #4194304 r1174 = ~r1174;
  always #8388608 r1175 = ~r1175;
  always #16777216 r1176 = ~r1176;
  always #33554432 r1177 = ~r1177;
  always #67108864 r1178 = ~r1178;
  always #134217728 r1179 = ~r1179;
  always #268435456 r1180 = ~r1180;
  always #536870912 r1181 = ~r1181;
  always #1073741824 r1182 = ~r1182;
  always #2147483648 r1183 = ~r1183;
  always #4294967296 r1184 = ~r1184;
  always #8589934592 r1185 = ~r1185;
  always #17179869184 r1186 = ~r1186;
  always #34359738368 r1187 = ~r1187;
  always #68719476736 r1188 = ~r1188;
  always #137438953472 r1189 = ~r1189;
  always #274877906944 r1190 = ~r1190;
  always #549755813888 r1191 = ~r1191;
  always #1099511627776 r1192 = ~r1192;
  always #2199023255552 r1193 = ~r1193;
  always #4398046511104 r1194 = ~r1194;
  always #8796093022208 r1195 = ~r1195;
  always #17592186044416 r1196 = ~r1196;
  always #35184372088832 r1197 = ~r1197;
  always #70368744177664 r1198 = ~r1198;
  always #140737488355328 r1199 = ~r1199;
  always #281474976710656 r1200 = ~r1200;
  always #562949953421312 r1201 = ~r1201;
  always #1125899906842624 r1202 = ~r1202;
  always #2251799813685248 r1203 = ~r1203;
  always #4503599627370496 r1204 = ~r1204;
  always #9007199254740992 r1205 = ~r1205;
  always #18014398509481984 r1206 = ~r1206;
  always #36028797018963968 r1207 = ~r1207;
  always #72057594037927936 r1208 = ~r1208;
  always #144115188075855872 r1209 = ~r1209;
  always #288230376151711744 r1210 = ~r1210;
  always #576460752303423488 r1211 = ~r1211;
  always #1152921504606846976 r1212 = ~r1212;
  always #2305843009213693952 r1213 = ~r1213;
  always #4611686018427387904 r1214 = ~r1214;
  always #9223372036854775808 r1215 = ~r1215;
  always #1 r1216 = ~r1216;
  always #2 r1217 = ~r1217;
  always #4 r1218 = ~r1218;
  always #8 r1219 = ~r1219;
  always #16 r1220 = ~r1220;
  always #32 r1221 = ~r1221;
  always #64 r1222 = ~r1222;
  always #128 r1223 = ~r1223;
  always #256 r1224 = ~r1224;
  always #512 r1225 = ~r1225;
  always #1024 r1226 = ~r1226;
  always #2048 r1227 = ~r1227;
  always #4096 r1228 = ~r1228;
  always #8192 r1229 = ~r1229;
  always #16384 r1230 = ~r1230;
  always #32768 r1231 = ~r1231;
  always #65536 r1232 = ~r1232;
  always #131072 r1233 = ~r1233;
  always #262144 r1234 = ~r1234;
  always #524288 r1235 = ~r1235;
  always #1048576 r1236 = ~r1236;
  always #2097152 r1237 = ~r1237;
  always #4194304 r1238 = ~r1238;
  always #8388608 r1239 = ~r1239;
  always #16777216 r1240 = ~r1240;
  always #33554432 r1241 = ~r1241;
  always #67108864 r1242 = ~r1242;
  always #134217728 r1243 = ~r1243;
  always #268435456 r1244 = ~r1244;
  always #536870912 r1245 = ~r1245;
  always #1073741824 r1246 = ~r1246;
  always #2147483648 r1247 = ~r1247;
  always #4294967296 r1248 = ~r1248;
  always #8589934592 r1249 = ~r1249;
  always #17179869184 r1250 = ~r1250;
  always #34359738368 r1251 = ~r1251;
  always #68719476736 r1252 = ~r1252;
  always #137438953472 r1253 = ~r1253;
  always #274877906944 r1254 = ~r1254;
  always #549755813888 r1255 = ~r1255;
  always #1099511627776 r1256 = ~r1256;
  always #2199023255552 r1257 = ~r1257;
  always #4398046511104 r1258 = ~r1258;
  always #8796093022208 r1259 = ~r1259;
  always #17592186044416 r1260 = ~r1260;
  always #35184372088832 r1261 = ~r1261;
  always #70368744177664 r1262 = ~r1262;
  always #140737488355328 r1263 = ~r1263;
  always #281474976710656 r1264 = ~r1264;
  always #562949953421312 r1265 = ~r1265;
  always #1125899906842624 r1266 = ~r1266;
  always #2251799813685248 r1267 = ~r1267;
  always #4503599627370496 r1268 = ~r1268;
  always #9007199254740992 r1269 = ~r1269;
  always #18014398509481984 r1270 = ~r1270;
  always #36028797018963968 r1271 = ~r1271;
  always #72057594037927936 r1272 = ~r1272;
  always #144115188075855872 r1273 = ~r1273;
  always #288230376151711744 r1274 = ~r1274;
  always #576460752303423488 r1275 = ~r1275;
  always #1152921504606846976 r1276 = ~r1276;
  always #2305843009213693952 r1277 = ~r1277;
  always #4611686018427387904 r1278 = ~r1278;
  always #9223372036854775808 r1279 = ~r1279;
  always #1 r1280 = ~r1280;
  always #2 r1281 = ~r1281;
  always #4 r1282 = ~r1282;
  always #8 r1283 = ~r1283;
  always #16 r1284 = ~r1284;
  always #32 r1285 = ~r1285;
  always #64 r1286 = ~r1286;
  always #128 r1287 = ~r1287;
  always #256 r1288 = ~r1288;
  always #512 r1289 = ~r1289;
  always #1024 r1290 = ~r1290;
  always #2048 r1291 = ~r1291;
  always #4096 r1292 = ~r1292;
  always #8192 r1293 = ~r1293;
  always #16384 r1294 = ~r1294;
  always #32768 r1295 = ~r1295;
  always #65536 r1296 = ~r1296;
  always #131072 r1297 = ~r1297;
  always #262144 r1298 = ~r1298;
  always #524288 r1299 = ~r1299;
  always #1048576 r1300 = ~r1300;
  always #2097152 r1301 = ~r1301;
  always #4194304 r1302 = ~r1302;
  always #8388608 r1303 = ~r1303;
  always #16777216 r1304 = ~r1304;
  always #33554432 r1305 = ~r1305;
  always #67108864 r1306 = ~r1306;
  always #134217728 r1307 = ~r1307;
  always #268435456 r1308 = ~r1308;
  always #536870912 r1309 = ~r1309;
  always #1073741824 r1310 = ~r1310;
  always #2147483648 r1311 = ~r1311;
  always #4294967296 r1312 = ~r1312;
  always #8589934592 r1313 = ~r1313;
  always #17179869184 r1314 = ~r1314;
  always #34359738368 r1315 = ~r1315;
  always #68719476736 r1316 = ~r1316;
  always #137438953472 r1317 = ~r1317;
  always #274877906944 r1318 = ~r1318;
  always #549755813888 r1319 = ~r1319;
  always #1099511627776 r1320 = ~r1320;
  always #2199023255552 r1321 = ~r1321;
  always #4398046511104 r1322 = ~r1322;
  always #8796093022208 r1323 = ~r1323;
  always #17592186044416 r1324 = ~r1324;
  always #35184372088832 r1325 = ~r1325;
  always #70368744177664 r1326 = ~r1326;
  always #140737488355328 r1327 = ~r1327;
  always #281474976710656 r1328 = ~r1328;
  always #562949953421312 r1329 = ~r1329;
  always #1125899906842624 r1330 = ~r1330;
  always #2251799813685248 r1331 = ~r1331;
  always #4503599627370496 r1332 = ~r1332;
  always #9007199254740992 r1333 = ~r1333;
  always #18014398509481984 r1334 = ~r1334;
  always #36028797018963968 r1335 = ~r1335;
  always #72057594037927936 r1336 = ~r1336;
  always #144115188075855872 r1337 = ~r1337;
  always #288230376151711744 r1338 = ~r1338;
  always #576460752303423488 r1339 = ~r1339;
  always #1152921504606846976 r1340 = ~r1340;
  always #2305843009213693952 r1341 = ~r1341;
  always #4611686018427387904 r1342 = ~r1342;
  always #9223372036854775808 r1343 = ~r1343;
  always #1 r1344 = ~r1344;
  always #2 r1345 = ~r1345;
  always #4 r1346 = ~r1346;
  always #8 r1347 = ~r1347;
  always #16 r1348 = ~r1348;
  always #32 r1349 = ~r1349;
  always #64 r1350 = ~r1350;
  always #128 r1351 = ~r1351;
  always #256 r1352 = ~r1352;
  always #512 r1353 = ~r1353;
  always #1024 r1354 = ~r1354;
  always #2048 r1355 = ~r1355;
  always #4096 r1356 = ~r1356;
  always #8192 r1357 = ~r1357;
  always #16384 r1358 = ~r1358;
  always #32768 r1359 = ~r1359;
  always #65536 r1360 = ~r1360;
  always #131072 r1361 = ~r1361;
  always #262144 r1362 = ~r1362;
  always #524288 r1363 = ~r1363;
  always #1048576 r1364 = ~r1364;
  always #2097152 r1365 = ~r1365;
  always #4194304 r1366 = ~r1366;
  always #8388608 r1367 = ~r1367;
  always #16777216 r1368 = ~r1368;
  always #33554432 r1369 = ~r1369;
  always #67108864 r1370 = ~r1370;
  always #134217728 r1371 = ~r1371;
  always #268435456 r1372 = ~r1372;
  always #536870912 r1373 = ~r1373;
  always #1073741824 r1374 = ~r1374;
  always #2147483648 r1375 = ~r1375;
  always #4294967296 r1376 = ~r1376;
  always #8589934592 r1377 = ~r1377;
  always #17179869184 r1378 = ~r1378;
  always #34359738368 r1379 = ~r1379;
  always #68719476736 r1380 = ~r1380;
  always #137438953472 r1381 = ~r1381;
  always #274877906944 r1382 = ~r1382;
  always #549755813888 r1383 = ~r1383;
  always #1099511627776 r1384 = ~r1384;
  always #2199023255552 r1385 = ~r1385;
  always #4398046511104 r1386 = ~r1386;
  always #8796093022208 r1387 = ~r1387;
  always #17592186044416 r1388 = ~r1388;
  always #35184372088832 r1389 = ~r1389;
  always #70368744177664 r1390 = ~r1390;
  always #140737488355328 r1391 = ~r1391;
  always #281474976710656 r1392 = ~r1392;
  always #562949953421312 r1393 = ~r1393;
  always #1125899906842624 r1394 = ~r1394;
  always #2251799813685248 r1395 = ~r1395;
  always #4503599627370496 r1396 = ~r1396;
  always #9007199254740992 r1397 = ~r1397;
  always #18014398509481984 r1398 = ~r1398;
  always #36028797018963968 r1399 = ~r1399;
  always #72057594037927936 r1400 = ~r1400;
  always #144115188075855872 r1401 = ~r1401;
  always #288230376151711744 r1402 = ~r1402;
  always #576460752303423488 r1403 = ~r1403;
  always #1152921504606846976 r1404 = ~r1404;
  always #2305843009213693952 r1405 = ~r1405;
  always #4611686018427387904 r1406 = ~r1406;
  always #9223372036854775808 r1407 = ~r1407;
  always #1 r1408 = ~r1408;
  always #2 r1409 = ~r1409;
  always #4 r1410 = ~r1410;
  always #8 r1411 = ~r1411;
  always #16 r1412 = ~r1412;
  always #32 r1413 = ~r1413;
  always #64 r1414 = ~r1414;
  always #128 r1415 = ~r1415;
  always #256 r1416 = ~r1416;
  always #512 r1417 = ~r1417;
  always #1024 r1418 = ~r1418;
  always #2048 r1419 = ~r1419;
  always #4096 r1420 = ~r1420;
  always #8192 r1421 = ~r1421;
  always #16384 r1422 = ~r1422;
  always #32768 r1423 = ~r1423;
  always #65536 r1424 = ~r1424;
  always #131072 r1425 = ~r1425;
  always #262144 r1426 = ~r1426;
  always #524288 r1427 = ~r1427;
  always #1048576 r1428 = ~r1428;
  always #2097152 r1429 = ~r1429;
  always #4194304 r1430 = ~r1430;
  always #8388608 r1431 = ~r1431;
  always #16777216 r1432 = ~r1432;
  always #33554432 r1433 = ~r1433;
  always #67108864 r1434 = ~r1434;
  always #134217728 r1435 = ~r1435;
  always #268435456 r1436 = ~r1436;
  always #536870912 r1437 = ~r1437;
  always #1073741824 r1438 = ~r1438;
  always #2147483648 r1439 = ~r1439;
  always #4294967296 r1440 = ~r1440;
  always #8589934592 r1441 = ~r1441;
  always #17179869184 r1442 = ~r1442;
  always #34359738368 r1443 = ~r1443;
  always #68719476736 r1444 = ~r1444;
  always #137438953472 r1445 = ~r1445;
  always #274877906944 r1446 = ~r1446;
  always #549755813888 r1447 = ~r1447;
  always #1099511627776 r1448 = ~r1448;
  always #2199023255552 r1449 = ~r1449;
  always #4398046511104 r1450 = ~r1450;
  always #8796093022208 r1451 = ~r1451;
  always #17592186044416 r1452 = ~r1452;
  always #35184372088832 r1453 = ~r1453;
  always #70368744177664 r1454 = ~r1454;
  always #140737488355328 r1455 = ~r1455;
  always #281474976710656 r1456 = ~r1456;
  always #562949953421312 r1457 = ~r1457;
  always #1125899906842624 r1458 = ~r1458;
  always #2251799813685248 r1459 = ~r1459;
  always #4503599627370496 r1460 = ~r1460;
  always #9007199254740992 r1461 = ~r1461;
  always #18014398509481984 r1462 = ~r1462;
  always #36028797018963968 r1463 = ~r1463;
  always #72057594037927936 r1464 = ~r1464;
  always #144115188075855872 r1465 = ~r1465;
  always #288230376151711744 r1466 = ~r1466;
  always #576460752303423488 r1467 = ~r1467;
  always #1152921504606846976 r1468 = ~r1468;
  always #2305843009213693952 r1469 = ~r1469;
  always #4611686018427387904 r1470 = ~r1470;
  always #9223372036854775808 r1471 = ~r1471;
  always #1 r1472 = ~r1472;
  always #2 r1473 = ~r1473;
  always #4 r1474 = ~r1474;
  always #8 r1475 = ~r1475;
  always #16 r1476 = ~r1476;
  always #32 r1477 = ~r1477;
  always #64 r1478 = ~r1478;
  always #128 r1479 = ~r1479;
  always #256 r1480 = ~r1480;
  always #512 r1481 = ~r1481;
  always #1024 r1482 = ~r1482;
  always #2048 r1483 = ~r1483;
  always #4096 r1484 = ~r1484;
  always #8192 r1485 = ~r1485;
  always #16384 r1486 = ~r1486;
  always #32768 r1487 = ~r1487;
  always #65536 r1488 = ~r1488;
  always #131072 r1489 = ~r1489;
  always #262144 r1490 = ~r1490;
  always #524288 r1491 = ~r1491;
  always #1048576 r1492 = ~r1492;
  always #2097152 r1493 = ~r1493;
  always #4194304 r1494 = ~r1494;
  always #8388608 r1495 = ~r1495;
  always #16777216 r1496 = ~r1496;
  always #33554432 r1497 = ~r1497;
  always #67108864 r1498 = ~r1498;
  always #134217728 r1499 = ~r1499;
  always #268435456 r1500 = ~r1500;
  always #536870912 r1501 = ~r1501;
  always #1073741824 r1502 = ~r1502;
  always #2147483648 r1503 = ~r1503;
  always #4294967296 r1504 = ~r1504;
  always #8589934592 r1505 = ~r1505;
  always #17179869184 r1506 = ~r1506;
  always #34359738368 r1507 = ~r1507;
  always #68719476736 r1508 = ~r1508;
  always #137438953472 r1509 = ~r1509;
  always #274877906944 r1510 = ~r1510;
  always #549755813888 r1511 = ~r1511;
  always #1099511627776 r1512 = ~r1512;
  always #2199023255552 r1513 = ~r1513;
  always #4398046511104 r1514 = ~r1514;
  always #8796093022208 r1515 = ~r1515;
  always #17592186044416 r1516 = ~r1516;
  always #35184372088832 r1517 = ~r1517;
  always #70368744177664 r1518 = ~r1518;
  always #140737488355328 r1519 = ~r1519;
  always #281474976710656 r1520 = ~r1520;
  always #562949953421312 r1521 = ~r1521;
  always #1125899906842624 r1522 = ~r1522;
  always #2251799813685248 r1523 = ~r1523;
  always #4503599627370496 r1524 = ~r1524;
  always #9007199254740992 r1525 = ~r1525;
  always #18014398509481984 r1526 = ~r1526;
  always #36028797018963968 r1527 = ~r1527;
  always #72057594037927936 r1528 = ~r1528;
  always #144115188075855872 r1529 = ~r1529;
  always #288230376151711744 r1530 = ~r1530;
  always #576460752303423488 r1531 = ~r1531;
  always #1152921504606846976 r1532 = ~r1532;
  always #2305843009213693952 r1533 = ~r1533;
  always #4611686018427387904 r1534 = ~r1534;
  always #9223372036854775808 r1535 = ~r1535;
  always #1 r1536 = ~r1536;
  always #2 r1537 = ~r1537;
  always #4 r1538 = ~r1538;
  always #8 r1539 = ~r1539;
  always #16 r1540 = ~r1540;
  always #32 r1541 = ~r1541;
  always #64 r1542 = ~r1542;
  always #128 r1543 = ~r1543;
  always #256 r1544 = ~r1544;
  always #512 r1545 = ~r1545;
  always #1024 r1546 = ~r1546;
  always #2048 r1547 = ~r1547;
  always #4096 r1548 = ~r1548;
  always #8192 r1549 = ~r1549;
  always #16384 r1550 = ~r1550;
  always #32768 r1551 = ~r1551;
  always #65536 r1552 = ~r1552;
  always #131072 r1553 = ~r1553;
  always #262144 r1554 = ~r1554;
  always #524288 r1555 = ~r1555;
  always #1048576 r1556 = ~r1556;
  always #2097152 r1557 = ~r1557;
  always #4194304 r1558 = ~r1558;
  always #8388608 r1559 = ~r1559;
  always #16777216 r1560 = ~r1560;
  always #33554432 r1561 = ~r1561;
  always #67108864 r1562 = ~r1562;
  always #134217728 r1563 = ~r1563;
  always #268435456 r1564 = ~r1564;
  always #536870912 r1565 = ~r1565;
  always #1073741824 r1566 = ~r1566;
  always #2147483648 r1567 = ~r1567;
  always #4294967296 r1568 = ~r1568;
  always #8589934592 r1569 = ~r1569;
  always #17179869184 r1570 = ~r1570;
  always #34359738368 r1571 = ~r1571;
  always #68719476736 r1572 = ~r1572;
  always #137438953472 r1573 = ~r1573;
  always #274877906944 r1574 = ~r1574;
  always #549755813888 r1575 = ~r1575;
  always #1099511627776 r1576 = ~r1576;
  always #2199023255552 r1577 = ~r1577;
  always #4398046511104 r1578 = ~r1578;
  always #8796093022208 r1579 = ~r1579;
  always #17592186044416 r1580 = ~r1580;
  always #35184372088832 r1581 = ~r1581;
  always #70368744177664 r1582 = ~r1582;
  always #140737488355328 r1583 = ~r1583;
  always #281474976710656 r1584 = ~r1584;
  always #562949953421312 r1585 = ~r1585;
  always #1125899906842624 r1586 = ~r1586;
  always #2251799813685248 r1587 = ~r1587;
  always #4503599627370496 r1588 = ~r1588;
  always #9007199254740992 r1589 = ~r1589;
  always #18014398509481984 r1590 = ~r1590;
  always #36028797018963968 r1591 = ~r1591;
  always #72057594037927936 r1592 = ~r1592;
  always #144115188075855872 r1593 = ~r1593;
  always #288230376151711744 r1594 = ~r1594;
  always #576460752303423488 r1595 = ~r1595;
  always #1152921504606846976 r1596 = ~r1596;
  always #2305843009213693952 r1597 = ~r1597;
  always #4611686018427387904 r1598 = ~r1598;
  always #9223372036854775808 r1599 = ~r1599;
  always #1 r1600 = ~r1600;
  always #2 r1601 = ~r1601;
  always #4 r1602 = ~r1602;
  always #8 r1603 = ~r1603;
  always #16 r1604 = ~r1604;
  always #32 r1605 = ~r1605;
  always #64 r1606 = ~r1606;
  always #128 r1607 = ~r1607;
  always #256 r1608 = ~r1608;
  always #512 r1609 = ~r1609;
  always #1024 r1610 = ~r1610;
  always #2048 r1611 = ~r1611;
  always #4096 r1612 = ~r1612;
  always #8192 r1613 = ~r1613;
  always #16384 r1614 = ~r1614;
  always #32768 r1615 = ~r1615;
  always #65536 r1616 = ~r1616;
  always #131072 r1617 = ~r1617;
  always #262144 r1618 = ~r1618;
  always #524288 r1619 = ~r1619;
  always #1048576 r1620 = ~r1620;
  always #2097152 r1621 = ~r1621;
  always #4194304 r1622 = ~r1622;
  always #8388608 r1623 = ~r1623;
  always #16777216 r1624 = ~r1624;
  always #33554432 r1625 = ~r1625;
  always #67108864 r1626 = ~r1626;
  always #134217728 r1627 = ~r1627;
  always #268435456 r1628 = ~r1628;
  always #536870912 r1629 = ~r1629;
  always #1073741824 r1630 = ~r1630;
  always #2147483648 r1631 = ~r1631;
  always #4294967296 r1632 = ~r1632;
  always #8589934592 r1633 = ~r1633;
  always #17179869184 r1634 = ~r1634;
  always #34359738368 r1635 = ~r1635;
  always #68719476736 r1636 = ~r1636;
  always #137438953472 r1637 = ~r1637;
  always #274877906944 r1638 = ~r1638;
  always #549755813888 r1639 = ~r1639;
  always #1099511627776 r1640 = ~r1640;
  always #2199023255552 r1641 = ~r1641;
  always #4398046511104 r1642 = ~r1642;
  always #8796093022208 r1643 = ~r1643;
  always #17592186044416 r1644 = ~r1644;
  always #35184372088832 r1645 = ~r1645;
  always #70368744177664 r1646 = ~r1646;
  always #140737488355328 r1647 = ~r1647;
  always #281474976710656 r1648 = ~r1648;
  always #562949953421312 r1649 = ~r1649;
  always #1125899906842624 r1650 = ~r1650;
  always #2251799813685248 r1651 = ~r1651;
  always #4503599627370496 r1652 = ~r1652;
  always #9007199254740992 r1653 = ~r1653;
  always #18014398509481984 r1654 = ~r1654;
  always #36028797018963968 r1655 = ~r1655;
  always #72057594037927936 r1656 = ~r1656;
  always #144115188075855872 r1657 = ~r1657;
  always #288230376151711744 r1658 = ~r1658;
  always #576460752303423488 r1659 = ~r1659;
  always #1152921504606846976 r1660 = ~r1660;
  always #2305843009213693952 r1661 = ~r1661;
  always #4611686018427387904 r1662 = ~r1662;
  always #9223372036854775808 r1663 = ~r1663;
  always #1 r1664 = ~r1664;
  always #2 r1665 = ~r1665;
  always #4 r1666 = ~r1666;
  always #8 r1667 = ~r1667;
  always #16 r1668 = ~r1668;
  always #32 r1669 = ~r1669;
  always #64 r1670 = ~r1670;
  always #128 r1671 = ~r1671;
  always #256 r1672 = ~r1672;
  always #512 r1673 = ~r1673;
  always #1024 r1674 = ~r1674;
  always #2048 r1675 = ~r1675;
  always #4096 r1676 = ~r1676;
  always #8192 r1677 = ~r1677;
  always #16384 r1678 = ~r1678;
  always #32768 r1679 = ~r1679;
  always #65536 r1680 = ~r1680;
  always #131072 r1681 = ~r1681;
  always #262144 r1682 = ~r1682;
  always #524288 r1683 = ~r1683;
  always #1048576 r1684 = ~r1684;
  always #2097152 r1685 = ~r1685;
  always #4194304 r1686 = ~r1686;
  always #8388608 r1687 = ~r1687;
  always #16777216 r1688 = ~r1688;
  always #33554432 r1689 = ~r1689;
  always #67108864 r1690 = ~r1690;
  always #134217728 r1691 = ~r1691;
  always #268435456 r1692 = ~r1692;
  always #536870912 r1693 = ~r1693;
  always #1073741824 r1694 = ~r1694;
  always #2147483648 r1695 = ~r1695;
  always #4294967296 r1696 = ~r1696;
  always #8589934592 r1697 = ~r1697;
  always #17179869184 r1698 = ~r1698;
  always #34359738368 r1699 = ~r1699;
  always #68719476736 r1700 = ~r1700;
  always #137438953472 r1701 = ~r1701;
  always #274877906944 r1702 = ~r1702;
  always #549755813888 r1703 = ~r1703;
  always #1099511627776 r1704 = ~r1704;
  always #2199023255552 r1705 = ~r1705;
  always #4398046511104 r1706 = ~r1706;
  always #8796093022208 r1707 = ~r1707;
  always #17592186044416 r1708 = ~r1708;
  always #35184372088832 r1709 = ~r1709;
  always #70368744177664 r1710 = ~r1710;
  always #140737488355328 r1711 = ~r1711;
  always #281474976710656 r1712 = ~r1712;
  always #562949953421312 r1713 = ~r1713;
  always #1125899906842624 r1714 = ~r1714;
  always #2251799813685248 r1715 = ~r1715;
  always #4503599627370496 r1716 = ~r1716;
  always #9007199254740992 r1717 = ~r1717;
  always #18014398509481984 r1718 = ~r1718;
  always #36028797018963968 r1719 = ~r1719;
  always #72057594037927936 r1720 = ~r1720;
  always #144115188075855872 r1721 = ~r1721;
  always #288230376151711744 r1722 = ~r1722;
  always #576460752303423488 r1723 = ~r1723;
  always #1152921504606846976 r1724 = ~r1724;
  always #2305843009213693952 r1725 = ~r1725;
  always #4611686018427387904 r1726 = ~r1726;
  always #9223372036854775808 r1727 = ~r1727;
  always #1 r1728 = ~r1728;
  always #2 r1729 = ~r1729;
  always #4 r1730 = ~r1730;
  always #8 r1731 = ~r1731;
  always #16 r1732 = ~r1732;
  always #32 r1733 = ~r1733;
  always #64 r1734 = ~r1734;
  always #128 r1735 = ~r1735;
  always #256 r1736 = ~r1736;
  always #512 r1737 = ~r1737;
  always #1024 r1738 = ~r1738;
  always #2048 r1739 = ~r1739;
  always #4096 r1740 = ~r1740;
  always #8192 r1741 = ~r1741;
  always #16384 r1742 = ~r1742;
  always #32768 r1743 = ~r1743;
  always #65536 r1744 = ~r1744;
  always #131072 r1745 = ~r1745;
  always #262144 r1746 = ~r1746;
  always #524288 r1747 = ~r1747;
  always #1048576 r1748 = ~r1748;
  always #2097152 r1749 = ~r1749;
  always #4194304 r1750 = ~r1750;
  always #8388608 r1751 = ~r1751;
  always #16777216 r1752 = ~r1752;
  always #33554432 r1753 = ~r1753;
  always #67108864 r1754 = ~r1754;
  always #134217728 r1755 = ~r1755;
  always #268435456 r1756 = ~r1756;
  always #536870912 r1757 = ~r1757;
  always #1073741824 r1758 = ~r1758;
  always #2147483648 r1759 = ~r1759;
  always #4294967296 r1760 = ~r1760;
  always #8589934592 r1761 = ~r1761;
  always #17179869184 r1762 = ~r1762;
  always #34359738368 r1763 = ~r1763;
  always #68719476736 r1764 = ~r1764;
  always #137438953472 r1765 = ~r1765;
  always #274877906944 r1766 = ~r1766;
  always #549755813888 r1767 = ~r1767;
  always #1099511627776 r1768 = ~r1768;
  always #2199023255552 r1769 = ~r1769;
  always #4398046511104 r1770 = ~r1770;
  always #8796093022208 r1771 = ~r1771;
  always #17592186044416 r1772 = ~r1772;
  always #35184372088832 r1773 = ~r1773;
  always #70368744177664 r1774 = ~r1774;
  always #140737488355328 r1775 = ~r1775;
  always #281474976710656 r1776 = ~r1776;
  always #562949953421312 r1777 = ~r1777;
  always #1125899906842624 r1778 = ~r1778;
  always #2251799813685248 r1779 = ~r1779;
  always #4503599627370496 r1780 = ~r1780;
  always #9007199254740992 r1781 = ~r1781;
  always #18014398509481984 r1782 = ~r1782;
  always #36028797018963968 r1783 = ~r1783;
  always #72057594037927936 r1784 = ~r1784;
  always #144115188075855872 r1785 = ~r1785;
  always #288230376151711744 r1786 = ~r1786;
  always #576460752303423488 r1787 = ~r1787;
  always #1152921504606846976 r1788 = ~r1788;
  always #2305843009213693952 r1789 = ~r1789;
  always #4611686018427387904 r1790 = ~r1790;
  always #9223372036854775808 r1791 = ~r1791;
  always #1 r1792 = ~r1792;
  always #2 r1793 = ~r1793;
  always #4 r1794 = ~r1794;
  always #8 r1795 = ~r1795;
  always #16 r1796 = ~r1796;
  always #32 r1797 = ~r1797;
  always #64 r1798 = ~r1798;
  always #128 r1799 = ~r1799;
  always #256 r1800 = ~r1800;
  always #512 r1801 = ~r1801;
  always #1024 r1802 = ~r1802;
  always #2048 r1803 = ~r1803;
  always #4096 r1804 = ~r1804;
  always #8192 r1805 = ~r1805;
  always #16384 r1806 = ~r1806;
  always #32768 r1807 = ~r1807;
  always #65536 r1808 = ~r1808;
  always #131072 r1809 = ~r1809;
  always #262144 r1810 = ~r1810;
  always #524288 r1811 = ~r1811;
  always #1048576 r1812 = ~r1812;
  always #2097152 r1813 = ~r1813;
  always #4194304 r1814 = ~r1814;
  always #8388608 r1815 = ~r1815;
  always #16777216 r1816 = ~r1816;
  always #33554432 r1817 = ~r1817;
  always #67108864 r1818 = ~r1818;
  always #134217728 r1819 = ~r1819;
  always #268435456 r1820 = ~r1820;
  always #536870912 r1821 = ~r1821;
  always #1073741824 r1822 = ~r1822;
  always #2147483648 r1823 = ~r1823;
  always #4294967296 r1824 = ~r1824;
  always #8589934592 r1825 = ~r1825;
  always #17179869184 r1826 = ~r1826;
  always #34359738368 r1827 = ~r1827;
  always #68719476736 r1828 = ~r1828;
  always #137438953472 r1829 = ~r1829;
  always #274877906944 r1830 = ~r1830;
  always #549755813888 r1831 = ~r1831;
  always #1099511627776 r1832 = ~r1832;
  always #2199023255552 r1833 = ~r1833;
  always #4398046511104 r1834 = ~r1834;
  always #8796093022208 r1835 = ~r1835;
  always #17592186044416 r1836 = ~r1836;
  always #35184372088832 r1837 = ~r1837;
  always #70368744177664 r1838 = ~r1838;
  always #140737488355328 r1839 = ~r1839;
  always #281474976710656 r1840 = ~r1840;
  always #562949953421312 r1841 = ~r1841;
  always #1125899906842624 r1842 = ~r1842;
  always #2251799813685248 r1843 = ~r1843;
  always #4503599627370496 r1844 = ~r1844;
  always #9007199254740992 r1845 = ~r1845;
  always #18014398509481984 r1846 = ~r1846;
  always #36028797018963968 r1847 = ~r1847;
  always #72057594037927936 r1848 = ~r1848;
  always #144115188075855872 r1849 = ~r1849;
  always #288230376151711744 r1850 = ~r1850;
  always #576460752303423488 r1851 = ~r1851;
  always #1152921504606846976 r1852 = ~r1852;
  always #2305843009213693952 r1853 = ~r1853;
  always #4611686018427387904 r1854 = ~r1854;
  always #9223372036854775808 r1855 = ~r1855;
  always #1 r1856 = ~r1856;
  always #2 r1857 = ~r1857;
  always #4 r1858 = ~r1858;
  always #8 r1859 = ~r1859;
  always #16 r1860 = ~r1860;
  always #32 r1861 = ~r1861;
  always #64 r1862 = ~r1862;
  always #128 r1863 = ~r1863;
  always #256 r1864 = ~r1864;
  always #512 r1865 = ~r1865;
  always #1024 r1866 = ~r1866;
  always #2048 r1867 = ~r1867;
  always #4096 r1868 = ~r1868;
  always #8192 r1869 = ~r1869;
  always #16384 r1870 = ~r1870;
  always #32768 r1871 = ~r1871;
  always #65536 r1872 = ~r1872;
  always #131072 r1873 = ~r1873;
  always #262144 r1874 = ~r1874;
  always #524288 r1875 = ~r1875;
  always #1048576 r1876 = ~r1876;
  always #2097152 r1877 = ~r1877;
  always #4194304 r1878 = ~r1878;
  always #8388608 r1879 = ~r1879;
  always #16777216 r1880 = ~r1880;
  always #33554432 r1881 = ~r1881;
  always #67108864 r1882 = ~r1882;
  always #134217728 r1883 = ~r1883;
  always #268435456 r1884 = ~r1884;
  always #536870912 r1885 = ~r1885;
  always #1073741824 r1886 = ~r1886;
  always #2147483648 r1887 = ~r1887;
  always #4294967296 r1888 = ~r1888;
  always #8589934592 r1889 = ~r1889;
  always #17179869184 r1890 = ~r1890;
  always #34359738368 r1891 = ~r1891;
  always #68719476736 r1892 = ~r1892;
  always #137438953472 r1893 = ~r1893;
  always #274877906944 r1894 = ~r1894;
  always #549755813888 r1895 = ~r1895;
  always #1099511627776 r1896 = ~r1896;
  always #2199023255552 r1897 = ~r1897;
  always #4398046511104 r1898 = ~r1898;
  always #8796093022208 r1899 = ~r1899;
  always #17592186044416 r1900 = ~r1900;
  always #35184372088832 r1901 = ~r1901;
  always #70368744177664 r1902 = ~r1902;
  always #140737488355328 r1903 = ~r1903;
  always #281474976710656 r1904 = ~r1904;
  always #562949953421312 r1905 = ~r1905;
  always #1125899906842624 r1906 = ~r1906;
  always #2251799813685248 r1907 = ~r1907;
  always #4503599627370496 r1908 = ~r1908;
  always #9007199254740992 r1909 = ~r1909;
  always #18014398509481984 r1910 = ~r1910;
  always #36028797018963968 r1911 = ~r1911;
  always #72057594037927936 r1912 = ~r1912;
  always #144115188075855872 r1913 = ~r1913;
  always #288230376151711744 r1914 = ~r1914;
  always #576460752303423488 r1915 = ~r1915;
  always #1152921504606846976 r1916 = ~r1916;
  always #2305843009213693952 r1917 = ~r1917;
  always #4611686018427387904 r1918 = ~r1918;
  always #9223372036854775808 r1919 = ~r1919;
  always #1 r1920 = ~r1920;
  always #2 r1921 = ~r1921;
  always #4 r1922 = ~r1922;
  always #8 r1923 = ~r1923;
  always #16 r1924 = ~r1924;
  always #32 r1925 = ~r1925;
  always #64 r1926 = ~r1926;
  always #128 r1927 = ~r1927;
  always #256 r1928 = ~r1928;
  always #512 r1929 = ~r1929;
  always #1024 r1930 = ~r1930;
  always #2048 r1931 = ~r1931;
  always #4096 r1932 = ~r1932;
  always #8192 r1933 = ~r1933;
  always #16384 r1934 = ~r1934;
  always #32768 r1935 = ~r1935;
  always #65536 r1936 = ~r1936;
  always #131072 r1937 = ~r1937;
  always #262144 r1938 = ~r1938;
  always #524288 r1939 = ~r1939;
  always #1048576 r1940 = ~r1940;
  always #2097152 r1941 = ~r1941;
  always #4194304 r1942 = ~r1942;
  always #8388608 r1943 = ~r1943;
  always #16777216 r1944 = ~r1944;
  always #33554432 r1945 = ~r1945;
  always #67108864 r1946 = ~r1946;
  always #134217728 r1947 = ~r1947;
  always #268435456 r1948 = ~r1948;
  always #536870912 r1949 = ~r1949;
  always #1073741824 r1950 = ~r1950;
  always #2147483648 r1951 = ~r1951;
  always #4294967296 r1952 = ~r1952;
  always #8589934592 r1953 = ~r1953;
  always #17179869184 r1954 = ~r1954;
  always #34359738368 r1955 = ~r1955;
  always #68719476736 r1956 = ~r1956;
  always #137438953472 r1957 = ~r1957;
  always #274877906944 r1958 = ~r1958;
  always #549755813888 r1959 = ~r1959;
  always #1099511627776 r1960 = ~r1960;
  always #2199023255552 r1961 = ~r1961;
  always #4398046511104 r1962 = ~r1962;
  always #8796093022208 r1963 = ~r1963;
  always #17592186044416 r1964 = ~r1964;
  always #35184372088832 r1965 = ~r1965;
  always #70368744177664 r1966 = ~r1966;
  always #140737488355328 r1967 = ~r1967;
  always #281474976710656 r1968 = ~r1968;
  always #562949953421312 r1969 = ~r1969;
  always #1125899906842624 r1970 = ~r1970;
  always #2251799813685248 r1971 = ~r1971;
  always #4503599627370496 r1972 = ~r1972;
  always #9007199254740992 r1973 = ~r1973;
  always #18014398509481984 r1974 = ~r1974;
  always #36028797018963968 r1975 = ~r1975;
  always #72057594037927936 r1976 = ~r1976;
  always #144115188075855872 r1977 = ~r1977;
  always #288230376151711744 r1978 = ~r1978;
  always #576460752303423488 r1979 = ~r1979;
  always #1152921504606846976 r1980 = ~r1980;
  always #2305843009213693952 r1981 = ~r1981;
  always #4611686018427387904 r1982 = ~r1982;
  always #9223372036854775808 r1983 = ~r1983;
  always #1 r1984 = ~r1984;
  always #2 r1985 = ~r1985;
  always #4 r1986 = ~r1986;
  always #8 r1987 = ~r1987;
  always #16 r1988 = ~r1988;
  always #32 r1989 = ~r1989;
  always #64 r1990 = ~r1990;
  always #128 r1991 = ~r1991;
  always #256 r1992 = ~r1992;
  always #512 r1993 = ~r1993;
  always #1024 r1994 = ~r1994;
  always #2048 r1995 = ~r1995;
  always #4096 r1996 = ~r1996;
  always #8192 r1997 = ~r1997;
endmodule
*/
// ****** TestBench Module Defination End ******

/*
// ******* The results for this case *********
******* result_1.txt *********
1)
  Loop Signals: w_894_586, w_894_587, w_894_588, w_894_589, w_894_590, w_894_591, 
  Loop Gates: I894_585.port1, I894_586.port2, I894_587.port2, I894_588.port2, I894_589.port1, I894_590.port1, 

2)
  Loop Signals: w_894_586, w_894_595, w_894_596, w_894_597, w_894_598, w_894_599, w_894_600, w_894_601, w_894_602, w_894_603, w_894_604, w_894_605, w_894_607, 
  Loop Gates: I894_590.port2, I894_591.port1, I894_592.port1, I894_593.port1, I894_594.port1, I894_595.port2, I894_596.port1, I894_597.port1, I894_598.port2, I894_599.port2, I894_600.port1, I894_601.port1, I894_602.port2, 

3)
  Loop Signals: w_102_1259, w_102_1260, w_102_1261, w_102_1262, w_102_1263, w_102_1264, 
  Loop Gates: I102_1258.port1, I102_1259.port2, I102_1260.port2, I102_1261.port2, I102_1262.port1, I102_1263.port1, 

4)
  Loop Signals: w_102_1259, w_102_1268, w_102_1269, w_102_1270, w_102_1271, w_102_1272, w_102_1273, w_102_1274, w_102_1275, w_102_1276, w_102_1278, 
  Loop Gates: I102_1263.port2, I102_1264.port1, I102_1265.port1, I102_1266.port2, I102_1267.port2, I102_1268.port2, I102_1269.port1, I102_1270.port2, I102_1271.port1, I102_1272.port1, I102_1273.port2, 

5)
  Loop Signals: w_054_628, w_054_629, w_054_630, w_054_631, w_054_632, w_054_633, w_054_634, w_054_635, w_054_636, w_054_637, 
  Loop Gates: I054_627.port2, I054_628.port1, I054_629.port1, I054_630.port2, I054_631.port1, I054_632.port1, I054_633.port1, I054_634.port2, I054_635.port1, I054_636.port2, 

6)
  Loop Signals: w_457_1221, w_457_1222, w_457_1223, w_457_1224, w_457_1225, w_457_1226, 
  Loop Gates: I457_1220.port2, I457_1221.port1, I457_1222.port1, I457_1223.port2, I457_1224.port1, I457_1225.port1, 

7)
  Loop Signals: w_484_492, w_484_493, w_484_494, 
  Loop Gates: I484_491.port1, I484_492.port1, I484_493.port1, 

8)
  Loop Signals: w_484_492, w_484_498, w_484_499, w_484_500, w_484_501, w_484_502, w_484_503, w_484_504, w_484_505, w_484_506, w_484_507, w_484_509, 
  Loop Gates: I484_493.port2, I484_494.port1, I484_495.port1, I484_496.port2, I484_497.port1, I484_498.port1, I484_499.port1, I484_500.port2, I484_501.port1, I484_502.port1, I484_503.port1, I484_504.port2, 

9)
  Loop Signals: w_1818_359, w_1818_360, w_1818_361, w_1818_362, 
  Loop Gates: I1818_358.port1, I1818_359.port2, I1818_360.port1, I1818_361.port1, 

10)
  Loop Signals: w_799_848, w_799_849, w_799_850, w_799_851, w_799_852, w_799_853, w_799_854, w_799_855, w_799_856, 
  Loop Gates: I799_847.port1, I799_848.port2, I799_849.port2, I799_850.port1, I799_851.port1, I799_852.port1, I799_853.port1, I799_854.port1, I799_855.port2, 

11)
  Loop Signals: w_799_855, w_799_860, w_799_861, w_799_862, w_799_863, w_799_865, 
  Loop Gates: I799_853.port2, I799_856.port1, I799_857.port1, I799_858.port1, I799_859.port1, I799_860.port2, 

12)
  Loop Signals: w_235_1042, w_235_1043, w_235_1044, w_235_1045, w_235_1046, w_235_1047, w_235_1048, 
  Loop Gates: I235_1041.port2, I235_1042.port2, I235_1043.port1, I235_1044.port2, I235_1045.port1, I235_1046.port1, I235_1047.port1, 

13)
  Loop Signals: w_235_1047, w_235_1052, w_235_1053, w_235_1054, w_235_1055, w_235_1056, w_235_1057, w_235_1058, w_235_1059, w_235_1060, w_235_1062, 
  Loop Gates: I235_1045.port2, I235_1048.port2, I235_1049.port2, I235_1050.port1, I235_1051.port1, I235_1052.port2, I235_1053.port2, I235_1054.port1, I235_1055.port1, I235_1056.port1, I235_1057.port2, 

14)
  Loop Signals: w_811_1656, w_811_1657, w_811_1658, 
  Loop Gates: I811_1655.port1, I811_1656.port1, I811_1657.port2, 

15)
  Loop Signals: w_811_1656, w_811_1662, w_811_1663, w_811_1664, w_811_1665, w_811_1666, w_811_1667, w_811_1668, w_811_1670, 
  Loop Gates: I811_1657.port1, I811_1658.port1, I811_1659.port1, I811_1660.port1, I811_1661.port2, I811_1662.port1, I811_1663.port1, I811_1664.port1, I811_1665.port2, 

16)
  Loop Signals: w_432_726, w_432_727, w_432_728, w_432_729, w_432_730, w_432_731, 
  Loop Gates: I432_725.port1, I432_726.port2, I432_727.port1, I432_728.port1, I432_729.port2, I432_730.port1, 

17)
  Loop Signals: w_432_726, w_432_735, w_432_736, w_432_737, w_432_738, w_432_739, w_432_741, 
  Loop Gates: I432_730.port2, I432_731.port2, I432_732.port2, I432_733.port2, I432_734.port1, I432_735.port1, I432_736.port2, 

18)
  Loop Signals: w_769_203, w_769_204, w_769_205, w_769_206, w_769_207, w_769_208, w_769_209, 
  Loop Gates: I769_202.port2, I769_203.port2, I769_204.port1, I769_205.port1, I769_206.port1, I769_207.port2, I769_208.port1, 

19)
  Loop Signals: w_1656_1927, w_1656_1928, w_1656_1929, w_1656_1930, 
  Loop Gates: I1656_1926.port2, I1656_1927.port1, I1656_1928.port1, I1656_1929.port1, 

20)
  Loop Signals: w_1692_766, w_1692_767, w_1692_768, w_1692_769, w_1692_770, 
  Loop Gates: I1692_765.port1, I1692_766.port1, I1692_767.port2, I1692_768.port1, I1692_769.port1, 

21)
  Loop Signals: w_1692_769, w_1692_774, w_1692_775, w_1692_776, w_1692_777, w_1692_778, w_1692_779, w_1692_780, w_1692_782, 
  Loop Gates: I1692_767.port1, I1692_770.port1, I1692_771.port2, I1692_772.port1, I1692_773.port2, I1692_774.port1, I1692_775.port1, I1692_776.port1, I1692_777.port2, 

22)
  Loop Signals: w_1298_518, w_1298_519, w_1298_520, 
  Loop Gates: I1298_517.port1, I1298_518.port2, I1298_519.port2, 

23)
  Loop Signals: w_1298_518, w_1298_524, w_1298_525, w_1298_526, w_1298_527, w_1298_529, 
  Loop Gates: I1298_519.port1, I1298_520.port1, I1298_521.port2, I1298_522.port1, I1298_523.port1, I1298_524.port2, 

24)
  Loop Signals: w_494_1931, w_494_1932, w_494_1933, w_494_1934, w_494_1935, w_494_1936, 
  Loop Gates: I494_1930.port1, I494_1931.port2, I494_1932.port2, I494_1933.port2, I494_1934.port2, I494_1935.port1, 

25)
  Loop Signals: w_563_960, w_563_961, w_563_962, w_563_963, 
  Loop Gates: I563_959.port1, I563_960.port1, I563_961.port2, I563_962.port2, 

26)
  Loop Signals: w_610_889, w_610_890, w_610_891, w_610_892, w_610_893, w_610_894, w_610_895, w_610_896, w_610_897, w_610_898, w_610_899, 
  Loop Gates: I610_888.port1, I610_889.port1, I610_890.port1, I610_891.port1, I610_892.port1, I610_893.port1, I610_894.port2, I610_895.port1, I610_896.port1, I610_897.port2, I610_898.port1, 

27)
  Loop Signals: w_1230_965, w_1230_966, w_1230_967, w_1230_968, w_1230_969, w_1230_970, 
  Loop Gates: I1230_964.port2, I1230_965.port1, I1230_966.port1, I1230_967.port1, I1230_968.port2, I1230_969.port1, 

28)
  Loop Signals: w_342_1768, w_342_1769, w_342_1770, w_342_1771, w_342_1772, w_342_1773, w_342_1774, w_342_1775, w_342_1776, w_342_1777, 
  Loop Gates: I342_1767.port2, I342_1768.port2, I342_1769.port1, I342_1770.port1, I342_1771.port2, I342_1772.port2, I342_1773.port1, I342_1774.port2, I342_1775.port2, I342_1776.port1, 

29)
  Loop Signals: w_342_1775, w_342_1781, w_342_1782, w_342_1783, w_342_1784, w_342_1785, w_342_1786, w_342_1788, 
  Loop Gates: I342_1773.port2, I342_1777.port2, I342_1778.port1, I342_1779.port1, I342_1780.port2, I342_1781.port2, I342_1782.port1, I342_1783.port2, 

30)
  Loop Signals: w_1288_1602, w_1288_1603, w_1288_1604, w_1288_1605, w_1288_1606, w_1288_1607, 
  Loop Gates: I1288_1601.port1, I1288_1602.port1, I1288_1603.port2, I1288_1604.port1, I1288_1605.port1, I1288_1606.port1, 

31)
  Loop Signals: w_1288_1604, w_1288_1611, w_1288_1612, w_1288_1613, w_1288_1614, w_1288_1615, w_1288_1616, w_1288_1617, w_1288_1618, w_1288_1619, w_1288_1620, w_1288_1622, 
  Loop Gates: I1288_1602.port2, I1288_1607.port2, I1288_1608.port1, I1288_1609.port1, I1288_1610.port1, I1288_1611.port1, I1288_1612.port1, I1288_1613.port1, I1288_1614.port2, I1288_1615.port2, I1288_1616.port1, I1288_1617.port2, 

32)
  Loop Signals: w_009_113, w_009_114, w_009_115, w_009_116, w_009_117, w_009_118, w_009_119, w_009_120, 
  Loop Gates: I009_112.port2, I009_113.port1, I009_114.port1, I009_115.port1, I009_116.port2, I009_117.port2, I009_118.port1, I009_119.port1, 

33)
  Loop Signals: w_009_118, w_009_124, w_009_125, w_009_126, w_009_127, w_009_128, w_009_129, w_009_131, 
  Loop Gates: I009_116.port1, I009_120.port1, I009_121.port1, I009_122.port2, I009_123.port1, I009_124.port1, I009_125.port1, I009_126.port2, 

34)
  Loop Signals: w_826_437, w_826_438, w_826_439, w_826_440, 
  Loop Gates: I826_436.port1, I826_437.port1, I826_438.port1, I826_439.port1, 

35)
  Loop Signals: w_826_440, w_826_444, w_826_445, w_826_446, w_826_447, w_826_448, w_826_449, w_826_450, w_826_452, 
  Loop Gates: I826_438.port2, I826_440.port1, I826_441.port1, I826_442.port2, I826_443.port1, I826_444.port1, I826_445.port1, I826_446.port1, I826_447.port2, 

36)
  Loop Signals: w_1132_1117, w_1132_1118, w_1132_1119, w_1132_1120, w_1132_1121, w_1132_1122, w_1132_1123, 
  Loop Gates: I1132_1116.port1, I1132_1117.port1, I1132_1118.port1, I1132_1119.port2, I1132_1120.port1, I1132_1121.port2, I1132_1122.port2, 

37)
  Loop Signals: w_1449_506, w_1449_507, w_1449_508, w_1449_509, 
  Loop Gates: I1449_505.port2, I1449_506.port2, I1449_507.port2, I1449_508.port1, 

38)
  Loop Signals: w_1423_462, w_1423_463, w_1423_464, w_1423_465, w_1423_466, w_1423_467, w_1423_468, w_1423_469, w_1423_470, w_1423_471, w_1423_472, 
  Loop Gates: I1423_461.port1, I1423_462.port1, I1423_463.port2, I1423_464.port1, I1423_465.port1, I1423_466.port2, I1423_467.port1, I1423_468.port2, I1423_469.port2, I1423_470.port1, I1423_471.port1, 

39)
  Loop Signals: w_1308_361, w_1308_362, w_1308_363, w_1308_364, w_1308_365, w_1308_366, w_1308_367, w_1308_368, w_1308_369, w_1308_370, w_1308_371, w_1308_372, 
  Loop Gates: I1308_360.port1, I1308_361.port1, I1308_362.port1, I1308_363.port1, I1308_364.port1, I1308_365.port1, I1308_366.port1, I1308_367.port1, I1308_368.port1, I1308_369.port1, I1308_370.port1, I1308_371.port1, 

40)
  Loop Signals: w_1308_362, w_1308_376, w_1308_377, w_1308_378, w_1308_379, w_1308_380, w_1308_381, w_1308_382, w_1308_384, 
  Loop Gates: I1308_360.port2, I1308_372.port1, I1308_373.port1, I1308_374.port2, I1308_375.port1, I1308_376.port1, I1308_377.port2, I1308_378.port1, I1308_379.port2, 

41)
  Loop Signals: w_531_1378, w_531_1379, w_531_1380, w_531_1381, w_531_1382, w_531_1383, w_531_1384, w_531_1385, w_531_1386, w_531_1387, w_531_1388, 
  Loop Gates: I531_1377.port1, I531_1378.port1, I531_1379.port1, I531_1380.port1, I531_1381.port1, I531_1382.port1, I531_1383.port1, I531_1384.port1, I531_1385.port1, I531_1386.port2, I531_1387.port1, 

42)
  Loop Signals: w_531_1388, w_531_1392, w_531_1393, w_531_1394, w_531_1395, w_531_1397, 
  Loop Gates: I531_1386.port1, I531_1388.port1, I531_1389.port2, I531_1390.port1, I531_1391.port1, I531_1392.port2, 

43)
  Loop Signals: w_1821_248, w_1821_249, w_1821_250, w_1821_251, w_1821_252, w_1821_253, 
  Loop Gates: I1821_247.port2, I1821_248.port2, I1821_249.port1, I1821_250.port1, I1821_251.port2, I1821_252.port1, 

44)
  Loop Signals: w_1821_251, w_1821_257, w_1821_258, w_1821_259, w_1821_260, w_1821_261, w_1821_262, w_1821_263, w_1821_264, w_1821_265, w_1821_266, w_1821_268, 
  Loop Gates: I1821_249.port2, I1821_253.port1, I1821_254.port1, I1821_255.port2, I1821_256.port2, I1821_257.port1, I1821_258.port1, I1821_259.port1, I1821_260.port2, I1821_261.port1, I1821_262.port1, I1821_263.port2, 

45)
  Loop Signals: w_1601_113, w_1601_114, w_1601_115, 
  Loop Gates: I1601_112.port1, I1601_113.port2, I1601_114.port1, 

46)
  Loop Signals: w_1601_115, w_1601_119, w_1601_120, w_1601_121, w_1601_122, w_1601_123, w_1601_124, w_1601_125, w_1601_127, 
  Loop Gates: I1601_113.port1, I1601_115.port1, I1601_116.port1, I1601_117.port1, I1601_118.port1, I1601_119.port1, I1601_120.port1, I1601_121.port1, I1601_122.port2, 

47)
  Loop Signals: w_1848_117, w_1848_118, w_1848_119, w_1848_120, 
  Loop Gates: I1848_116.port1, I1848_117.port1, I1848_118.port1, I1848_119.port1, 

48)
  Loop Signals: w_305_018, w_305_019, w_305_020, w_305_021, w_305_022, w_305_023, w_305_024, 
  Loop Gates: I305_017.port2, I305_018.port1, I305_019.port2, I305_020.port1, I305_021.port1, I305_022.port2, I305_023.port2, 

49)
  Loop Signals: w_1836_1757, w_1836_1758, w_1836_1759, w_1836_1760, w_1836_1761, w_1836_1762, w_1836_1763, w_1836_1764, w_1836_1765, w_1836_1766, w_1836_1767, w_1836_1768, 
  Loop Gates: I1836_1756.port1, I1836_1757.port2, I1836_1758.port1, I1836_1759.port2, I1836_1760.port1, I1836_1761.port1, I1836_1762.port1, I1836_1763.port1, I1836_1764.port2, I1836_1765.port1, I1836_1766.port2, I1836_1767.port1, 

50)
  Loop Signals: w_1836_1768, w_1836_1772, w_1836_1773, w_1836_1774, w_1836_1775, w_1836_1776, w_1836_1778, 
  Loop Gates: I1836_1766.port1, I1836_1768.port1, I1836_1769.port2, I1836_1770.port1, I1836_1771.port2, I1836_1772.port1, I1836_1773.port2, 

51)
  Loop Signals: w_1911_1096, w_1911_1097, w_1911_1098, w_1911_1099, w_1911_1100, w_1911_1101, w_1911_1102, w_1911_1103, w_1911_1104, w_1911_1105, w_1911_1106, w_1911_1107, 
  Loop Gates: I1911_1095.port1, I1911_1096.port1, I1911_1097.port2, I1911_1098.port2, I1911_1099.port1, I1911_1100.port1, I1911_1101.port1, I1911_1102.port1, I1911_1103.port2, I1911_1104.port2, I1911_1105.port1, I1911_1106.port2, 

52)
  Loop Signals: w_1579_1708, w_1579_1709, w_1579_1710, w_1579_1711, w_1579_1712, w_1579_1713, w_1579_1714, w_1579_1715, 
  Loop Gates: I1579_1707.port1, I1579_1708.port1, I1579_1709.port1, I1579_1710.port1, I1579_1711.port1, I1579_1712.port2, I1579_1713.port1, I1579_1714.port1, 

53)
  Loop Signals: w_851_1288, w_851_1289, w_851_1290, w_851_1291, w_851_1292, w_851_1293, w_851_1294, w_851_1295, w_851_1296, w_851_1297, 
  Loop Gates: I851_1287.port1, I851_1288.port1, I851_1289.port2, I851_1290.port1, I851_1291.port1, I851_1292.port1, I851_1293.port1, I851_1294.port1, I851_1295.port1, I851_1296.port1, 

54)
  Loop Signals: w_1176_1251, w_1176_1252, w_1176_1253, w_1176_1254, w_1176_1255, w_1176_1256, w_1176_1257, w_1176_1258, w_1176_1259, w_1176_1260, w_1176_1261, w_1176_1262, 
  Loop Gates: I1176_1250.port2, I1176_1251.port1, I1176_1252.port1, I1176_1253.port2, I1176_1254.port2, I1176_1255.port1, I1176_1256.port1, I1176_1257.port2, I1176_1258.port1, I1176_1259.port2, I1176_1260.port2, I1176_1261.port1, 

55)
  Loop Signals: w_299_1759, w_299_1760, w_299_1761, 
  Loop Gates: I299_1758.port1, I299_1759.port2, I299_1760.port1, 

56)
  Loop Signals: w_1075_1904, w_1075_1905, w_1075_1906, w_1075_1907, w_1075_1908, w_1075_1909, w_1075_1910, w_1075_1911, 
  Loop Gates: I1075_1903.port1, I1075_1904.port1, I1075_1905.port2, I1075_1906.port2, I1075_1907.port1, I1075_1908.port2, I1075_1909.port1, I1075_1910.port1, 

57)
  Loop Signals: w_1075_1910, w_1075_1915, w_1075_1916, w_1075_1917, w_1075_1918, w_1075_1919, w_1075_1920, w_1075_1921, w_1075_1922, w_1075_1924, 
  Loop Gates: I1075_1908.port1, I1075_1911.port2, I1075_1912.port1, I1075_1913.port2, I1075_1914.port2, I1075_1915.port1, I1075_1916.port1, I1075_1917.port2, I1075_1918.port1, I1075_1919.port2, 

58)
  Loop Signals: w_919_1871, w_919_1872, w_919_1873, w_919_1874, w_919_1875, w_919_1876, w_919_1877, w_919_1878, 
  Loop Gates: I919_1870.port1, I919_1871.port1, I919_1872.port1, I919_1873.port1, I919_1874.port2, I919_1875.port1, I919_1876.port2, I919_1877.port1, 

59)
  Loop Signals: w_209_1547, w_209_1548, w_209_1549, w_209_1550, w_209_1551, w_209_1552, w_209_1553, w_209_1554, w_209_1555, 
  Loop Gates: I209_1546.port2, I209_1547.port2, I209_1548.port2, I209_1549.port2, I209_1550.port2, I209_1551.port1, I209_1552.port1, I209_1553.port1, I209_1554.port1, 

60)
  Loop Signals: w_669_137, w_669_138, w_669_139, w_669_140, w_669_141, w_669_142, w_669_143, w_669_144, w_669_145, 
  Loop Gates: I669_136.port1, I669_137.port1, I669_138.port2, I669_139.port1, I669_140.port2, I669_141.port2, I669_142.port1, I669_143.port1, I669_144.port2, 

61)
  Loop Signals: w_897_1329, w_897_1330, w_897_1331, w_897_1332, w_897_1333, w_897_1334, w_897_1335, w_897_1336, w_897_1337, w_897_1338, 
  Loop Gates: I897_1328.port2, I897_1329.port1, I897_1330.port1, I897_1331.port1, I897_1332.port1, I897_1333.port2, I897_1334.port2, I897_1335.port1, I897_1336.port2, I897_1337.port1, 

62)
  Loop Signals: w_941_1118, w_941_1119, w_941_1120, 
  Loop Gates: I941_1117.port1, I941_1118.port1, I941_1119.port2, 

63)
  Loop Signals: w_116_1549, w_116_1550, w_116_1551, w_116_1552, w_116_1553, w_116_1554, w_116_1555, w_116_1556, w_116_1557, w_116_1558, 
  Loop Gates: I116_1548.port2, I116_1549.port1, I116_1550.port2, I116_1551.port1, I116_1552.port2, I116_1553.port2, I116_1554.port1, I116_1555.port1, I116_1556.port1, I116_1557.port2, 

64)
  Loop Signals: w_116_1550, w_116_1562, w_116_1563, w_116_1564, w_116_1565, w_116_1566, w_116_1567, w_116_1568, w_116_1569, w_116_1570, w_116_1571, w_116_1572, w_116_1574, 
  Loop Gates: I116_1548.port1, I116_1558.port1, I116_1559.port1, I116_1560.port2, I116_1561.port1, I116_1562.port1, I116_1563.port2, I116_1564.port1, I116_1565.port1, I116_1566.port2, I116_1567.port2, I116_1568.port1, I116_1569.port2, 

65)
  Loop Signals: w_1666_1997, w_1666_1998, w_1666_1999, w_1666_2000, w_1666_2001, w_1666_2002, w_1666_2003, w_1666_2004, w_1666_2005, w_1666_2006, w_1666_2007, w_1666_2008, 
  Loop Gates: I1666_1996.port1, I1666_1997.port1, I1666_1998.port1, I1666_1999.port2, I1666_2000.port2, I1666_2001.port1, I1666_2002.port1, I1666_2003.port2, I1666_2004.port2, I1666_2005.port1, I1666_2006.port1, I1666_2007.port1, 

66)
  Loop Signals: w_1666_2002, w_1666_2012, w_1666_2013, w_1666_2014, w_1666_2016, 
  Loop Gates: I1666_2000.port1, I1666_2008.port1, I1666_2009.port2, I1666_2010.port1, I1666_2011.port2, 

67)
  Loop Signals: w_1199_1954, w_1199_1955, w_1199_1956, 
  Loop Gates: I1199_1953.port1, I1199_1954.port1, I1199_1955.port1, 

68)
  Loop Signals: w_1199_1954, w_1199_1960, w_1199_1961, w_1199_1962, w_1199_1963, w_1199_1964, w_1199_1965, w_1199_1966, w_1199_1967, w_1199_1968, w_1199_1969, w_1199_1970, w_1199_1971, w_1199_1973, 
  Loop Gates: I1199_1955.port2, I1199_1956.port1, I1199_1957.port1, I1199_1958.port1, I1199_1959.port2, I1199_1960.port1, I1199_1961.port1, I1199_1962.port1, I1199_1963.port1, I1199_1964.port2, I1199_1965.port1, I1199_1966.port1, I1199_1967.port1, I1199_1968.port2, 

69)
  Loop Signals: w_1598_1875, w_1598_1876, w_1598_1877, w_1598_1878, w_1598_1879, w_1598_1880, w_1598_1881, w_1598_1882, w_1598_1883, w_1598_1884, w_1598_1885, 
  Loop Gates: I1598_1874.port2, I1598_1875.port1, I1598_1876.port2, I1598_1877.port1, I1598_1878.port1, I1598_1879.port2, I1598_1880.port1, I1598_1881.port1, I1598_1882.port2, I1598_1883.port2, I1598_1884.port1, 

70)
  Loop Signals: w_1055_453, w_1055_454, w_1055_455, w_1055_456, w_1055_457, w_1055_458, w_1055_459, w_1055_460, w_1055_461, w_1055_462, w_1055_463, w_1055_464, 
  Loop Gates: I1055_452.port1, I1055_453.port1, I1055_454.port1, I1055_455.port1, I1055_456.port1, I1055_457.port2, I1055_458.port1, I1055_459.port2, I1055_460.port2, I1055_461.port2, I1055_462.port2, I1055_463.port1, 

71)
  Loop Signals: w_110_1611, w_110_1612, w_110_1613, w_110_1614, w_110_1615, w_110_1616, w_110_1617, 
  Loop Gates: I110_1610.port1, I110_1611.port1, I110_1612.port2, I110_1613.port2, I110_1614.port1, I110_1615.port2, I110_1616.port2, 

72)
  Loop Signals: w_110_1612, w_110_1621, w_110_1622, w_110_1623, w_110_1624, w_110_1625, w_110_1626, w_110_1627, w_110_1628, w_110_1629, w_110_1630, w_110_1631, w_110_1633, 
  Loop Gates: I110_1610.port2, I110_1617.port2, I110_1618.port1, I110_1619.port1, I110_1620.port1, I110_1621.port2, I110_1622.port1, I110_1623.port2, I110_1624.port1, I110_1625.port1, I110_1626.port2, I110_1627.port1, I110_1628.port2, 

73)
  Loop Signals: w_1312_969, w_1312_970, w_1312_971, w_1312_972, w_1312_973, w_1312_974, w_1312_975, w_1312_976, w_1312_977, w_1312_978, w_1312_979, w_1312_980, 
  Loop Gates: I1312_968.port1, I1312_969.port1, I1312_970.port1, I1312_971.port1, I1312_972.port2, I1312_973.port1, I1312_974.port1, I1312_975.port1, I1312_976.port2, I1312_977.port1, I1312_978.port2, I1312_979.port2, 

74)
  Loop Signals: w_1312_969, w_1312_984, w_1312_985, w_1312_986, w_1312_988, 
  Loop Gates: I1312_979.port1, I1312_980.port1, I1312_981.port1, I1312_982.port1, I1312_983.port2, 

75)
  Loop Signals: w_1422_540, w_1422_541, w_1422_542, w_1422_543, w_1422_544, 
  Loop Gates: I1422_539.port2, I1422_540.port1, I1422_541.port1, I1422_542.port1, I1422_543.port1, 

76)
  Loop Signals: w_976_287, w_976_288, w_976_289, w_976_290, w_976_291, w_976_292, w_976_293, w_976_294, w_976_295, 
  Loop Gates: I976_286.port1, I976_287.port2, I976_288.port1, I976_289.port2, I976_290.port1, I976_291.port2, I976_292.port2, I976_293.port2, I976_294.port2, 

77)
  Loop Signals: w_976_295, w_976_299, w_976_300, w_976_301, w_976_303, 
  Loop Gates: I976_293.port1, I976_295.port2, I976_296.port1, I976_297.port1, I976_298.port2, 

78)
  Loop Signals: w_1078_081, w_1078_082, w_1078_083, w_1078_084, w_1078_085, w_1078_086, w_1078_087, w_1078_088, w_1078_089, w_1078_090, w_1078_091, w_1078_092, 
  Loop Gates: I1078_080.port1, I1078_081.port2, I1078_082.port2, I1078_083.port1, I1078_084.port1, I1078_085.port1, I1078_086.port1, I1078_087.port1, I1078_088.port1, I1078_089.port1, I1078_090.port1, I1078_091.port1, 

79)
  Loop Signals: w_1118_1455, w_1118_1456, w_1118_1457, w_1118_1458, w_1118_1459, w_1118_1460, w_1118_1461, w_1118_1462, w_1118_1463, w_1118_1464, 
  Loop Gates: I1118_1454.port2, I1118_1455.port1, I1118_1456.port2, I1118_1457.port1, I1118_1458.port1, I1118_1459.port2, I1118_1460.port1, I1118_1461.port1, I1118_1462.port1, I1118_1463.port1, 

80)
  Loop Signals: w_863_389, w_863_390, w_863_391, w_863_392, w_863_393, w_863_394, 
  Loop Gates: I863_388.port2, I863_389.port2, I863_390.port1, I863_391.port2, I863_392.port2, I863_393.port2, 

81)
  Loop Signals: w_863_389, w_863_398, w_863_399, w_863_400, w_863_401, w_863_402, w_863_403, w_863_404, w_863_405, w_863_406, w_863_407, w_863_408, w_863_409, w_863_411, 
  Loop Gates: I863_393.port1, I863_394.port1, I863_395.port1, I863_396.port1, I863_397.port1, I863_398.port1, I863_399.port1, I863_400.port1, I863_401.port1, I863_402.port1, I863_403.port2, I863_404.port1, I863_405.port1, I863_406.port2, 

82)
  Loop Signals: w_996_1460, w_996_1461, w_996_1462, w_996_1463, w_996_1464, w_996_1465, w_996_1466, w_996_1467, 
  Loop Gates: I996_1459.port1, I996_1460.port1, I996_1461.port1, I996_1462.port1, I996_1463.port2, I996_1464.port1, I996_1465.port2, I996_1466.port2, 

83)
  Loop Signals: w_996_1465, w_996_1471, w_996_1472, w_996_1473, w_996_1474, w_996_1475, w_996_1476, w_996_1477, w_996_1478, w_996_1479, w_996_1480, w_996_1482, 
  Loop Gates: I996_1463.port1, I996_1467.port2, I996_1468.port1, I996_1469.port1, I996_1470.port1, I996_1471.port2, I996_1472.port1, I996_1473.port1, I996_1474.port1, I996_1475.port1, I996_1476.port1, I996_1477.port2, 

84)
  Loop Signals: w_399_1788, w_399_1789, w_399_1790, w_399_1791, w_399_1792, w_399_1793, w_399_1794, w_399_1795, w_399_1796, w_399_1797, w_399_1798, 
  Loop Gates: I399_1787.port1, I399_1788.port1, I399_1789.port2, I399_1790.port1, I399_1791.port1, I399_1792.port1, I399_1793.port1, I399_1794.port1, I399_1795.port1, I399_1796.port1, I399_1797.port1, 

85)
  Loop Signals: w_399_1791, w_399_1802, w_399_1803, w_399_1804, w_399_1806, 
  Loop Gates: I399_1789.port1, I399_1798.port1, I399_1799.port1, I399_1800.port1, I399_1801.port2, 

86)
  Loop Signals: w_1112_1748, w_1112_1749, w_1112_1750, w_1112_1751, w_1112_1752, w_1112_1753, w_1112_1754, w_1112_1755, w_1112_1756, 
  Loop Gates: I1112_1747.port2, I1112_1748.port1, I1112_1749.port1, I1112_1750.port2, I1112_1751.port1, I1112_1752.port1, I1112_1753.port2, I1112_1754.port1, I1112_1755.port1, 

87)
  Loop Signals: w_1289_456, w_1289_457, w_1289_458, w_1289_459, w_1289_460, w_1289_461, w_1289_462, w_1289_463, 
  Loop Gates: I1289_456.port1, I1289_457.port1, I1289_458.port1, I1289_459.port1, I1289_460.port1, I1289_461.port2, I1289_462.port1, I1289_463.port2, 

88)
  Loop Signals: w_966_461, w_966_462, w_966_463, w_966_464, w_966_465, w_966_466, 
  Loop Gates: I966_460.port1, I966_461.port2, I966_462.port2, I966_463.port1, I966_464.port1, I966_465.port2, 

89)
  Loop Signals: w_966_462, w_966_470, w_966_471, w_966_472, w_966_473, w_966_474, w_966_475, w_966_476, w_966_477, w_966_478, w_966_480, 
  Loop Gates: I966_460.port2, I966_466.port1, I966_467.port2, I966_468.port1, I966_469.port1, I966_470.port1, I966_471.port1, I966_472.port1, I966_473.port2, I966_474.port1, I966_475.port2, 

90)
  Loop Signals: w_1824_1452, w_1824_1453, w_1824_1454, 
  Loop Gates: I1824_1451.port1, I1824_1452.port1, I1824_1453.port2, 

91)
  Loop Signals: w_148_1915, w_148_1916, w_148_1917, w_148_1918, w_148_1919, w_148_1920, w_148_1921, w_148_1922, w_148_1923, w_148_1924, w_148_1925, 
  Loop Gates: I148_1914.port1, I148_1915.port1, I148_1916.port1, I148_1917.port2, I148_1918.port1, I148_1919.port1, I148_1920.port1, I148_1921.port2, I148_1922.port1, I148_1923.port1, I148_1924.port2, 

92)
  Loop Signals: w_1275_1432, w_1275_1433, w_1275_1434, w_1275_1435, w_1275_1436, w_1275_1437, w_1275_1438, w_1275_1439, w_1275_1440, 
  Loop Gates: I1275_1431.port2, I1275_1432.port1, I1275_1433.port1, I1275_1434.port1, I1275_1435.port1, I1275_1436.port1, I1275_1437.port2, I1275_1438.port1, I1275_1439.port1, 

93)
  Loop Signals: w_1275_1436, w_1275_1444, w_1275_1445, w_1275_1446, w_1275_1447, w_1275_1448, w_1275_1449, w_1275_1450, w_1275_1451, w_1275_1452, w_1275_1453, w_1275_1454, w_1275_1456, 
  Loop Gates: I1275_1434.port2, I1275_1440.port1, I1275_1441.port1, I1275_1442.port2, I1275_1443.port1, I1275_1444.port1, I1275_1445.port1, I1275_1446.port1, I1275_1447.port1, I1275_1448.port2, I1275_1449.port1, I1275_1450.port1, I1275_1451.port2, 

94)
  Loop Signals: w_493_572, w_493_573, w_493_574, w_493_575, w_493_576, w_493_577, w_493_578, 
  Loop Gates: I493_571.port2, I493_572.port1, I493_573.port1, I493_574.port2, I493_575.port1, I493_576.port1, I493_577.port1, 

95)
  Loop Signals: w_493_573, w_493_582, w_493_583, w_493_584, w_493_585, w_493_586, w_493_587, w_493_589, 
  Loop Gates: I493_571.port1, I493_578.port1, I493_579.port1, I493_580.port1, I493_581.port2, I493_582.port1, I493_583.port1, I493_584.port2, 

96)
  Loop Signals: w_1688_1681, w_1688_1682, w_1688_1683, w_1688_1684, w_1688_1685, w_1688_1686, w_1688_1687, w_1688_1688, 
  Loop Gates: I1688_1680.port1, I1688_1681.port1, I1688_1682.port1, I1688_1683.port1, I1688_1684.port1, I1688_1685.port1, I1688_1686.port1, I1688_1687.port2, 

97)
  Loop Signals: w_022_440, w_022_441, w_022_442, w_022_443, w_022_444, w_022_445, w_022_446, w_022_447, 
  Loop Gates: I022_439.port2, I022_440.port1, I022_441.port2, I022_442.port1, I022_443.port1, I022_444.port1, I022_445.port1, I022_446.port1, 

98)
  Loop Signals: w_022_451, w_022_452, w_022_453, w_022_454, w_022_455, w_022_456, w_022_457, w_022_458, w_022_459, 
  Loop Gates: I022_447.port2, I022_448.port2, I022_449.port2, I022_450.port1, I022_451.port1, I022_452.port2, I022_453.port2, I022_454.port2, I022_455.port2, 

99)
  Loop Signals: w_722_1621, w_722_1622, w_722_1623, w_722_1624, w_722_1625, w_722_1626, w_722_1627, w_722_1628, 
  Loop Gates: I722_1620.port2, I722_1621.port2, I722_1622.port2, I722_1623.port1, I722_1624.port2, I722_1625.port1, I722_1626.port1, I722_1627.port2, 

******* result_2.txt *********
1)
  Loop Signals: w_054_628, w_054_629, w_054_630, w_054_631, w_054_632, w_054_633, w_054_634, w_054_635, w_054_636, w_054_637, 
  Loop Gates: I054_627.port2, I054_628.port1, I054_629.port1, I054_630.port2, I054_631.port1, I054_632.port1, I054_633.port1, I054_634.port2, I054_635.port1, I054_636.port2, 

2)
  Loop Signals: w_457_1221, w_457_1222, w_457_1223, w_457_1224, w_457_1225, w_457_1226, 
  Loop Gates: I457_1220.port2, I457_1221.port1, I457_1222.port1, I457_1223.port2, I457_1224.port1, I457_1225.port1, 

3)
  Loop Signals: w_484_492, w_484_493, w_484_494, 
  Loop Gates: I484_491.port1, I484_492.port1, I484_493.port1, 

4)
  Loop Signals: w_484_492, w_484_498, w_484_499, w_484_500, w_484_501, w_484_502, w_484_503, w_484_504, w_484_505, w_484_506, w_484_507, w_484_509, 
  Loop Gates: I484_493.port2, I484_494.port1, I484_495.port1, I484_496.port2, I484_497.port1, I484_498.port1, I484_499.port1, I484_500.port2, I484_501.port1, I484_502.port1, I484_503.port1, I484_504.port2, 

5)
  Loop Signals: w_1818_359, w_1818_360, w_1818_361, w_1818_362, 
  Loop Gates: I1818_358.port1, I1818_359.port2, I1818_360.port1, I1818_361.port1, 

6)
  Loop Signals: w_799_855, w_799_860, w_799_861, w_799_862, w_799_863, w_799_865, 
  Loop Gates: I799_853.port2, I799_856.port1, I799_857.port1, I799_858.port1, I799_859.port1, I799_860.port2, 

7)
  Loop Signals: w_235_1042, w_235_1043, w_235_1044, w_235_1045, w_235_1046, w_235_1047, w_235_1048, 
  Loop Gates: I235_1041.port2, I235_1042.port2, I235_1043.port1, I235_1044.port2, I235_1045.port1, I235_1046.port1, I235_1047.port1, 

8)
  Loop Signals: w_235_1047, w_235_1052, w_235_1053, w_235_1054, w_235_1055, w_235_1056, w_235_1057, w_235_1058, w_235_1059, w_235_1060, w_235_1062, 
  Loop Gates: I235_1045.port2, I235_1048.port2, I235_1049.port2, I235_1050.port1, I235_1051.port1, I235_1052.port2, I235_1053.port2, I235_1054.port1, I235_1055.port1, I235_1056.port1, I235_1057.port2, 

9)
  Loop Signals: w_811_1656, w_811_1657, w_811_1658, 
  Loop Gates: I811_1655.port1, I811_1656.port1, I811_1657.port2, 

10)
  Loop Signals: w_432_726, w_432_727, w_432_728, w_432_729, w_432_730, w_432_731, 
  Loop Gates: I432_725.port1, I432_726.port2, I432_727.port1, I432_728.port1, I432_729.port2, I432_730.port1, 

11)
  Loop Signals: w_769_203, w_769_204, w_769_205, w_769_206, w_769_207, w_769_208, w_769_209, 
  Loop Gates: I769_202.port2, I769_203.port2, I769_204.port1, I769_205.port1, I769_206.port1, I769_207.port2, I769_208.port1, 

12)
  Loop Signals: w_1656_1927, w_1656_1928, w_1656_1929, w_1656_1930, 
  Loop Gates: I1656_1926.port2, I1656_1927.port1, I1656_1928.port1, I1656_1929.port1, 

13)
  Loop Signals: w_1692_766, w_1692_767, w_1692_768, w_1692_769, w_1692_770, 
  Loop Gates: I1692_765.port1, I1692_766.port1, I1692_767.port2, I1692_768.port1, I1692_769.port1, 

14)
  Loop Signals: w_1298_518, w_1298_519, w_1298_520, 
  Loop Gates: I1298_517.port1, I1298_518.port2, I1298_519.port2, 

15)
  Loop Signals: w_494_1931, w_494_1932, w_494_1933, w_494_1934, w_494_1935, w_494_1936, 
  Loop Gates: I494_1930.port1, I494_1931.port2, I494_1932.port2, I494_1933.port2, I494_1934.port2, I494_1935.port1, 

16)
  Loop Signals: w_563_960, w_563_961, w_563_962, w_563_963, 
  Loop Gates: I563_959.port1, I563_960.port1, I563_961.port2, I563_962.port2, 

17)
  Loop Signals: w_342_1768, w_342_1769, w_342_1770, w_342_1771, w_342_1772, w_342_1773, w_342_1774, w_342_1775, w_342_1776, w_342_1777, 
  Loop Gates: I342_1767.port2, I342_1768.port2, I342_1769.port1, I342_1770.port1, I342_1771.port2, I342_1772.port2, I342_1773.port1, I342_1774.port2, I342_1775.port2, I342_1776.port1, 

18)
  Loop Signals: w_342_1775, w_342_1781, w_342_1782, w_342_1783, w_342_1784, w_342_1785, w_342_1786, w_342_1788, 
  Loop Gates: I342_1773.port2, I342_1777.port2, I342_1778.port1, I342_1779.port1, I342_1780.port2, I342_1781.port2, I342_1782.port1, I342_1783.port2, 

19)
  Loop Signals: w_1288_1604, w_1288_1611, w_1288_1612, w_1288_1613, w_1288_1614, w_1288_1615, w_1288_1616, w_1288_1617, w_1288_1618, w_1288_1619, w_1288_1620, w_1288_1622, 
  Loop Gates: I1288_1602.port2, I1288_1607.port2, I1288_1608.port1, I1288_1609.port1, I1288_1610.port1, I1288_1611.port1, I1288_1612.port1, I1288_1613.port1, I1288_1614.port2, I1288_1615.port2, I1288_1616.port1, I1288_1617.port2, 

20)
  Loop Signals: w_009_113, w_009_114, w_009_115, w_009_116, w_009_117, w_009_118, w_009_119, w_009_120, 
  Loop Gates: I009_112.port2, I009_113.port1, I009_114.port1, I009_115.port1, I009_116.port2, I009_117.port2, I009_118.port1, I009_119.port1, 

21)
  Loop Signals: w_009_118, w_009_124, w_009_125, w_009_126, w_009_127, w_009_128, w_009_129, w_009_131, 
  Loop Gates: I009_116.port1, I009_120.port1, I009_121.port1, I009_122.port2, I009_123.port1, I009_124.port1, I009_125.port1, I009_126.port2, 

22)
  Loop Signals: w_1423_462, w_1423_463, w_1423_464, w_1423_465, w_1423_466, w_1423_467, w_1423_468, w_1423_469, w_1423_470, w_1423_471, w_1423_472, 
  Loop Gates: I1423_461.port1, I1423_462.port1, I1423_463.port2, I1423_464.port1, I1423_465.port1, I1423_466.port2, I1423_467.port1, I1423_468.port2, I1423_469.port2, I1423_470.port1, I1423_471.port1, 

23)
  Loop Signals: w_531_1378, w_531_1379, w_531_1380, w_531_1381, w_531_1382, w_531_1383, w_531_1384, w_531_1385, w_531_1386, w_531_1387, w_531_1388, 
  Loop Gates: I531_1377.port1, I531_1378.port1, I531_1379.port1, I531_1380.port1, I531_1381.port1, I531_1382.port1, I531_1383.port1, I531_1384.port1, I531_1385.port1, I531_1386.port2, I531_1387.port1, 

24)
  Loop Signals: w_1601_113, w_1601_114, w_1601_115, 
  Loop Gates: I1601_112.port1, I1601_113.port2, I1601_114.port1, 

25)
  Loop Signals: w_1848_117, w_1848_118, w_1848_119, w_1848_120, 
  Loop Gates: I1848_116.port1, I1848_117.port1, I1848_118.port1, I1848_119.port1, 

26)
  Loop Signals: w_1836_1757, w_1836_1758, w_1836_1759, w_1836_1760, w_1836_1761, w_1836_1762, w_1836_1763, w_1836_1764, w_1836_1765, w_1836_1766, w_1836_1767, w_1836_1768, 
  Loop Gates: I1836_1756.port1, I1836_1757.port2, I1836_1758.port1, I1836_1759.port2, I1836_1760.port1, I1836_1761.port1, I1836_1762.port1, I1836_1763.port1, I1836_1764.port2, I1836_1765.port1, I1836_1766.port2, I1836_1767.port1, 

27)
  Loop Signals: w_1836_1768, w_1836_1772, w_1836_1773, w_1836_1774, w_1836_1775, w_1836_1776, w_1836_1778, 
  Loop Gates: I1836_1766.port1, I1836_1768.port1, I1836_1769.port2, I1836_1770.port1, I1836_1771.port2, I1836_1772.port1, I1836_1773.port2, 

28)
  Loop Signals: w_1579_1708, w_1579_1709, w_1579_1710, w_1579_1711, w_1579_1712, w_1579_1713, w_1579_1714, w_1579_1715, 
  Loop Gates: I1579_1707.port1, I1579_1708.port1, I1579_1709.port1, I1579_1710.port1, I1579_1711.port1, I1579_1712.port2, I1579_1713.port1, I1579_1714.port1, 

29)
  Loop Signals: w_851_1288, w_851_1289, w_851_1290, w_851_1291, w_851_1292, w_851_1293, w_851_1294, w_851_1295, w_851_1296, w_851_1297, 
  Loop Gates: I851_1287.port1, I851_1288.port1, I851_1289.port2, I851_1290.port1, I851_1291.port1, I851_1292.port1, I851_1293.port1, I851_1294.port1, I851_1295.port1, I851_1296.port1, 

30)
  Loop Signals: w_1176_1251, w_1176_1252, w_1176_1253, w_1176_1254, w_1176_1255, w_1176_1256, w_1176_1257, w_1176_1258, w_1176_1259, w_1176_1260, w_1176_1261, w_1176_1262, 
  Loop Gates: I1176_1250.port2, I1176_1251.port1, I1176_1252.port1, I1176_1253.port2, I1176_1254.port2, I1176_1255.port1, I1176_1256.port1, I1176_1257.port2, I1176_1258.port1, I1176_1259.port2, I1176_1260.port2, I1176_1261.port1, 

31)
  Loop Signals: w_919_1871, w_919_1872, w_919_1873, w_919_1874, w_919_1875, w_919_1876, w_919_1877, w_919_1878, 
  Loop Gates: I919_1870.port1, I919_1871.port1, I919_1872.port1, I919_1873.port1, I919_1874.port2, I919_1875.port1, I919_1876.port2, I919_1877.port1, 

32)
  Loop Signals: w_209_1547, w_209_1548, w_209_1549, w_209_1550, w_209_1551, w_209_1552, w_209_1553, w_209_1554, w_209_1555, 
  Loop Gates: I209_1546.port2, I209_1547.port2, I209_1548.port2, I209_1549.port2, I209_1550.port2, I209_1551.port1, I209_1552.port1, I209_1553.port1, I209_1554.port1, 

33)
  Loop Signals: w_669_137, w_669_138, w_669_139, w_669_140, w_669_141, w_669_142, w_669_143, w_669_144, w_669_145, 
  Loop Gates: I669_136.port1, I669_137.port1, I669_138.port2, I669_139.port1, I669_140.port2, I669_141.port2, I669_142.port1, I669_143.port1, I669_144.port2, 

34)
  Loop Signals: w_941_1118, w_941_1119, w_941_1120, 
  Loop Gates: I941_1117.port1, I941_1118.port1, I941_1119.port2, 

35)
  Loop Signals: w_1666_1997, w_1666_1998, w_1666_1999, w_1666_2000, w_1666_2001, w_1666_2002, w_1666_2003, w_1666_2004, w_1666_2005, w_1666_2006, w_1666_2007, w_1666_2008, 
  Loop Gates: I1666_1996.port1, I1666_1997.port1, I1666_1998.port1, I1666_1999.port2, I1666_2000.port2, I1666_2001.port1, I1666_2002.port1, I1666_2003.port2, I1666_2004.port2, I1666_2005.port1, I1666_2006.port1, I1666_2007.port1, 

36)
  Loop Signals: w_1666_2002, w_1666_2012, w_1666_2013, w_1666_2014, w_1666_2016, 
  Loop Gates: I1666_2000.port1, I1666_2008.port1, I1666_2009.port2, I1666_2010.port1, I1666_2011.port2, 

37)
  Loop Signals: w_1199_1954, w_1199_1955, w_1199_1956, 
  Loop Gates: I1199_1953.port1, I1199_1954.port1, I1199_1955.port1, 

38)
  Loop Signals: w_1199_1954, w_1199_1960, w_1199_1961, w_1199_1962, w_1199_1963, w_1199_1964, w_1199_1965, w_1199_1966, w_1199_1967, w_1199_1968, w_1199_1969, w_1199_1970, w_1199_1971, w_1199_1973, 
  Loop Gates: I1199_1955.port2, I1199_1956.port1, I1199_1957.port1, I1199_1958.port1, I1199_1959.port2, I1199_1960.port1, I1199_1961.port1, I1199_1962.port1, I1199_1963.port1, I1199_1964.port2, I1199_1965.port1, I1199_1966.port1, I1199_1967.port1, I1199_1968.port2, 

39)
  Loop Signals: w_1598_1875, w_1598_1876, w_1598_1877, w_1598_1878, w_1598_1879, w_1598_1880, w_1598_1881, w_1598_1882, w_1598_1883, w_1598_1884, w_1598_1885, 
  Loop Gates: I1598_1874.port2, I1598_1875.port1, I1598_1876.port2, I1598_1877.port1, I1598_1878.port1, I1598_1879.port2, I1598_1880.port1, I1598_1881.port1, I1598_1882.port2, I1598_1883.port2, I1598_1884.port1, 

40)
  Loop Signals: w_1055_453, w_1055_454, w_1055_455, w_1055_456, w_1055_457, w_1055_458, w_1055_459, w_1055_460, w_1055_461, w_1055_462, w_1055_463, w_1055_464, 
  Loop Gates: I1055_452.port1, I1055_453.port1, I1055_454.port1, I1055_455.port1, I1055_456.port1, I1055_457.port2, I1055_458.port1, I1055_459.port2, I1055_460.port2, I1055_461.port2, I1055_462.port2, I1055_463.port1, 

41)
  Loop Signals: w_110_1612, w_110_1621, w_110_1622, w_110_1623, w_110_1624, w_110_1625, w_110_1626, w_110_1627, w_110_1628, w_110_1629, w_110_1630, w_110_1631, w_110_1633, 
  Loop Gates: I110_1610.port2, I110_1617.port2, I110_1618.port1, I110_1619.port1, I110_1620.port1, I110_1621.port2, I110_1622.port1, I110_1623.port2, I110_1624.port1, I110_1625.port1, I110_1626.port2, I110_1627.port1, I110_1628.port2, 

42)
  Loop Signals: w_1312_969, w_1312_970, w_1312_971, w_1312_972, w_1312_973, w_1312_974, w_1312_975, w_1312_976, w_1312_977, w_1312_978, w_1312_979, w_1312_980, 
  Loop Gates: I1312_968.port1, I1312_969.port1, I1312_970.port1, I1312_971.port1, I1312_972.port2, I1312_973.port1, I1312_974.port1, I1312_975.port1, I1312_976.port2, I1312_977.port1, I1312_978.port2, I1312_979.port2, 

43)
  Loop Signals: w_1422_540, w_1422_541, w_1422_542, w_1422_543, w_1422_544, 
  Loop Gates: I1422_539.port2, I1422_540.port1, I1422_541.port1, I1422_542.port1, I1422_543.port1, 

44)
  Loop Signals: w_863_389, w_863_390, w_863_391, w_863_392, w_863_393, w_863_394, 
  Loop Gates: I863_388.port2, I863_389.port2, I863_390.port1, I863_391.port2, I863_392.port2, I863_393.port2, 

45)
  Loop Signals: w_863_389, w_863_398, w_863_399, w_863_400, w_863_401, w_863_402, w_863_403, w_863_404, w_863_405, w_863_406, w_863_407, w_863_408, w_863_409, w_863_411, 
  Loop Gates: I863_393.port1, I863_394.port1, I863_395.port1, I863_396.port1, I863_397.port1, I863_398.port1, I863_399.port1, I863_400.port1, I863_401.port1, I863_402.port1, I863_403.port2, I863_404.port1, I863_405.port1, I863_406.port2, 

46)
  Loop Signals: w_1824_1452, w_1824_1453, w_1824_1454, 
  Loop Gates: I1824_1451.port1, I1824_1452.port1, I1824_1453.port2, 

47)
  Loop Signals: w_1275_1432, w_1275_1433, w_1275_1434, w_1275_1435, w_1275_1436, w_1275_1437, w_1275_1438, w_1275_1439, w_1275_1440, 
  Loop Gates: I1275_1431.port2, I1275_1432.port1, I1275_1433.port1, I1275_1434.port1, I1275_1435.port1, I1275_1436.port1, I1275_1437.port2, I1275_1438.port1, I1275_1439.port1, 

48)
  Loop Signals: w_493_573, w_493_582, w_493_583, w_493_584, w_493_585, w_493_586, w_493_587, w_493_589, 
  Loop Gates: I493_571.port1, I493_578.port1, I493_579.port1, I493_580.port1, I493_581.port2, I493_582.port1, I493_583.port1, I493_584.port2, 

49)
  Loop Signals: w_1688_1681, w_1688_1682, w_1688_1683, w_1688_1684, w_1688_1685, w_1688_1686, w_1688_1687, w_1688_1688, 
  Loop Gates: I1688_1680.port1, I1688_1681.port1, I1688_1682.port1, I1688_1683.port1, I1688_1684.port1, I1688_1685.port1, I1688_1686.port1, I1688_1687.port2, 

******* result_3.txt *********
1)
  Loop Signals: w_894_586, w_894_587, w_894_588, w_894_589, w_894_590, w_894_591, 
  Loop Gates: I894_585.port1, I894_586.port2, I894_587.port2, I894_588.port2, I894_589.port1, I894_590.port1, 
  Loop Conditions: I894_585.port2=1, I894_586.port1=1, I894_587.port1=1, I894_588.port1=0, I894_589.port2=1, I894_590.port2=1, 
  (Signal Values: w_083_015=1, w_116_454=1, w_164_146=0, w_489_1324=1, w_570_1461=1, w_894_607=1, )

2)
  Loop Signals: w_894_586, w_894_595, w_894_596, w_894_597, w_894_598, w_894_599, w_894_600, w_894_601, w_894_602, w_894_603, w_894_604, w_894_605, w_894_607, 
  Loop Gates: I894_590.port2, I894_591.port1, I894_592.port1, I894_593.port1, I894_594.port1, I894_595.port2, I894_596.port1, I894_597.port1, I894_598.port2, I894_599.port2, I894_600.port1, I894_601.port1, I894_602.port2, 
  Loop Conditions: I894_590.port2=1, I894_593.port2=1, I894_594.port2=1, I894_595.port1=1, I894_597.port2=0, I894_598.port1=1, I894_599.port1=1, I894_600.port2=0, I894_602.port2=1, 
  (Signal Values: w_144_763=1, w_178_586=1, w_252_382=1, w_451_632=0, w_525_366=1, w_762_973=1, w_789_059=0, w_894_605=1, w_894_607=1, )

3)
  Loop Signals: w_102_1259, w_102_1260, w_102_1261, w_102_1262, w_102_1263, w_102_1264, 
  Loop Gates: I102_1258.port1, I102_1259.port2, I102_1260.port2, I102_1261.port2, I102_1262.port1, I102_1263.port1, 
  Loop Conditions: I102_1258.port2=1, I102_1259.port1=1, I102_1260.port1=1, I102_1261.port1=0, I102_1262.port2=1, I102_1263.port2=1, 
  (Signal Values: w_018_055=1, w_026_1029=0, w_026_838=1, w_040_724=1, w_058_054=1, w_102_1278=1, )

4)
  Loop Signals: w_102_1259, w_102_1268, w_102_1269, w_102_1270, w_102_1271, w_102_1272, w_102_1273, w_102_1274, w_102_1275, w_102_1276, w_102_1278, 
  Loop Gates: I102_1263.port2, I102_1264.port1, I102_1265.port1, I102_1266.port2, I102_1267.port2, I102_1268.port2, I102_1269.port1, I102_1270.port2, I102_1271.port1, I102_1272.port1, I102_1273.port2, 
  Loop Conditions: I102_1263.port2=1, I102_1264.port2=1, I102_1265.port2=1, I102_1266.port1=0, I102_1267.port1=1, I102_1268.port1=1, I102_1269.port2=1, I102_1270.port1=1, I102_1273.port2=1, 
  (Signal Values: w_003_114=1, w_007_874=0, w_045_405=1, w_046_119=1, w_073_073=1, w_076_138=1, w_086_1093=1, w_102_1276=1, w_102_1278=1, )

5)
  Loop Signals: w_799_848, w_799_849, w_799_850, w_799_851, w_799_852, w_799_853, w_799_854, w_799_855, w_799_856, 
  Loop Gates: I799_847.port1, I799_848.port2, I799_849.port2, I799_850.port1, I799_851.port1, I799_852.port1, I799_853.port1, I799_854.port1, I799_855.port2, 
  Loop Conditions: I799_847.port2=0, I799_848.port1=0, I799_849.port1=0, I799_850.port2=1, I799_852.port2=1, I799_853.port2=1, I799_855.port1=1, 
  (Signal Values: w_024_882=1, w_271_175=1, w_496_495=0, w_651_012=1, w_674_050=0, w_773_158=0, w_799_865=1, )

6)
  Loop Signals: w_811_1656, w_811_1662, w_811_1663, w_811_1664, w_811_1665, w_811_1666, w_811_1667, w_811_1668, w_811_1670, 
  Loop Gates: I811_1657.port1, I811_1658.port1, I811_1659.port1, I811_1660.port1, I811_1661.port2, I811_1662.port1, I811_1663.port1, I811_1664.port1, I811_1665.port2, 
  Loop Conditions: I811_1657.port2=1, I811_1659.port2=1, I811_1661.port1=0, I811_1665.port2=1, 
  (Signal Values: w_232_480=0, w_674_041=1, w_811_1658=1, w_811_1668=1, )

7)
  Loop Signals: w_432_726, w_432_735, w_432_736, w_432_737, w_432_738, w_432_739, w_432_741, 
  Loop Gates: I432_730.port2, I432_731.port2, I432_732.port2, I432_733.port2, I432_734.port1, I432_735.port1, I432_736.port2, 
  Loop Conditions: I432_730.port2=1, I432_731.port1=0, I432_732.port1=1, I432_733.port1=1, I432_736.port2=1, 
  (Signal Values: w_059_353=0, w_068_126=1, w_144_1040=1, w_432_739=1, w_432_741=1, )

8)
  Loop Signals: w_1692_769, w_1692_774, w_1692_775, w_1692_776, w_1692_777, w_1692_778, w_1692_779, w_1692_780, w_1692_782, 
  Loop Gates: I1692_767.port1, I1692_770.port1, I1692_771.port2, I1692_772.port1, I1692_773.port2, I1692_774.port1, I1692_775.port1, I1692_776.port1, I1692_777.port2, 
  Loop Conditions: I1692_767.port2=0, I1692_770.port2=0, I1692_771.port1=0, I1692_773.port1=1, I1692_774.port2=1, I1692_777.port2=1, 
  (Signal Values: w_186_165=1, w_336_1630=1, w_1239_502=0, w_1629_026=0, w_1692_768=0, w_1692_780=1, )

9)
  Loop Signals: w_1298_518, w_1298_524, w_1298_525, w_1298_526, w_1298_527, w_1298_529, 
  Loop Gates: I1298_519.port1, I1298_520.port1, I1298_521.port2, I1298_522.port1, I1298_523.port1, I1298_524.port2, 
  Loop Conditions: I1298_519.port2=1, I1298_520.port2=1, I1298_521.port1=1, I1298_522.port2=0, I1298_524.port2=1, 
  (Signal Values: w_310_019=1, w_855_946=0, w_978_267=1, w_1298_520=1, w_1298_527=1, )

10)
  Loop Signals: w_610_889, w_610_890, w_610_891, w_610_892, w_610_893, w_610_894, w_610_895, w_610_896, w_610_897, w_610_898, w_610_899, 
  Loop Gates: I610_888.port1, I610_889.port1, I610_890.port1, I610_891.port1, I610_892.port1, I610_893.port1, I610_894.port2, I610_895.port1, I610_896.port1, I610_897.port2, I610_898.port1, 
  Loop Conditions: I610_892.port2=1, I610_894.port1=1, I610_896.port2=1, I610_897.port1=0, I610_898.port2=1, 
  (Signal Values: w_041_158=1, w_089_1226=1, w_160_041=1, w_396_560=0, w_463_172=1, )

11)
  Loop Signals: w_1230_965, w_1230_966, w_1230_967, w_1230_968, w_1230_969, w_1230_970, 
  Loop Gates: I1230_964.port2, I1230_965.port1, I1230_966.port1, I1230_967.port1, I1230_968.port2, I1230_969.port1, 
  Loop Conditions: I1230_964.port1=1, I1230_965.port2=0, I1230_966.port2=1, I1230_968.port1=1, I1230_969.port2=1, 
  (Signal Values: w_010_376=1, w_066_007=1, w_563_905=0, w_585_360=1, w_1227_414=1, )

12)
  Loop Signals: w_1288_1602, w_1288_1603, w_1288_1604, w_1288_1605, w_1288_1606, w_1288_1607, 
  Loop Gates: I1288_1601.port1, I1288_1602.port1, I1288_1603.port2, I1288_1604.port1, I1288_1605.port1, I1288_1606.port1, 
  Loop Conditions: I1288_1601.port2=1, I1288_1602.port2=1, I1288_1603.port1=1, 
  (Signal Values: w_576_511=1, w_1033_020=1, w_1288_1622=1, )

13)
  Loop Signals: w_826_437, w_826_438, w_826_439, w_826_440, 
  Loop Gates: I826_436.port1, I826_437.port1, I826_438.port1, I826_439.port1, 
  Loop Conditions: I826_436.port2=0, I826_437.port2=0, I826_438.port2=1, I826_439.port2=1, 
  (Signal Values: w_105_1459=0, w_161_455=0, w_796_506=1, w_826_452=1, )

14)
  Loop Signals: w_826_440, w_826_444, w_826_445, w_826_446, w_826_447, w_826_448, w_826_449, w_826_450, w_826_452, 
  Loop Gates: I826_438.port2, I826_440.port1, I826_441.port1, I826_442.port2, I826_443.port1, I826_444.port1, I826_445.port1, I826_446.port1, I826_447.port2, 
  Loop Conditions: I826_438.port2=1, I826_440.port2=1, I826_441.port2=0, I826_442.port1=1, I826_443.port2=1, I826_444.port2=1, I826_445.port2=1, I826_447.port2=1, 
  (Signal Values: w_016_013=0, w_059_023=1, w_181_1114=1, w_277_292=1, w_501_352=1, w_807_337=1, w_826_450=1, w_826_452=1, )

15)
  Loop Signals: w_1132_1117, w_1132_1118, w_1132_1119, w_1132_1120, w_1132_1121, w_1132_1122, w_1132_1123, 
  Loop Gates: I1132_1116.port1, I1132_1117.port1, I1132_1118.port1, I1132_1119.port2, I1132_1120.port1, I1132_1121.port2, I1132_1122.port2, 
  Loop Conditions: I1132_1116.port2=1, I1132_1118.port2=1, I1132_1119.port1=0, I1132_1121.port1=1, I1132_1122.port1=1, 
  (Signal Values: w_259_272=1, w_287_271=1, w_416_364=1, w_745_034=1, w_796_1386=0, )

16)
  Loop Signals: w_1449_506, w_1449_507, w_1449_508, w_1449_509, 
  Loop Gates: I1449_505.port2, I1449_506.port2, I1449_507.port2, I1449_508.port1, 
  Loop Conditions: I1449_505.port1=0, I1449_506.port1=0, I1449_507.port1=1, I1449_508.port2=0, 
  (Signal Values: w_105_1248=1, w_555_1335=0, w_832_266=0, w_1165_045=0, )

17)
  Loop Signals: w_1308_361, w_1308_362, w_1308_363, w_1308_364, w_1308_365, w_1308_366, w_1308_367, w_1308_368, w_1308_369, w_1308_370, w_1308_371, w_1308_372, 
  Loop Gates: I1308_360.port1, I1308_361.port1, I1308_362.port1, I1308_363.port1, I1308_364.port1, I1308_365.port1, I1308_366.port1, I1308_367.port1, I1308_368.port1, I1308_369.port1, I1308_370.port1, I1308_371.port1, 
  Loop Conditions: I1308_360.port2=0, I1308_363.port2=1, I1308_365.port2=1, I1308_367.port2=1, I1308_368.port2=1, I1308_370.port2=0, 
  (Signal Values: w_204_1002=0, w_332_063=1, w_877_632=1, w_1117_515=1, w_1212_003=1, w_1308_384=0, )

18)
  Loop Signals: w_1308_362, w_1308_376, w_1308_377, w_1308_378, w_1308_379, w_1308_380, w_1308_381, w_1308_382, w_1308_384, 
  Loop Gates: I1308_360.port2, I1308_372.port1, I1308_373.port1, I1308_374.port2, I1308_375.port1, I1308_376.port1, I1308_377.port2, I1308_378.port1, I1308_379.port2, 
  Loop Conditions: I1308_360.port2=0, I1308_372.port2=0, I1308_374.port1=1, I1308_375.port2=1, I1308_377.port1=1, I1308_379.port2=1, 
  (Signal Values: w_107_888=0, w_326_1155=1, w_633_068=1, w_1203_345=1, w_1308_382=1, w_1308_384=0, )

19)
  Loop Signals: w_531_1388, w_531_1392, w_531_1393, w_531_1394, w_531_1395, w_531_1397, 
  Loop Gates: I531_1386.port1, I531_1388.port1, I531_1389.port2, I531_1390.port1, I531_1391.port1, I531_1392.port2, 
  Loop Conditions: I531_1386.port2=1, I531_1389.port1=1, I531_1392.port2=1, 
  (Signal Values: w_386_011=1, w_531_1387=1, w_531_1395=1, )

20)
  Loop Signals: w_1821_248, w_1821_249, w_1821_250, w_1821_251, w_1821_252, w_1821_253, 
  Loop Gates: I1821_247.port2, I1821_248.port2, I1821_249.port1, I1821_250.port1, I1821_251.port2, I1821_252.port1, 
  Loop Conditions: I1821_247.port1=1, I1821_248.port1=1, I1821_249.port2=1, I1821_250.port2=0, I1821_251.port1=1, I1821_252.port2=1, 
  (Signal Values: w_054_544=0, w_514_955=1, w_819_190=1, w_820_664=1, w_1252_023=1, w_1821_268=1, )

21)
  Loop Signals: w_1821_251, w_1821_257, w_1821_258, w_1821_259, w_1821_260, w_1821_261, w_1821_262, w_1821_263, w_1821_264, w_1821_265, w_1821_266, w_1821_268, 
  Loop Gates: I1821_249.port2, I1821_253.port1, I1821_254.port1, I1821_255.port2, I1821_256.port2, I1821_257.port1, I1821_258.port1, I1821_259.port1, I1821_260.port2, I1821_261.port1, I1821_262.port1, I1821_263.port2, 
  Loop Conditions: I1821_249.port2=1, I1821_253.port2=0, I1821_255.port1=1, I1821_256.port1=1, I1821_260.port1=1, I1821_261.port2=1, I1821_263.port2=1, 
  (Signal Values: w_310_477=1, w_352_672=0, w_731_059=1, w_1199_581=1, w_1463_482=1, w_1821_266=1, w_1821_268=1, )

22)
  Loop Signals: w_1601_115, w_1601_119, w_1601_120, w_1601_121, w_1601_122, w_1601_123, w_1601_124, w_1601_125, w_1601_127, 
  Loop Gates: I1601_113.port1, I1601_115.port1, I1601_116.port1, I1601_117.port1, I1601_118.port1, I1601_119.port1, I1601_120.port1, I1601_121.port1, I1601_122.port2, 
  Loop Conditions: I1601_113.port2=0, I1601_115.port2=1, I1601_116.port2=0, I1601_117.port2=1, I1601_118.port2=0, I1601_119.port2=1, I1601_120.port2=1, I1601_122.port2=1, 
  (Signal Values: w_466_103=1, w_901_607=1, w_975_669=0, w_1259_894=1, w_1468_475=1, w_1534_349=0, w_1601_114=0, w_1601_125=1, )

23)
  Loop Signals: w_305_018, w_305_019, w_305_020, w_305_021, w_305_022, w_305_023, w_305_024, 
  Loop Gates: I305_017.port2, I305_018.port1, I305_019.port2, I305_020.port1, I305_021.port1, I305_022.port2, I305_023.port2, 
  Loop Conditions: I305_017.port1=0, I305_019.port1=0, I305_022.port1=0, I305_023.port1=1, 
  (Signal Values: w_003_006=0, w_071_312=0, w_185_1853=1, w_209_638=0, )

24)
  Loop Signals: w_1911_1096, w_1911_1097, w_1911_1098, w_1911_1099, w_1911_1100, w_1911_1101, w_1911_1102, w_1911_1103, w_1911_1104, w_1911_1105, w_1911_1106, w_1911_1107, 
  Loop Gates: I1911_1095.port1, I1911_1096.port1, I1911_1097.port2, I1911_1098.port2, I1911_1099.port1, I1911_1100.port1, I1911_1101.port1, I1911_1102.port1, I1911_1103.port2, I1911_1104.port2, I1911_1105.port1, I1911_1106.port2, 
  Loop Conditions: I1911_1097.port1=1, I1911_1098.port1=1, I1911_1099.port2=1, I1911_1100.port2=1, I1911_1101.port2=0, I1911_1103.port1=0, I1911_1104.port1=1, I1911_1106.port1=0, 
  (Signal Values: w_051_992=0, w_510_177=0, w_798_611=1, w_810_657=1, w_1503_257=1, w_1687_828=1, w_1787_1409=0, w_1801_026=1, )

25)
  Loop Signals: w_299_1759, w_299_1760, w_299_1761, 
  Loop Gates: I299_1758.port1, I299_1759.port2, I299_1760.port1, 
  Loop Conditions: I299_1759.port1=1, 
  (Signal Values: w_235_733=1, )

26)
  Loop Signals: w_1075_1904, w_1075_1905, w_1075_1906, w_1075_1907, w_1075_1908, w_1075_1909, w_1075_1910, w_1075_1911, 
  Loop Gates: I1075_1903.port1, I1075_1904.port1, I1075_1905.port2, I1075_1906.port2, I1075_1907.port1, I1075_1908.port2, I1075_1909.port1, I1075_1910.port1, 
  Loop Conditions: I1075_1905.port1=1, I1075_1906.port1=1, I1075_1907.port2=1, I1075_1908.port2=1, I1075_1910.port2=1, 
  (Signal Values: w_087_1603=1, w_357_083=1, w_697_644=1, w_781_1927=1, w_1075_1909=1, )

27)
  Loop Signals: w_1075_1910, w_1075_1915, w_1075_1916, w_1075_1917, w_1075_1918, w_1075_1919, w_1075_1920, w_1075_1921, w_1075_1922, w_1075_1924, 
  Loop Gates: I1075_1908.port1, I1075_1911.port2, I1075_1912.port1, I1075_1913.port2, I1075_1914.port2, I1075_1915.port1, I1075_1916.port1, I1075_1917.port2, I1075_1918.port1, I1075_1919.port2, 
  Loop Conditions: I1075_1908.port2=1, I1075_1911.port1=1, I1075_1912.port2=1, I1075_1913.port1=1, I1075_1914.port1=0, I1075_1915.port2=1, I1075_1917.port1=1, I1075_1919.port2=1, 
  (Signal Values: w_570_560=1, w_671_330=0, w_809_1170=1, w_827_820=1, w_925_563=1, w_1041_374=1, w_1075_1909=1, w_1075_1922=1, )

28)
  Loop Signals: w_897_1329, w_897_1330, w_897_1331, w_897_1332, w_897_1333, w_897_1334, w_897_1335, w_897_1336, w_897_1337, w_897_1338, 
  Loop Gates: I897_1328.port2, I897_1329.port1, I897_1330.port1, I897_1331.port1, I897_1332.port1, I897_1333.port2, I897_1334.port2, I897_1335.port1, I897_1336.port2, I897_1337.port1, 
  Loop Conditions: I897_1328.port1=1, I897_1329.port2=1, I897_1330.port2=0, I897_1332.port2=1, I897_1333.port1=1, I897_1334.port1=1, I897_1335.port2=1, I897_1336.port1=0, I897_1337.port2=1, 
  (Signal Values: w_087_1494=1, w_093_070=1, w_163_147=1, w_184_002=1, w_211_212=1, w_214_230=1, w_249_423=0, w_354_1250=0, w_650_173=1, )

29)
  Loop Signals: w_116_1549, w_116_1550, w_116_1551, w_116_1552, w_116_1553, w_116_1554, w_116_1555, w_116_1556, w_116_1557, w_116_1558, 
  Loop Gates: I116_1548.port2, I116_1549.port1, I116_1550.port2, I116_1551.port1, I116_1552.port2, I116_1553.port2, I116_1554.port1, I116_1555.port1, I116_1556.port1, I116_1557.port2, 
  Loop Conditions: I116_1548.port2=0, I116_1549.port2=0, I116_1550.port1=1, I116_1551.port2=1, I116_1552.port1=0, I116_1553.port1=1, I116_1554.port2=0, I116_1555.port2=1, I116_1556.port2=1, I116_1557.port1=1, 
  (Signal Values: w_001_1454=0, w_009_036=1, w_022_056=1, w_027_348=1, w_043_059=1, w_059_272=1, w_060_013=0, w_073_101=0, w_077_170=1, w_116_1549=0, )

30)
  Loop Signals: w_116_1550, w_116_1562, w_116_1563, w_116_1564, w_116_1565, w_116_1566, w_116_1567, w_116_1568, w_116_1569, w_116_1570, w_116_1571, w_116_1572, w_116_1574, 
  Loop Gates: I116_1548.port1, I116_1558.port1, I116_1559.port1, I116_1560.port2, I116_1561.port1, I116_1562.port1, I116_1563.port2, I116_1564.port1, I116_1565.port1, I116_1566.port2, I116_1567.port2, I116_1568.port1, I116_1569.port2, 
  Loop Conditions: I116_1548.port2=0, I116_1558.port2=0, I116_1560.port1=1, I116_1562.port2=1, I116_1563.port1=1, I116_1565.port2=1, I116_1566.port1=1, I116_1567.port1=1, I116_1569.port2=1, 
  (Signal Values: w_029_547=1, w_039_1509=1, w_063_590=1, w_071_531=0, w_092_767=1, w_095_279=1, w_115_559=1, w_116_1549=0, w_116_1572=1, )

31)
  Loop Signals: w_110_1611, w_110_1612, w_110_1613, w_110_1614, w_110_1615, w_110_1616, w_110_1617, 
  Loop Gates: I110_1610.port1, I110_1611.port1, I110_1612.port2, I110_1613.port2, I110_1614.port1, I110_1615.port2, I110_1616.port2, 
  Loop Conditions: I110_1610.port2=1, I110_1611.port2=1, I110_1612.port1=1, I110_1613.port1=0, I110_1615.port1=0, I110_1616.port1=1, 
  (Signal Values: w_004_1051=0, w_006_208=1, w_054_073=0, w_072_010=1, w_095_845=1, w_110_1633=1, )

32)
  Loop Signals: w_1312_969, w_1312_984, w_1312_985, w_1312_986, w_1312_988, 
  Loop Gates: I1312_979.port1, I1312_980.port1, I1312_981.port1, I1312_982.port1, I1312_983.port2, 
  Loop Conditions: I1312_979.port2=0, I1312_980.port2=1, I1312_981.port2=0, I1312_983.port2=1, 
  (Signal Values: w_530_1605=1, w_614_388=0, w_1312_980=0, w_1312_986=1, )

33)
  Loop Signals: w_976_287, w_976_288, w_976_289, w_976_290, w_976_291, w_976_292, w_976_293, w_976_294, w_976_295, 
  Loop Gates: I976_286.port1, I976_287.port2, I976_288.port1, I976_289.port2, I976_290.port1, I976_291.port2, I976_292.port2, I976_293.port2, I976_294.port2, 
  Loop Conditions: I976_287.port1=1, I976_288.port2=0, I976_289.port1=1, I976_290.port2=1, I976_291.port1=0, I976_292.port1=0, I976_293.port2=1, I976_294.port1=1, 
  (Signal Values: w_137_112=1, w_164_498=0, w_299_113=0, w_341_249=1, w_427_055=1, w_599_010=0, w_834_1377=1, w_976_294=1, )

34)
  Loop Signals: w_976_295, w_976_299, w_976_300, w_976_301, w_976_303, 
  Loop Gates: I976_293.port1, I976_295.port2, I976_296.port1, I976_297.port1, I976_298.port2, 
  Loop Conditions: I976_293.port2=1, I976_295.port1=0, I976_296.port2=1, I976_298.port2=1, 
  (Signal Values: w_271_056=0, w_660_223=1, w_976_294=1, w_976_301=1, )

35)
  Loop Signals: w_1078_081, w_1078_082, w_1078_083, w_1078_084, w_1078_085, w_1078_086, w_1078_087, w_1078_088, w_1078_089, w_1078_090, w_1078_091, w_1078_092, 
  Loop Gates: I1078_080.port1, I1078_081.port2, I1078_082.port2, I1078_083.port1, I1078_084.port1, I1078_085.port1, I1078_086.port1, I1078_087.port1, I1078_088.port1, I1078_089.port1, I1078_090.port1, I1078_091.port1, 
  Loop Conditions: I1078_080.port2=1, I1078_081.port1=0, I1078_082.port1=1, I1078_085.port2=0, I1078_087.port2=0, I1078_088.port2=0, I1078_089.port2=1, I1078_090.port2=1, 
  (Signal Values: w_026_1287=0, w_498_636=1, w_549_164=1, w_638_1113=0, w_845_041=1, w_1017_151=1, w_1018_190=0, w_1069_579=0, )

36)
  Loop Signals: w_1118_1455, w_1118_1456, w_1118_1457, w_1118_1458, w_1118_1459, w_1118_1460, w_1118_1461, w_1118_1462, w_1118_1463, w_1118_1464, 
  Loop Gates: I1118_1454.port2, I1118_1455.port1, I1118_1456.port2, I1118_1457.port1, I1118_1458.port1, I1118_1459.port2, I1118_1460.port1, I1118_1461.port1, I1118_1462.port1, I1118_1463.port1, 
  Loop Conditions: I1118_1454.port1=0, I1118_1455.port2=0, I1118_1456.port1=1, I1118_1458.port2=1, I1118_1459.port1=1, I1118_1460.port2=0, I1118_1463.port2=0, 
  (Signal Values: w_135_304=1, w_420_1439=0, w_510_260=0, w_560_1382=0, w_794_021=1, w_811_1380=1, w_916_191=0, )

37)
  Loop Signals: w_996_1460, w_996_1461, w_996_1462, w_996_1463, w_996_1464, w_996_1465, w_996_1466, w_996_1467, 
  Loop Gates: I996_1459.port1, I996_1460.port1, I996_1461.port1, I996_1462.port1, I996_1463.port2, I996_1464.port1, I996_1465.port2, I996_1466.port2, 
  Loop Conditions: I996_1459.port2=0, I996_1460.port2=0, I996_1463.port2=0, I996_1465.port1=0, I996_1466.port1=0, 
  (Signal Values: w_252_658=0, w_356_068=0, w_696_431=0, w_797_284=0, w_996_1464=0, )

38)
  Loop Signals: w_996_1465, w_996_1471, w_996_1472, w_996_1473, w_996_1474, w_996_1475, w_996_1476, w_996_1477, w_996_1478, w_996_1479, w_996_1480, w_996_1482, 
  Loop Gates: I996_1463.port1, I996_1467.port2, I996_1468.port1, I996_1469.port1, I996_1470.port1, I996_1471.port2, I996_1472.port1, I996_1473.port1, I996_1474.port1, I996_1475.port1, I996_1476.port1, I996_1477.port2, 
  Loop Conditions: I996_1463.port2=0, I996_1467.port1=1, I996_1469.port2=0, I996_1471.port1=1, I996_1473.port2=1, I996_1475.port2=0, I996_1477.port2=1, 
  (Signal Values: w_311_453=0, w_373_465=1, w_691_509=0, w_797_000=1, w_817_481=1, w_996_1464=0, w_996_1480=1, )

39)
  Loop Signals: w_399_1788, w_399_1789, w_399_1790, w_399_1791, w_399_1792, w_399_1793, w_399_1794, w_399_1795, w_399_1796, w_399_1797, w_399_1798, 
  Loop Gates: I399_1787.port1, I399_1788.port1, I399_1789.port2, I399_1790.port1, I399_1791.port1, I399_1792.port1, I399_1793.port1, I399_1794.port1, I399_1795.port1, I399_1796.port1, I399_1797.port1, 
  Loop Conditions: I399_1789.port2=1, I399_1791.port2=0, I399_1793.port2=0, I399_1797.port2=1, 
  (Signal Values: w_079_747=0, w_141_123=1, w_368_455=0, w_399_1790=1, )

40)
  Loop Signals: w_399_1791, w_399_1802, w_399_1803, w_399_1804, w_399_1806, 
  Loop Gates: I399_1789.port1, I399_1798.port1, I399_1799.port1, I399_1800.port1, I399_1801.port2, 
  Loop Conditions: I399_1789.port2=1, I399_1801.port2=1, 
  (Signal Values: w_399_1790=1, w_399_1804=1, )

41)
  Loop Signals: w_1112_1748, w_1112_1749, w_1112_1750, w_1112_1751, w_1112_1752, w_1112_1753, w_1112_1754, w_1112_1755, w_1112_1756, 
  Loop Gates: I1112_1747.port2, I1112_1748.port1, I1112_1749.port1, I1112_1750.port2, I1112_1751.port1, I1112_1752.port1, I1112_1753.port2, I1112_1754.port1, I1112_1755.port1, 
  Loop Conditions: I1112_1747.port1=1, I1112_1750.port1=1, I1112_1752.port2=1, I1112_1753.port1=1, I1112_1754.port2=0, I1112_1755.port2=1, 
  (Signal Values: w_057_632=1, w_276_134=0, w_499_436=1, w_591_1100=1, w_1055_134=1, w_1087_369=1, )

42)
  Loop Signals: w_1289_456, w_1289_457, w_1289_458, w_1289_459, w_1289_460, w_1289_461, w_1289_462, w_1289_463, 
  Loop Gates: I1289_456.port1, I1289_457.port1, I1289_458.port1, I1289_459.port1, I1289_460.port1, I1289_461.port2, I1289_462.port1, I1289_463.port2, 
  Loop Conditions: I1289_456.port2=1, I1289_458.port2=1, I1289_459.port2=0, I1289_461.port1=1, I1289_462.port2=1, I1289_463.port1=0, 
  (Signal Values: w_036_355=0, w_326_737=0, w_549_222=1, w_606_070=1, w_620_074=1, w_860_1045=1, )

43)
  Loop Signals: w_966_461, w_966_462, w_966_463, w_966_464, w_966_465, w_966_466, 
  Loop Gates: I966_460.port1, I966_461.port2, I966_462.port2, I966_463.port1, I966_464.port1, I966_465.port2, 
  Loop Conditions: I966_460.port2=1, I966_461.port1=1, I966_462.port1=0, I966_463.port2=1, I966_464.port2=1, I966_465.port1=1, 
  (Signal Values: w_032_140=1, w_267_432=1, w_487_1069=0, w_830_022=1, w_876_063=1, w_966_480=1, )

44)
  Loop Signals: w_966_462, w_966_470, w_966_471, w_966_472, w_966_473, w_966_474, w_966_475, w_966_476, w_966_477, w_966_478, w_966_480, 
  Loop Gates: I966_460.port2, I966_466.port1, I966_467.port2, I966_468.port1, I966_469.port1, I966_470.port1, I966_471.port1, I966_472.port1, I966_473.port2, I966_474.port1, I966_475.port2, 
  Loop Conditions: I966_460.port2=1, I966_466.port2=0, I966_467.port1=1, I966_468.port2=1, I966_469.port2=0, I966_470.port2=1, I966_471.port2=1, I966_472.port2=0, I966_473.port1=0, I966_475.port2=1, 
  (Signal Values: w_016_028=1, w_047_545=0, w_213_512=0, w_259_070=1, w_481_1485=0, w_510_180=0, w_512_268=1, w_690_753=1, w_966_478=1, w_966_480=1, )

45)
  Loop Signals: w_148_1915, w_148_1916, w_148_1917, w_148_1918, w_148_1919, w_148_1920, w_148_1921, w_148_1922, w_148_1923, w_148_1924, w_148_1925, 
  Loop Gates: I148_1914.port1, I148_1915.port1, I148_1916.port1, I148_1917.port2, I148_1918.port1, I148_1919.port1, I148_1920.port1, I148_1921.port2, I148_1922.port1, I148_1923.port1, I148_1924.port2, 
  Loop Conditions: I148_1916.port2=0, I148_1917.port1=1, I148_1919.port2=0, I148_1920.port2=1, I148_1921.port1=1, I148_1923.port2=1, I148_1924.port1=1, 
  (Signal Values: w_041_110=0, w_041_288=1, w_058_1347=0, w_075_187=1, w_110_905=1, w_137_417=1, w_139_1723=1, )

46)
  Loop Signals: w_1275_1436, w_1275_1444, w_1275_1445, w_1275_1446, w_1275_1447, w_1275_1448, w_1275_1449, w_1275_1450, w_1275_1451, w_1275_1452, w_1275_1453, w_1275_1454, w_1275_1456, 
  Loop Gates: I1275_1434.port2, I1275_1440.port1, I1275_1441.port1, I1275_1442.port2, I1275_1443.port1, I1275_1444.port1, I1275_1445.port1, I1275_1446.port1, I1275_1447.port1, I1275_1448.port2, I1275_1449.port1, I1275_1450.port1, I1275_1451.port2, 
  Loop Conditions: I1275_1434.port2=1, I1275_1440.port2=1, I1275_1441.port2=1, I1275_1442.port1=1, I1275_1443.port2=0, I1275_1446.port2=0, I1275_1447.port2=1, I1275_1448.port1=0, I1275_1451.port2=1, 
  (Signal Values: w_011_702=0, w_063_1040=1, w_421_269=0, w_504_152=1, w_626_1103=1, w_942_113=1, w_1246_814=0, w_1275_1454=1, w_1275_1456=1, )

47)
  Loop Signals: w_493_572, w_493_573, w_493_574, w_493_575, w_493_576, w_493_577, w_493_578, 
  Loop Gates: I493_571.port2, I493_572.port1, I493_573.port1, I493_574.port2, I493_575.port1, I493_576.port1, I493_577.port1, 
  Loop Conditions: I493_571.port2=1, I493_572.port2=1, I493_574.port1=1, I493_577.port2=1, 
  (Signal Values: w_262_184=1, w_349_104=1, w_476_312=1, w_493_572=1, )

48)
  Loop Signals: w_022_440, w_022_441, w_022_442, w_022_443, w_022_444, w_022_445, w_022_446, w_022_447, 
  Loop Gates: I022_439.port2, I022_440.port1, I022_441.port2, I022_442.port1, I022_443.port1, I022_444.port1, I022_445.port1, I022_446.port1, 
  Loop Conditions: I022_439.port1=1, I022_441.port1=1, I022_442.port2=1, I022_444.port2=1, I022_446.port2=1, 
  (Signal Values: w_003_271=1, w_009_009=1, w_010_322=1, w_011_011=1, w_018_200=1, )

49)
  Loop Signals: w_022_451, w_022_452, w_022_453, w_022_454, w_022_455, w_022_456, w_022_457, w_022_458, w_022_459, 
  Loop Gates: I022_447.port2, I022_448.port2, I022_449.port2, I022_450.port1, I022_451.port1, I022_452.port2, I022_453.port2, I022_454.port2, I022_455.port2, 
  Loop Conditions: I022_447.port1=1, I022_448.port1=1, I022_449.port1=1, I022_450.port2=0, I022_451.port2=1, I022_452.port1=1, I022_453.port1=0, I022_454.port1=1, I022_455.port1=0, 
  (Signal Values: w_003_289=0, w_003_319=0, w_010_135=1, w_010_295=0, w_011_256=1, w_013_302=1, w_015_048=1, w_017_1231=1, w_009_129=1, )

50)
  Loop Signals: w_722_1621, w_722_1622, w_722_1623, w_722_1624, w_722_1625, w_722_1626, w_722_1627, w_722_1628, 
  Loop Gates: I722_1620.port2, I722_1621.port2, I722_1622.port2, I722_1623.port1, I722_1624.port2, I722_1625.port1, I722_1626.port1, I722_1627.port2, 
  Loop Conditions: I722_1620.port1=1, I722_1621.port1=1, I722_1622.port1=0, I722_1624.port1=1, I722_1625.port2=1, I722_1626.port2=0, I722_1627.port1=0, 
  (Signal Values: w_184_004=0, w_246_1608=0, w_298_828=1, w_316_915=1, w_320_484=0, w_611_122=1, w_670_353=1, )

******* result_4.txt *********
1)
  Loop Breaker: I894_590.port0-w_894_586-Register-w_894_586'-I894_585.port1 

2)
  Loop Breaker: I894_590.port0-w_894_586-Register-w_894_586'-I894_601.port1 

3)
  Loop Breaker: I102_1263.port0-w_102_1259-Register-w_102_1259'-I102_1258.port1 

4)
  Loop Breaker: I102_1263.port0-w_102_1259-Register-w_102_1259'-I102_1272.port1 

5)
  Loop Breaker: I799_853.port0-w_799_855-Register-w_799_855'-I799_854.port1 

6)
  Loop Breaker: I811_1657.port0-w_811_1656-Register-w_811_1656'-I811_1664.port1 

7)
  Loop Breaker: I432_730.port0-w_432_726-Register-w_432_726'-I432_735.port1 

8)
  Loop Breaker: I1692_767.port0-w_1692_769-Register-w_1692_769'-I1692_776.port1 

9)
  Loop Breaker: I1298_519.port0-w_1298_518-Register-w_1298_518'-I1298_523.port1 

10)
  Loop Breaker: I610_888.port0-w_610_890-Register-w_610_890'-I610_889.port1 

11)
  Loop Breaker: I1230_964.port0-w_1230_966-Register-w_1230_966'-I1230_965.port1 

12)
  Loop Breaker: I1288_1602.port0-w_1288_1604-Register-w_1288_1604'-I1288_1603.port2 

13)
  Loop Breaker: I826_438.port0-w_826_440-Register-w_826_440'-I826_439.port1 

14)
  Loop Breaker: I826_438.port0-w_826_440-Register-w_826_440'-I826_446.port1 

15)
  Loop Breaker: I1132_1116.port0-w_1132_1118-Register-w_1132_1118'-I1132_1117.port1 

16)
  Loop Breaker: I1449_505.port0-w_1449_507-Register-w_1449_507'-I1449_506.port2 

17)
  Loop Breaker: I1308_360.port0-w_1308_362-Register-w_1308_362'-I1308_361.port1 

18)
  Loop Breaker: I1308_360.port0-w_1308_362-Register-w_1308_362'-I1308_378.port1 

19)
  Loop Breaker: I531_1386.port0-w_531_1388-Register-w_531_1388'-I531_1391.port1 

20)
  Loop Breaker: I1821_249.port0-w_1821_251-Register-w_1821_251'-I1821_250.port1 

21)
  Loop Breaker: I1821_249.port0-w_1821_251-Register-w_1821_251'-I1821_262.port1 

22)
  Loop Breaker: I1601_113.port0-w_1601_115-Register-w_1601_115'-I1601_121.port1 

23)
  Loop Breaker: I305_017.port0-w_305_019-Register-w_305_019'-I305_018.port1 

24)
  Loop Breaker: I1911_1095.port0-w_1911_1097-Register-w_1911_1097'-I1911_1096.port1 

25)
  Loop Breaker: I299_1758.port0-w_299_1760-Register-w_299_1760'-I299_1759.port2 

26)
  Loop Breaker: I1075_1908.port0-w_1075_1910-Register-w_1075_1910'-I1075_1909.port1 

27)
  Loop Breaker: I1075_1908.port0-w_1075_1910-Register-w_1075_1910'-I1075_1918.port1 

28)
  Loop Breaker: I897_1328.port0-w_897_1330-Register-w_897_1330'-I897_1329.port1 

29)
  Loop Breaker: I116_1548.port0-w_116_1550-Register-w_116_1550'-I116_1549.port1 

30)
  Loop Breaker: I116_1548.port0-w_116_1550-Register-w_116_1550'-I116_1568.port1 

31)
  Loop Breaker: I110_1610.port0-w_110_1612-Register-w_110_1612'-I110_1611.port1 

32)
  Loop Breaker: I1312_979.port0-w_1312_969-Register-w_1312_969'-I1312_982.port1 

33)
  Loop Breaker: I976_293.port0-w_976_295-Register-w_976_295'-I976_294.port2 

34)
  Loop Breaker: I976_293.port0-w_976_295-Register-w_976_295'-I976_297.port1 

35)
  Loop Breaker: I1078_080.port0-w_1078_082-Register-w_1078_082'-I1078_081.port2 

36)
  Loop Breaker: I1118_1454.port0-w_1118_1456-Register-w_1118_1456'-I1118_1455.port1 

37)
  Loop Breaker: I996_1463.port0-w_996_1465-Register-w_996_1465'-I996_1464.port1 

38)
  Loop Breaker: I996_1463.port0-w_996_1465-Register-w_996_1465'-I996_1476.port1 

39)
  Loop Breaker: I399_1789.port0-w_399_1791-Register-w_399_1791'-I399_1790.port1 

40)
  Loop Breaker: I399_1789.port0-w_399_1791-Register-w_399_1791'-I399_1800.port1 

41)
  Loop Breaker: I1112_1747.port0-w_1112_1749-Register-w_1112_1749'-I1112_1748.port1 

42)
  Loop Breaker: I1289_456.port0-w_1289_457-Register-w_1289_457'-I1289_457.port1 

43)
  Loop Breaker: I966_460.port0-w_966_462-Register-w_966_462'-I966_461.port2 

44)
  Loop Breaker: I966_460.port0-w_966_462-Register-w_966_462'-I966_474.port1 

45)
  Loop Breaker: I148_1914.port0-w_148_1916-Register-w_148_1916'-I148_1915.port1 

46)
  Loop Breaker: I1275_1434.port0-w_1275_1436-Register-w_1275_1436'-I1275_1450.port1 

47)
  Loop Breaker: I493_571.port0-w_493_573-Register-w_493_573'-I493_572.port1 

48)
  Loop Breaker: I022_439.port0-w_022_441-Register-w_022_441'-I022_440.port1 

49)
  Loop Breaker: I022_447.port0-w_022_452-Register-w_022_452'-I022_448.port2 

50)
  Loop Breaker: I722_1620.port0-w_722_1622-Register-w_722_1622'-I722_1621.port2 

// ******* The results for this case End *********
*/

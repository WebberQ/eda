// ****** Basic Gate Module Defination ******
module or2(out, in1, in2);
  output out;
  input in1, in2;
  wire in1, in2, out;
  assign out = in1 || in2;
endmodule

module and2(out, in1, in2);
  output out;
  input in1, in2;
  wire in1, in2, out;
  assign out = in1 && in2;
endmodule

module not1(out, in);
  output out;
  input in;
  wire in,out;
  assign out = ~in;
endmodule

module nand2(out, in1, in2);
  output out;
  input in1, in2;
  wire in1, in2, out;
  assign out = ~(in1 && in2);
endmodule
// ****** Basic Gate Module Defination End ******

// ****** Combined Logic Module Defination ******
module combLogic( w_000_000, w_000_001, w_000_002, w_000_003, w_000_004, w_000_005, w_000_006, w_000_007, w_000_008, w_000_009, w_000_010, w_000_011, w_000_012, w_000_013, w_000_014, w_000_015, w_000_016, w_000_017, w_000_018, w_000_019, w_000_020, w_000_021, w_000_022, w_000_023, w_000_024, w_000_025, w_000_026, w_000_027, w_000_028, w_000_029, w_000_030, w_000_031, w_000_032, w_000_033, w_000_034, w_000_035, w_000_036, w_000_037, w_000_038, w_000_039, w_000_040, w_000_041, w_000_042, w_000_043, w_000_044, w_000_045, w_000_046, w_000_047, w_000_048, w_000_050, w_000_051, w_000_053, w_000_054, w_000_055, w_000_056, w_000_057, w_000_058, w_000_059, w_000_060, w_000_061, w_000_064, w_000_065, w_000_066, w_000_067, w_000_068, w_000_069, w_000_070, w_000_071, w_000_072, w_000_073, w_000_074, w_000_075, w_080_000, w_080_001, w_080_002, w_080_003, w_080_004 );
  inout w_000_000, w_000_001, w_000_002, w_000_003, w_000_004, w_000_005, w_000_006, w_000_007, w_000_008, w_000_009, w_000_010, w_000_011, w_000_012, w_000_013, w_000_014, w_000_015, w_000_016, w_000_017, w_000_018, w_000_019, w_000_020, w_000_021, w_000_022, w_000_023, w_000_024, w_000_025, w_000_026, w_000_027, w_000_028, w_000_029, w_000_030, w_000_031, w_000_032, w_000_033, w_000_034, w_000_035, w_000_036, w_000_037, w_000_038, w_000_039, w_000_040, w_000_041, w_000_042, w_000_043, w_000_044, w_000_045, w_000_046, w_000_047, w_000_048, w_000_050, w_000_051, w_000_053, w_000_054, w_000_055, w_000_056, w_000_057, w_000_058, w_000_059, w_000_060, w_000_061, w_000_064, w_000_065, w_000_066, w_000_067, w_000_068, w_000_069, w_000_070, w_000_071, w_000_072, w_000_073, w_000_074, w_000_075;
  output w_080_000, w_080_001, w_080_002, w_080_003, w_080_004;
  wire w_000_000, w_000_001, w_000_002, w_000_003, w_000_004, w_000_005, w_000_006, w_000_007, w_000_008, w_000_009, w_000_010, w_000_011, w_000_012, w_000_013, w_000_014, w_000_015, w_000_016, w_000_017, w_000_018, w_000_019, w_000_020, w_000_021, w_000_022, w_000_023, w_000_024, w_000_025, w_000_026, w_000_027, w_000_028, w_000_029, w_000_030, w_000_031, w_000_032, w_000_033, w_000_034, w_000_035, w_000_036, w_000_037, w_000_038, w_000_039, w_000_040, w_000_041, w_000_042, w_000_043, w_000_044, w_000_045, w_000_046, w_000_047, w_000_048, w_000_050, w_000_051, w_000_053, w_000_054, w_000_055, w_000_056, w_000_057, w_000_058, w_000_059, w_000_060, w_000_061, w_000_064, w_000_065, w_000_066, w_000_067, w_000_068, w_000_069, w_000_070, w_000_071, w_000_072, w_000_073, w_000_074, w_000_075;
  wire w_001_000, w_001_001, w_001_002, w_001_003, w_001_004, w_001_005, w_001_007, w_001_008, w_001_009, w_001_010, w_001_011, w_001_012, w_001_013, w_001_014, w_001_015, w_001_016, w_001_017, w_001_018, w_001_019, w_001_020, w_001_021, w_001_022, w_001_024, w_001_025, w_001_026, w_001_027, w_001_028, w_001_029, w_001_030, w_001_031, w_001_032, w_001_033, w_001_034, w_001_035, w_001_037, w_001_040, w_001_041, w_001_042, w_001_043, w_001_044;
  wire w_002_000, w_002_001, w_002_004, w_002_005, w_002_006, w_002_007, w_002_010, w_002_011, w_002_012, w_002_013, w_002_014, w_002_017, w_002_018, w_002_019, w_002_020, w_002_021, w_002_022, w_002_023, w_002_024, w_002_026, w_002_027, w_002_028, w_002_030, w_002_033, w_002_036, w_002_037, w_002_038, w_002_039, w_002_040, w_002_041, w_002_042, w_002_043, w_002_046, w_002_047, w_002_048, w_002_050, w_002_051, w_002_052, w_002_055, w_002_056, w_002_057, w_002_058, w_002_060, w_002_061, w_002_065;
  wire w_003_000, w_003_001, w_003_002, w_003_003, w_003_004, w_003_006, w_003_007, w_003_008, w_003_009, w_003_010, w_003_011, w_003_013, w_003_015, w_003_016, w_003_017, w_003_018, w_003_019, w_003_021, w_003_022, w_003_024, w_003_025, w_003_026, w_003_030, w_003_031, w_003_033, w_003_034, w_003_040, w_003_043, w_003_044, w_003_045;
  wire w_004_000, w_004_001, w_004_002, w_004_004, w_004_006, w_004_009, w_004_010, w_004_011, w_004_012, w_004_013, w_004_014, w_004_015, w_004_017, w_004_018, w_004_019, w_004_020, w_004_021, w_004_023, w_004_024, w_004_026, w_004_027, w_004_028;
  wire w_005_000, w_005_001, w_005_002, w_005_003, w_005_005, w_005_008, w_005_009, w_005_010, w_005_011, w_005_012, w_005_013, w_005_015, w_005_016, w_005_017, w_005_018, w_005_022, w_005_024, w_005_025, w_005_026, w_005_027, w_005_028, w_005_030, w_005_031, w_005_033;
  wire w_006_000;
  wire w_007_000, w_007_001, w_007_002, w_007_003, w_007_004, w_007_005, w_007_006, w_007_009, w_007_010, w_007_012, w_007_013, w_007_015, w_007_016, w_007_017, w_007_018, w_007_019;
  wire w_008_000, w_008_003, w_008_004, w_008_006, w_008_009, w_008_010, w_008_011, w_008_013, w_008_016, w_008_019, w_008_023, w_008_026, w_008_027, w_008_030, w_008_031, w_008_032, w_008_033;
  wire w_009_000, w_009_001, w_009_002, w_009_003, w_009_004, w_009_005, w_009_008, w_009_009, w_009_011;
  wire w_010_000, w_010_001, w_010_002, w_010_004, w_010_008, w_010_009, w_010_014, w_010_015, w_010_016, w_010_018, w_010_019;
  wire w_011_001, w_011_003, w_011_004, w_011_010, w_011_013, w_011_014, w_011_015, w_011_016, w_011_017, w_011_018, w_011_019, w_011_021, w_011_023, w_011_024;
  wire w_012_000, w_012_010, w_012_014, w_012_023, w_012_024, w_012_025, w_012_030, w_012_034, w_012_039, w_012_045, w_012_046, w_012_049, w_012_050, w_012_059, w_012_060, w_012_061, w_012_062, w_012_063, w_012_064, w_012_065, w_012_066, w_012_067, w_012_068;
  wire w_013_014, w_013_015, w_013_020, w_013_041, w_013_042, w_013_052, w_013_058, w_013_067;
  wire w_014_007, w_014_014, w_014_019, w_014_021, w_014_031;
  wire w_015_001, w_015_002, w_015_003, w_015_005, w_015_006, w_015_007, w_015_008;
  wire w_016_004, w_016_005, w_016_006, w_016_007, w_016_009, w_016_014, w_016_015, w_016_017, w_016_018, w_016_020, w_016_022;
  wire w_017_007, w_017_013, w_017_020, w_017_023, w_017_026, w_017_046, w_017_057, w_017_064, w_017_067, w_017_070;
  wire w_018_001, w_018_002, w_018_005, w_018_006, w_018_012, w_018_030, w_018_036, w_018_049, w_018_055;
  wire w_019_000;
  wire w_020_024, w_020_027, w_020_038, w_020_046, w_020_053, w_020_056, w_020_057, w_020_059, w_020_060, w_020_061, w_020_062, w_020_063, w_020_064, w_020_065, w_020_066, w_020_067, w_020_069, w_020_071, w_020_072, w_020_073, w_020_074, w_020_075, w_020_076, w_020_077, w_020_078, w_020_079, w_020_080, w_020_081, w_020_083, w_020_085;
  wire w_021_000, w_021_009, w_021_010, w_021_011, w_021_014, w_021_015;
  wire w_022_000, w_022_001, w_022_004, w_022_007, w_022_008, w_022_010, w_022_011, w_022_012, w_022_014, w_022_017, w_022_023, w_022_024, w_022_025, w_022_026, w_022_027, w_022_028, w_022_029, w_022_030, w_022_031, w_022_032, w_022_033, w_022_034, w_022_036, w_022_038, w_022_039, w_022_040, w_022_041, w_022_042, w_022_043, w_022_045, w_022_047, w_022_049;
  wire w_023_000, w_023_001, w_023_002, w_023_004;
  wire w_024_002, w_024_018, w_024_031, w_024_032, w_024_033, w_024_034, w_024_038, w_024_039, w_024_040, w_024_041, w_024_042, w_024_043, w_024_044, w_024_045, w_024_047;
  wire w_025_005, w_025_050;
  wire w_026_026, w_026_046;
  wire w_027_011, w_027_015, w_027_016;
  wire w_029_006, w_029_013, w_029_019;
  wire w_030_030;
  wire w_031_025, w_031_028, w_031_034, w_031_038;
  wire w_033_002, w_033_003, w_033_004, w_033_005, w_033_006, w_033_009;
  wire w_034_023, w_034_030, w_034_071;
  wire w_036_000;
  wire w_037_008, w_037_055, w_037_074, w_037_075, w_037_076, w_037_077, w_037_078, w_037_079;
  wire w_038_038, w_038_062, w_038_081, w_038_082, w_038_083, w_038_084, w_038_088, w_038_089, w_038_090, w_038_091, w_038_093;
  wire w_039_023, w_039_024, w_039_029;
  wire w_040_001;
  wire w_041_002, w_041_008;
  wire w_042_002, w_042_007;
  wire w_043_000;
  wire w_044_004, w_044_006, w_044_007, w_044_010;
  wire w_047_008, w_047_030, w_047_038, w_047_045, w_047_058;
  wire w_048_031, w_048_042, w_048_043, w_048_044, w_048_045, w_048_046, w_048_047, w_048_048, w_048_049, w_048_050, w_048_051, w_048_052, w_048_056, w_048_057, w_048_058, w_048_060;
  wire w_049_001;
  wire w_050_017;
  wire w_051_000, w_051_001, w_051_024, w_051_025, w_051_026, w_051_027, w_051_028, w_051_029, w_051_030, w_051_031, w_051_032;
  wire w_052_026, w_052_027, w_052_028, w_052_029, w_052_030, w_052_031, w_052_032, w_052_033, w_052_034, w_052_038, w_052_039, w_052_040, w_052_041, w_052_042, w_052_044;
  wire w_054_015, w_054_035;
  wire w_055_018;
  wire w_056_039;
  wire w_057_029, w_057_063, w_057_064, w_057_065;
  wire w_060_016;
  wire w_061_014, w_061_023;
  wire w_062_003;
  wire w_064_008, w_064_024;
  wire w_065_034, w_065_035, w_065_036, w_065_037, w_065_038, w_065_039, w_065_040, w_065_041, w_065_042, w_065_043, w_065_044, w_065_045, w_065_049, w_065_050, w_065_051, w_065_052, w_065_053, w_065_054, w_065_055, w_065_056, w_065_057, w_065_059;
  wire w_069_000;
  wire w_075_004;
  wire w_076_002, w_076_033, w_076_034, w_076_035, w_076_036, w_076_037, w_076_038, w_076_039, w_076_043, w_076_044, w_076_045, w_076_046, w_076_047, w_076_048, w_076_049, w_076_050, w_076_051, w_076_052, w_076_054;
  wire w_077_000;
  wire w_080_000, w_080_001, w_080_002, w_080_003, w_080_004;
  not1 I001_000(w_001_000, w_000_000);
  nand2 I001_001(w_001_001, w_000_001, w_000_002);
  not1 I001_002(w_001_002, w_000_003);
  or2  I001_003(w_001_003, w_000_004, w_000_005);
  nand2 I001_004(w_001_004, w_000_006, w_000_007);
  nand2 I001_005(w_001_005, w_000_006, w_000_008);
  and2 I001_007(w_001_007, w_000_010, w_000_008);
  nand2 I001_008(w_001_008, w_000_011, w_000_012);
  not1 I001_009(w_001_009, w_000_013);
  nand2 I001_010(w_001_010, w_000_014, w_000_015);
  or2  I001_011(w_001_011, w_000_016, w_000_017);
  not1 I001_012(w_001_012, w_000_018);
  nand2 I001_013(w_001_013, w_000_019, w_000_020);
  nand2 I001_014(w_001_014, w_000_021, w_000_022);
  or2  I001_015(w_001_015, w_000_021, w_000_023);
  and2 I001_016(w_001_016, w_000_024, w_000_025);
  and2 I001_017(w_001_017, w_000_026, w_000_027);
  or2  I001_018(w_001_018, w_000_006, w_000_011);
  and2 I001_019(w_001_019, w_000_028, w_000_029);
  not1 I001_020(w_001_020, w_000_030);
  and2 I001_021(w_001_021, w_000_001, w_000_031);
  or2  I001_022(w_001_022, w_000_032, w_000_007);
  or2  I001_024(w_001_024, w_000_033, w_000_017);
  and2 I001_025(w_001_025, w_000_034, w_000_035);
  or2  I001_026(w_001_026, w_000_014, w_000_007);
  not1 I001_027(w_001_027, w_000_036);
  nand2 I001_028(w_001_028, w_000_037, w_000_038);
  and2 I001_029(w_001_029, w_000_039, w_000_040);
  and2 I001_030(w_001_030, w_000_041, w_000_042);
  nand2 I001_031(w_001_031, w_000_034, w_000_043);
  and2 I001_032(w_001_032, w_000_020, w_000_044);
  and2 I001_033(w_001_033, w_000_045, w_000_012);
  not1 I001_034(w_001_034, w_000_026);
  not1 I001_035(w_001_035, w_000_019);
  not1 I001_037(w_001_037, w_000_027);
  or2  I001_040(w_001_040, w_000_040, w_000_046);
  or2  I001_041(w_001_041, w_000_025, w_000_009);
  and2 I001_042(w_001_042, w_000_047, w_000_040);
  or2  I001_043(w_001_043, w_000_031, w_000_037);
  or2  I001_044(w_001_044, w_000_011, w_000_001);
  and2 I002_000(w_002_000, w_001_033, w_000_005);
  not1 I002_001(w_002_001, w_001_013);
  nand2 I002_004(w_002_004, w_000_050, w_000_003);
  not1 I002_005(w_002_005, w_001_000);
  nand2 I002_006(w_002_006, w_001_035, w_001_002);
  and2 I002_007(w_002_007, w_000_001, w_000_051);
  or2  I002_010(w_002_010, w_001_016, w_000_053);
  or2  I002_011(w_002_011, w_000_054, w_001_034);
  or2  I002_012(w_002_012, w_000_055, w_001_037);
  nand2 I002_013(w_002_013, w_001_012, w_000_056);
  nand2 I002_014(w_002_014, w_000_009, w_000_004);
  or2  I002_017(w_002_017, w_001_031, w_000_044);
  nand2 I002_018(w_002_018, w_000_023, w_000_057);
  and2 I002_019(w_002_019, w_001_044, w_000_058);
  nand2 I002_020(w_002_020, w_000_026, w_001_002);
  not1 I002_021(w_002_021, w_000_037);
  nand2 I002_022(w_002_022, w_001_004, w_000_051);
  not1 I002_023(w_002_023, w_000_019);
  nand2 I002_024(w_002_024, w_000_048, w_000_059);
  not1 I002_026(w_002_026, w_000_025);
  and2 I002_027(w_002_027, w_000_004, w_000_042);
  or2  I002_028(w_002_028, w_000_056, w_000_058);
  and2 I002_030(w_002_030, w_000_059, w_001_030);
  and2 I002_033(w_002_033, w_001_033, w_001_019);
  not1 I002_036(w_002_036, w_000_060);
  not1 I002_037(w_002_037, w_000_016);
  not1 I002_038(w_002_038, w_000_061);
  or2  I002_039(w_002_039, w_000_059, w_000_007);
  and2 I002_040(w_002_040, w_000_012, w_001_009);
  and2 I002_041(w_002_041, w_000_022, w_001_000);
  or2  I002_042(w_002_042, w_001_012, w_001_009);
  nand2 I002_043(w_002_043, w_001_041, w_000_019);
  and2 I002_046(w_002_046, w_000_064, w_000_001);
  not1 I002_047(w_002_047, w_000_012);
  and2 I002_048(w_002_048, w_000_010, w_001_025);
  not1 I002_050(w_002_050, w_000_065);
  not1 I002_051(w_002_051, w_000_044);
  not1 I002_052(w_002_052, w_001_021);
  not1 I002_055(w_002_055, w_001_020);
  not1 I002_056(w_002_056, w_001_044);
  or2  I002_057(w_002_057, w_001_021, w_001_024);
  or2  I002_058(w_002_058, w_001_034, w_000_019);
  or2  I002_060(w_002_060, w_000_066, w_000_067);
  and2 I002_061(w_002_061, w_000_038, w_000_036);
  and2 I002_065(w_002_065, w_000_028, w_001_009);
  nand2 I003_000(w_003_000, w_001_003, w_002_013);
  and2 I003_001(w_003_001, w_000_005, w_002_010);
  nand2 I003_002(w_003_002, w_002_037, w_000_068);
  and2 I003_003(w_003_003, w_002_001, w_000_064);
  and2 I003_004(w_003_004, w_001_004, w_002_036);
  nand2 I003_006(w_003_006, w_001_033, w_002_028);
  nand2 I003_007(w_003_007, w_002_041, w_002_058);
  nand2 I003_008(w_003_008, w_002_055, w_002_019);
  and2 I003_009(w_003_009, w_000_047, w_000_029);
  or2  I003_010(w_003_010, w_000_045, w_001_017);
  nand2 I003_011(w_003_011, w_000_020, w_001_005);
  nand2 I003_013(w_003_013, w_002_024, w_000_069);
  or2  I003_015(w_003_015, w_002_006, w_002_042);
  and2 I003_016(w_003_016, w_000_023, w_002_001);
  or2  I003_017(w_003_017, w_000_065, w_002_047);
  or2  I003_018(w_003_018, w_000_050, w_001_044);
  or2  I003_019(w_003_019, w_002_048, w_000_038);
  not1 I003_021(w_003_021, w_001_026);
  not1 I003_022(w_003_022, w_001_020);
  nand2 I003_024(w_003_024, w_000_031, w_001_011);
  nand2 I003_025(w_003_025, w_002_046, w_000_035);
  and2 I003_026(w_003_026, w_002_012, w_000_010);
  and2 I003_030(w_003_030, w_000_046, w_001_009);
  or2  I003_031(w_003_031, w_000_019, w_002_038);
  or2  I003_033(w_003_033, w_000_003, w_001_032);
  or2  I003_034(w_003_034, w_001_025, w_000_060);
  nand2 I003_040(w_003_040, w_001_042, w_002_052);
  nand2 I003_043(w_003_043, w_000_061, w_002_060);
  not1 I003_044(w_003_044, w_002_018);
  or2  I003_045(w_003_045, w_001_030, w_001_042);
  nand2 I004_000(w_004_000, w_000_044, w_002_020);
  not1 I004_001(w_004_001, w_001_004);
  not1 I004_002(w_004_002, w_000_019);
  nand2 I004_004(w_004_004, w_003_033, w_001_018);
  and2 I004_006(w_004_006, w_002_065, w_003_003);
  or2  I004_009(w_004_009, w_002_005, w_002_022);
  not1 I004_010(w_004_010, w_001_030);
  or2  I004_011(w_004_011, w_002_046, w_001_000);
  or2  I004_012(w_004_012, w_003_034, w_002_007);
  nand2 I004_013(w_004_013, w_001_042, w_003_002);
  nand2 I004_014(w_004_014, w_002_012, w_002_057);
  not1 I004_015(w_004_015, w_003_017);
  or2  I004_017(w_004_017, w_003_024, w_002_017);
  and2 I004_018(w_004_018, w_003_015, w_002_018);
  not1 I004_019(w_004_019, w_000_011);
  or2  I004_020(w_004_020, w_001_005, w_001_033);
  and2 I004_021(w_004_021, w_003_045, w_002_028);
  or2  I004_023(w_004_023, w_000_007, w_002_043);
  or2  I004_024(w_004_024, w_000_061, w_001_040);
  not1 I004_026(w_004_026, w_000_071);
  nand2 I004_027(w_004_027, w_001_030, w_000_012);
  nand2 I004_028(w_004_028, w_002_040, w_003_026);
  not1 I005_000(w_005_000, w_000_013);
  not1 I005_001(w_005_001, w_004_002);
  nand2 I005_002(w_005_002, w_004_012, w_000_032);
  and2 I005_003(w_005_003, w_004_013, w_003_000);
  nand2 I005_005(w_005_005, w_001_008, w_003_004);
  or2  I005_008(w_005_008, w_003_015, w_003_013);
  or2  I005_009(w_005_009, w_002_039, w_003_006);
  or2  I005_010(w_005_010, w_000_044, w_003_008);
  not1 I005_011(w_005_011, w_001_010);
  not1 I005_012(w_005_012, w_000_012);
  nand2 I005_013(w_005_013, w_004_009, w_001_010);
  not1 I005_015(w_005_015, w_004_013);
  or2  I005_016(w_005_016, w_004_028, w_004_006);
  nand2 I005_017(w_005_017, w_002_023, w_002_005);
  and2 I005_018(w_005_018, w_002_001, w_000_050);
  nand2 I005_022(w_005_022, w_000_016, w_000_044);
  or2  I005_024(w_005_024, w_002_014, w_001_026);
  nand2 I005_025(w_005_025, w_002_028, w_000_072);
  not1 I005_026(w_005_026, w_002_043);
  and2 I005_027(w_005_027, w_004_017, w_004_027);
  and2 I005_028(w_005_028, w_002_061, w_001_043);
  or2  I005_030(w_005_030, w_000_070, w_003_034);
  and2 I005_031(w_005_031, w_001_014, w_002_005);
  and2 I005_033(w_005_033, w_003_043, w_002_048);
  and2 I006_000(w_006_000, w_005_015, w_004_017);
  and2 I007_000(w_007_000, w_004_023, w_001_017);
  or2  I007_001(w_007_001, w_004_006, w_004_011);
  nand2 I007_002(w_007_002, w_000_030, w_000_073);
  not1 I007_003(w_007_003, w_005_015);
  or2  I007_004(w_007_004, w_004_020, w_001_033);
  and2 I007_005(w_007_005, w_003_007, w_004_019);
  or2  I007_006(w_007_006, w_005_002, w_001_001);
  and2 I007_009(w_007_009, w_001_027, w_005_002);
  nand2 I007_010(w_007_010, w_006_000, w_005_005);
  not1 I007_012(w_007_012, w_005_018);
  not1 I007_013(w_007_013, w_000_054);
  or2  I007_015(w_007_015, w_005_012, w_002_036);
  and2 I007_016(w_007_016, w_004_002, w_005_009);
  or2  I007_017(w_007_017, w_004_023, w_000_026);
  nand2 I007_018(w_007_018, w_001_024, w_005_011);
  and2 I007_019(w_007_019, w_002_017, w_000_028);
  and2 I008_000(w_008_000, w_003_016, w_006_000);
  nand2 I008_003(w_008_003, w_000_020, w_002_038);
  nand2 I008_004(w_008_004, w_004_019, w_000_074);
  not1 I008_006(w_008_006, w_001_030);
  not1 I008_009(w_008_009, w_006_000);
  nand2 I008_010(w_008_010, w_001_015, w_000_061);
  or2  I008_011(w_008_011, w_006_000, w_005_031);
  or2  I008_013(w_008_013, w_001_033, w_006_000);
  not1 I008_016(w_008_016, w_005_025);
  nand2 I008_019(w_008_019, w_004_012, w_000_019);
  not1 I008_023(w_008_023, w_003_007);
  and2 I008_026(w_008_026, w_007_017, w_007_012);
  or2  I008_027(w_008_027, w_005_022, w_005_013);
  or2  I008_030(w_008_030, w_005_028, w_001_030);
  or2  I008_031(w_008_031, w_007_018, w_000_002);
  and2 I008_032(w_008_032, w_007_000, w_001_022);
  not1 I008_033(w_008_033, w_000_006);
  not1 I009_000(w_009_000, w_005_030);
  not1 I009_001(w_009_001, w_005_031);
  not1 I009_002(w_009_002, w_001_015);
  nand2 I009_003(w_009_003, w_006_000, w_004_018);
  not1 I009_004(w_009_004, w_003_009);
  and2 I009_005(w_009_005, w_008_030, w_008_027);
  not1 I009_008(w_009_008, w_004_009);
  nand2 I009_009(w_009_009, w_000_041, w_003_034);
  nand2 I009_011(w_009_011, w_006_000, w_004_004);
  nand2 I010_000(w_010_000, w_009_003, w_008_033);
  and2 I010_001(w_010_001, w_009_005, w_004_013);
  nand2 I010_002(w_010_002, w_004_019, w_005_000);
  not1 I010_004(w_010_004, w_007_002);
  nand2 I010_008(w_010_008, w_001_008, w_008_011);
  and2 I010_009(w_010_009, w_005_002, w_007_019);
  or2  I010_014(w_010_014, w_003_044, w_007_012);
  nand2 I010_015(w_010_015, w_007_009, w_005_001);
  and2 I010_016(w_010_016, w_009_005, w_005_027);
  and2 I010_018(w_010_018, w_002_011, w_000_045);
  nand2 I010_019(w_010_019, w_002_051, w_009_011);
  and2 I011_001(w_011_001, w_006_000, w_008_030);
  or2  I011_003(w_011_003, w_002_013, w_008_023);
  not1 I011_004(w_011_004, w_006_000);
  not1 I011_010(w_011_010, w_003_031);
  not1 I011_013(w_011_013, w_004_014);
  or2  I011_014(w_011_014, w_002_039, w_003_010);
  and2 I011_015(w_011_015, w_002_036, w_000_070);
  or2  I011_016(w_011_016, w_004_015, w_002_027);
  or2  I011_017(w_011_017, w_005_010, w_004_000);
  and2 I011_018(w_011_018, w_005_003, w_008_016);
  or2  I011_019(w_011_019, w_006_000, w_001_043);
  nand2 I011_021(w_011_021, w_007_009, w_007_010);
  or2  I011_023(w_011_023, w_009_011, w_002_007);
  and2 I011_024(w_011_024, w_000_041, w_005_011);
  and2 I012_000(w_012_000, w_003_008, w_011_023);
  nand2 I012_010(w_012_010, w_010_009, w_010_001);
  or2  I012_014(w_012_014, w_009_008, w_005_008);
  not1 I012_023(w_012_023, w_004_020);
  and2 I012_024(w_012_024, w_010_018, w_001_034);
  nand2 I012_025(w_012_025, w_002_026, w_004_013);
  or2  I012_030(w_012_030, w_007_016, w_005_028);
  not1 I012_034(w_012_034, w_002_030);
  not1 I012_039(w_012_039, w_002_004);
  nand2 I012_045(w_012_045, w_004_011, w_003_021);
  or2  I012_046(w_012_046, w_004_013, w_011_001);
  or2  I012_049(w_012_049, w_008_031, w_010_015);
  or2  I012_050(w_012_050, w_002_017, w_000_029);
  and2 I012_058(w_012_060, w_004_001, w_012_059);
  or2  I012_059(w_012_061, w_012_060, w_005_011);
  and2 I012_060(w_012_062, w_002_056, w_012_061);
  and2 I012_061(w_012_063, w_012_062, w_007_012);
  and2 I012_062(w_012_064, w_012_063, w_005_033);
  nand2 I012_063(w_012_065, w_006_000, w_012_064);
  not1 I012_064(w_012_066, w_012_065);
  or2  I012_065(w_012_067, w_012_066, w_005_000);
  and2 I012_066(w_012_068, w_012_067, w_003_016);
  not1 I012_067(w_012_059, w_012_068);
  nand2 I013_014(w_013_014, w_001_043, w_008_000);
  and2 I013_015(w_013_015, w_012_014, w_000_024);
  or2  I013_020(w_013_020, w_010_000, w_008_030);
  not1 I013_041(w_013_041, w_012_045);
  or2  I013_042(w_013_042, w_000_042, w_008_032);
  not1 I013_052(w_013_052, w_012_023);
  or2  I013_058(w_013_058, w_005_016, w_009_001);
  not1 I013_067(w_013_067, w_003_030);
  nand2 I014_007(w_014_007, w_010_009, w_009_000);
  not1 I014_014(w_014_014, w_010_019);
  nand2 I014_019(w_014_019, w_006_000, w_005_027);
  nand2 I014_021(w_014_021, w_000_075, w_013_014);
  and2 I014_031(w_014_031, w_012_024, w_000_055);
  or2  I015_001(w_015_001, w_004_024, w_013_052);
  nand2 I015_002(w_015_002, w_006_000, w_002_056);
  and2 I015_003(w_015_003, w_006_000, w_011_018);
  or2  I015_005(w_015_005, w_010_014, w_014_031);
  not1 I015_006(w_015_006, w_000_045);
  or2  I015_007(w_015_007, w_004_011, w_005_005);
  and2 I015_008(w_015_008, w_009_004, w_007_004);
  and2 I016_004(w_016_004, w_002_021, w_003_001);
  not1 I016_005(w_016_005, w_008_006);
  or2  I016_006(w_016_006, w_011_013, w_005_024);
  nand2 I016_007(w_016_007, w_004_015, w_010_002);
  not1 I016_009(w_016_009, w_005_026);
  and2 I016_014(w_016_014, w_015_001, w_008_026);
  nand2 I016_015(w_016_015, w_015_006, w_011_013);
  nand2 I016_017(w_016_017, w_001_003, w_015_005);
  not1 I016_018(w_016_018, w_000_017);
  not1 I016_020(w_016_020, w_000_068);
  or2  I016_022(w_016_022, w_002_065, w_007_013);
  not1 I017_007(w_017_007, w_011_019);
  and2 I017_013(w_017_013, w_000_051, w_003_018);
  nand2 I017_020(w_017_020, w_007_017, w_004_018);
  not1 I017_023(w_017_023, w_012_025);
  or2  I017_026(w_017_026, w_015_002, w_010_004);
  not1 I017_046(w_017_046, w_005_009);
  not1 I017_057(w_017_057, w_006_000);
  or2  I017_064(w_017_064, w_004_012, w_016_018);
  not1 I017_067(w_017_067, w_002_014);
  or2  I017_070(w_017_070, w_007_015, w_007_006);
  nand2 I018_001(w_018_001, w_011_017, w_013_042);
  nand2 I018_002(w_018_002, w_003_011, w_006_000);
  or2  I018_005(w_018_005, w_002_018, w_005_031);
  or2  I018_006(w_018_006, w_005_026, w_015_003);
  or2  I018_012(w_018_012, w_013_058, w_014_019);
  not1 I018_030(w_018_030, w_006_000);
  not1 I018_036(w_018_036, w_001_007);
  nand2 I018_049(w_018_049, w_011_014, w_004_001);
  nand2 I018_055(w_018_055, w_004_000, w_011_004);
  not1 I019_000(w_019_000, w_004_013);
  not1 I020_024(w_020_024, w_009_004);
  and2 I020_027(w_020_027, w_007_000, w_007_018);
  and2 I020_038(w_020_038, w_012_049, w_001_003);
  and2 I020_046(w_020_046, w_006_000, w_001_028);
  nand2 I020_053(w_020_053, w_001_000, w_003_018);
  nand2 I020_056(w_020_056, w_007_001, w_016_005);
  or2  I020_057(w_020_057, w_004_006, w_018_001);
  nand2 I020_058(w_020_060, w_020_059, w_018_030);
  or2  I020_059(w_020_061, w_010_018, w_020_060);
  not1 I020_060(w_020_062, w_020_061);
  not1 I020_061(w_020_063, w_020_062);
  nand2 I020_062(w_020_064, w_020_063, w_020_083);
  not1 I020_063(w_020_065, w_020_064);
  or2  I020_064(w_020_066, w_002_022, w_020_065);
  and2 I020_065(w_020_067, w_020_085, w_020_066);
  not1 I020_066(w_020_059, w_020_067);
  or2  I020_067(w_020_072, w_020_071, w_010_001);
  nand2 I020_068(w_020_073, w_017_046, w_020_072);
  and2 I020_069(w_020_074, w_020_073, w_017_023);
  or2  I020_070(w_020_075, w_007_016, w_020_074);
  not1 I020_071(w_020_076, w_020_075);
  not1 I020_072(w_020_077, w_020_076);
  not1 I020_073(w_020_078, w_020_077);
  nand2 I020_074(w_020_079, w_004_015, w_020_078);
  nand2 I020_075(w_020_080, w_020_079, w_018_002);
  and2 I020_076(w_020_081, w_020_080, w_018_055);
  not1 I020_077(w_020_071, w_020_064);
  and2 I020_078(w_020_083, w_017_026, w_020_081);
  not1 I020_079(w_020_085, w_007_016);
  or2  I021_000(w_021_000, w_012_010, w_009_011);
  and2 I021_009(w_021_009, w_016_009, w_012_039);
  nand2 I021_010(w_021_010, w_001_025, w_015_006);
  and2 I021_011(w_021_011, w_000_022, w_011_003);
  or2  I021_014(w_021_014, w_001_013, w_000_010);
  and2 I021_015(w_021_015, w_006_000, w_005_015);
  and2 I021_016(w_020_069, w_013_020, w_020_059);
  or2  I022_000(w_022_000, w_008_009, w_018_055);
  or2  I022_001(w_022_001, w_001_029, w_002_017);
  nand2 I022_004(w_022_004, w_008_013, w_011_024);
  not1 I022_007(w_022_007, w_000_018);
  and2 I022_008(w_022_008, w_021_000, w_008_010);
  or2  I022_010(w_022_010, w_018_036, w_017_057);
  nand2 I022_011(w_022_011, w_001_026, w_001_030);
  and2 I022_012(w_022_012, w_009_009, w_018_012);
  not1 I022_014(w_022_014, w_007_003);
  and2 I022_017(w_022_017, w_020_069, w_011_015);
  and2 I022_022(w_022_024, w_010_001, w_022_023);
  nand2 I022_023(w_022_025, w_022_024, w_022_047);
  and2 I022_024(w_022_026, w_009_001, w_022_025);
  not1 I022_025(w_022_027, w_022_026);
  not1 I022_026(w_022_028, w_022_027);
  nand2 I022_027(w_022_029, w_022_028, w_008_003);
  nand2 I022_028(w_022_030, w_022_029, w_011_015);
  and2 I022_029(w_022_031, w_022_030, w_010_016);
  or2  I022_030(w_022_032, w_022_031, w_022_045);
  and2 I022_031(w_022_033, w_022_049, w_022_032);
  and2 I022_032(w_022_034, w_022_033, w_019_000);
  not1 I022_033(w_022_023, w_022_034);
  and2 I022_034(w_022_039, w_022_038, w_020_053);
  not1 I022_035(w_022_040, w_022_039);
  and2 I022_036(w_022_041, w_007_017, w_022_040);
  or2  I022_037(w_022_042, w_022_041, w_003_007);
  and2 I022_038(w_022_043, w_004_011, w_022_042);
  not1 I022_039(w_022_038, w_022_032);
  and2 I022_040(w_022_045, w_006_000, w_022_043);
  not1 I022_041(w_022_047, w_006_000);
  not1 I022_042(w_022_049, w_006_000);
  nand2 I023_000(w_023_000, w_018_006, w_007_006);
  not1 I023_001(w_023_001, w_012_000);
  or2  I023_002(w_023_002, w_003_018, w_018_049);
  and2 I023_004(w_023_004, w_021_015, w_001_015);
  and2 I023_005(w_022_036, w_016_018, w_022_023);
  and2 I024_002(w_024_002, w_012_050, w_018_005);
  nand2 I024_018(w_024_018, w_020_057, w_014_007);
  or2  I024_030(w_024_032, w_024_031, w_024_047);
  and2 I024_031(w_024_033, w_024_032, w_007_006);
  and2 I024_032(w_024_034, w_007_013, w_024_033);
  nand2 I024_033(w_024_031, w_013_041, w_024_034);
  nand2 I024_034(w_024_039, w_024_038, w_010_004);
  and2 I024_035(w_024_040, w_024_039, w_022_036);
  or2  I024_036(w_024_041, w_024_040, w_004_021);
  or2  I024_037(w_024_042, w_004_006, w_024_041);
  nand2 I024_038(w_024_043, w_024_042, w_004_026);
  nand2 I024_039(w_024_044, w_021_009, w_024_043);
  and2 I024_040(w_024_045, w_024_044, w_005_001);
  not1 I024_041(w_024_038, w_024_032);
  and2 I024_042(w_024_047, w_007_005, w_024_045);
  and2 I025_005(w_025_005, w_020_038, w_002_012);
  or2  I025_050(w_025_050, w_002_020, w_020_056);
  not1 I026_026(w_026_026, w_002_000);
  not1 I026_046(w_026_046, w_016_022);
  not1 I027_011(w_027_011, w_024_018);
  nand2 I027_015(w_027_015, w_023_000, w_023_002);
  and2 I027_016(w_027_016, w_022_007, w_016_007);
  or2  I029_006(w_029_006, w_023_004, w_012_046);
  nand2 I029_013(w_029_013, w_023_002, w_010_014);
  nand2 I029_019(w_029_019, w_016_020, w_015_001);
  not1 I030_030(w_030_030, w_015_007);
  or2  I031_025(w_031_025, w_023_001, w_005_025);
  or2  I031_028(w_031_028, w_004_017, w_026_046);
  not1 I031_034(w_031_034, w_008_004);
  nand2 I031_038(w_031_038, w_020_027, w_008_006);
  not1 I033_002(w_033_002, w_019_000);
  not1 I033_003(w_033_003, w_007_000);
  and2 I033_004(w_033_004, w_001_014, w_003_031);
  or2  I033_005(w_033_005, w_026_026, w_001_013);
  and2 I033_006(w_033_006, w_000_060, w_008_010);
  not1 I033_009(w_033_009, w_003_021);
  not1 I034_023(w_034_023, w_033_002);
  nand2 I034_030(w_034_030, w_022_001, w_002_033);
  or2  I034_071(w_034_071, w_022_007, w_017_007);
  not1 I036_000(w_036_000, w_011_021);
  and2 I037_008(w_037_008, w_015_008, w_014_014);
  and2 I037_055(w_037_055, w_022_010, w_034_071);
  nand2 I037_073(w_037_075, w_037_074, w_011_010);
  and2 I037_074(w_037_076, w_027_015, w_037_075);
  nand2 I037_075(w_037_077, w_009_008, w_037_076);
  or2  I037_076(w_037_078, w_012_030, w_037_077);
  and2 I037_077(w_037_079, w_020_046, w_037_078);
  or2  I037_078(w_037_074, w_037_079, w_021_015);
  and2 I038_038(w_038_038, w_002_011, w_000_035);
  not1 I038_062(w_038_062, w_029_019);
  or2  I038_080(w_038_082, w_038_093, w_038_081);
  not1 I038_081(w_038_083, w_038_082);
  and2 I038_082(w_038_084, w_038_083, w_012_034);
  not1 I038_083(w_038_081, w_038_084);
  and2 I038_084(w_038_089, w_038_088, w_007_009);
  and2 I038_085(w_038_090, w_038_089, w_016_014);
  and2 I038_086(w_038_091, w_016_004, w_038_090);
  not1 I038_087(w_038_088, w_038_082);
  and2 I038_088(w_038_093, w_016_006, w_038_091);
  nand2 I039_023(w_039_023, w_034_023, w_021_011);
  not1 I039_024(w_039_024, w_036_000);
  not1 I039_029(w_039_029, w_034_030);
  or2  I040_001(w_040_001, w_027_016, w_022_008);
  or2  I041_002(w_041_002, w_025_005, w_003_022);
  nand2 I041_008(w_041_008, w_008_003, w_013_015);
  or2  I042_002(w_042_002, w_002_050, w_031_034);
  nand2 I042_007(w_042_007, w_021_011, w_038_038);
  nand2 I043_000(w_043_000, w_036_000, w_014_021);
  or2  I044_004(w_044_004, w_022_012, w_020_038);
  and2 I044_006(w_044_006, w_038_062, w_009_003);
  and2 I044_007(w_044_007, w_000_071, w_025_050);
  not1 I044_010(w_044_010, w_000_073);
  nand2 I047_008(w_047_008, w_022_004, w_015_001);
  nand2 I047_030(w_047_030, w_011_019, w_039_029);
  and2 I047_038(w_047_038, w_002_030, w_022_000);
  and2 I047_045(w_047_045, w_033_005, w_036_000);
  and2 I047_058(w_047_058, w_033_004, w_017_064);
  nand2 I048_031(w_048_031, w_047_038, w_022_011);
  and2 I048_041(w_048_043, w_048_042, w_017_070);
  and2 I048_042(w_048_044, w_048_043, w_016_017);
  and2 I048_043(w_048_045, w_021_014, w_048_044);
  or2  I048_044(w_048_046, w_041_008, w_048_045);
  and2 I048_045(w_048_047, w_048_060, w_048_046);
  not1 I048_046(w_048_048, w_048_047);
  nand2 I048_047(w_048_049, w_041_002, w_048_048);
  nand2 I048_048(w_048_050, w_001_019, w_048_049);
  not1 I048_049(w_048_051, w_048_050);
  and2 I048_050(w_048_052, w_044_007, w_048_051);
  not1 I048_051(w_048_042, w_048_052);
  nand2 I048_052(w_048_057, w_003_040, w_048_056);
  and2 I048_053(w_048_058, w_011_018, w_048_057);
  not1 I048_054(w_048_056, w_048_047);
  and2 I048_055(w_048_060, w_044_010, w_048_058);
  and2 I049_001(w_049_001, w_014_021, w_040_001);
  nand2 I050_017(w_050_017, w_004_028, w_012_050);
  nand2 I051_000(w_051_000, w_009_002, w_011_015);
  and2 I051_001(w_051_001, w_006_000, w_033_003);
  not1 I051_023(w_051_025, w_051_024);
  and2 I051_024(w_051_026, w_051_025, w_024_002);
  not1 I051_025(w_051_027, w_051_026);
  and2 I051_026(w_051_028, w_051_027, w_008_019);
  and2 I051_027(w_051_029, w_051_028, w_033_004);
  or2  I051_028(w_051_030, w_051_029, w_039_024);
  not1 I051_029(w_051_031, w_051_030);
  and2 I051_030(w_051_032, w_017_020, w_051_031);
  or2  I051_031(w_051_024, w_010_008, w_051_032);
  not1 I052_025(w_052_027, w_052_026);
  or2  I052_026(w_052_028, w_044_004, w_052_027);
  not1 I052_027(w_052_029, w_052_028);
  not1 I052_028(w_052_030, w_052_029);
  and2 I052_029(w_052_031, w_052_030, w_017_067);
  and2 I052_030(w_052_032, w_052_031, w_017_013);
  and2 I052_031(w_052_033, w_052_044, w_052_032);
  and2 I052_032(w_052_034, w_042_002, w_052_033);
  nand2 I052_033(w_052_026, w_015_005, w_052_034);
  and2 I052_034(w_052_039, w_052_038, w_007_017);
  not1 I052_035(w_052_040, w_052_039);
  not1 I052_036(w_052_041, w_052_040);
  and2 I052_037(w_052_042, w_052_041, w_043_000);
  not1 I052_038(w_052_038, w_052_033);
  and2 I052_039(w_052_044, w_022_017, w_052_042);
  and2 I054_015(w_054_015, w_027_011, w_001_042);
  not1 I054_035(w_054_035, w_047_045);
  nand2 I055_018(w_055_018, w_009_000, w_004_010);
  not1 I056_039(w_056_039, w_029_013);
  not1 I057_029(w_057_029, w_030_030);
  or2  I057_062(w_057_064, w_057_063, w_015_002);
  and2 I057_063(w_057_065, w_056_039, w_057_064);
  or2  I057_064(w_057_063, w_033_009, w_057_065);
  not1 I060_016(w_060_016, w_036_000);
  and2 I061_014(w_061_014, w_015_006, w_047_058);
  or2  I061_023(w_061_023, w_051_000, w_021_010);
  nand2 I062_003(w_062_003, w_051_001, w_003_025);
  or2  I064_008(w_064_008, w_047_008, w_049_001);
  or2  I064_024(w_064_024, w_062_003, w_054_015);
  or2  I065_033(w_065_035, w_043_000, w_065_034);
  not1 I065_034(w_065_036, w_065_035);
  and2 I065_035(w_065_037, w_022_047, w_065_036);
  nand2 I065_036(w_065_038, w_044_007, w_065_037);
  or2  I065_037(w_065_039, w_006_000, w_065_038);
  not1 I065_038(w_065_040, w_065_039);
  not1 I065_039(w_065_041, w_065_040);
  or2  I065_040(w_065_042, w_065_059, w_065_041);
  and2 I065_041(w_065_043, w_064_024, w_065_042);
  or2  I065_042(w_065_044, w_065_043, w_055_018);
  and2 I065_043(w_065_045, w_065_044, w_037_008);
  or2  I065_044(w_065_034, w_065_045, w_020_024);
  or2  I065_045(w_065_050, w_065_049, w_050_017);
  nand2 I065_046(w_065_051, w_060_016, w_065_050);
  and2 I065_047(w_065_052, w_016_015, w_065_051);
  nand2 I065_048(w_065_053, w_065_052, w_015_008);
  nand2 I065_049(w_065_054, w_061_014, w_065_053);
  and2 I065_050(w_065_055, w_064_008, w_065_054);
  not1 I065_051(w_065_056, w_065_055);
  and2 I065_052(w_065_057, w_021_015, w_065_056);
  not1 I065_053(w_065_049, w_065_042);
  and2 I065_054(w_065_059, w_031_038, w_065_057);
  and2 I069_000(w_069_000, w_047_030, w_031_025);
  or2  I075_004(w_075_004, w_022_014, w_069_000);
  nand2 I076_002(w_076_002, w_061_023, w_044_006);
  or2  I076_032(w_076_034, w_076_054, w_076_033);
  not1 I076_033(w_076_035, w_076_034);
  nand2 I076_034(w_076_036, w_076_035, w_033_006);
  and2 I076_035(w_076_037, w_076_036, w_057_029);
  not1 I076_036(w_076_038, w_076_037);
  and2 I076_037(w_076_039, w_015_005, w_076_038);
  and2 I076_038(w_076_033, w_023_001, w_076_039);
  nand2 I076_039(w_076_044, w_036_000, w_076_043);
  not1 I076_040(w_076_045, w_076_044);
  nand2 I076_041(w_076_046, w_039_023, w_076_045);
  and2 I076_042(w_076_047, w_019_000, w_076_046);
  not1 I076_043(w_076_048, w_076_047);
  and2 I076_044(w_076_049, w_076_048, w_021_011);
  or2  I076_045(w_076_050, w_076_049, w_005_017);
  and2 I076_046(w_076_051, w_076_050, w_031_028);
  and2 I076_047(w_076_052, w_076_051, w_075_004);
  not1 I076_048(w_076_043, w_076_034);
  and2 I076_049(w_076_054, w_048_031, w_076_052);
  nand2 I077_000(w_077_000, w_042_007, w_011_016);
  nand2 I080_000(w_080_000, w_076_002, w_003_019);
  and2 I080_001(w_080_001, w_054_035, w_011_014);
  or2  I080_002(w_080_002, w_010_014, w_029_006);
  nand2 I080_003(w_080_003, w_011_010, w_013_067);
  or2  I080_004(w_080_004, w_077_000, w_037_055);

  initial begin
    $get_module_info();
  end
endmodule

// ****** Combined Logic Module Defination ******

// ****** TestBench Module Defination ******

/*
module tb();
  wire  w_000_000, w_000_001, w_000_002, w_000_003, w_000_004, w_000_005, w_000_006, w_000_007, w_000_008, w_000_009, w_000_010, w_000_011, w_000_012, w_000_013, w_000_014, w_000_015, w_000_016, w_000_017, w_000_018, w_000_019, w_000_020, w_000_021, w_000_022, w_000_023, w_000_024, w_000_025, w_000_026, w_000_027, w_000_028, w_000_029, w_000_030, w_000_031, w_000_032, w_000_033, w_000_034, w_000_035, w_000_036, w_000_037, w_000_038, w_000_039, w_000_040, w_000_041, w_000_042, w_000_043, w_000_044, w_000_045, w_000_046, w_000_047, w_000_048, w_000_050, w_000_051, w_000_053, w_000_054, w_000_055, w_000_056, w_000_057, w_000_058, w_000_059, w_000_060, w_000_061, w_000_064, w_000_065, w_000_066, w_000_067, w_000_068, w_000_069, w_000_070, w_000_071, w_000_072, w_000_073, w_000_074, w_000_075, w_080_000, w_080_001, w_080_002, w_080_003, w_080_004 ;
  combLogic I0(  w_000_000, w_000_001, w_000_002, w_000_003, w_000_004, w_000_005, w_000_006, w_000_007, w_000_008, w_000_009, w_000_010, w_000_011, w_000_012, w_000_013, w_000_014, w_000_015, w_000_016, w_000_017, w_000_018, w_000_019, w_000_020, w_000_021, w_000_022, w_000_023, w_000_024, w_000_025, w_000_026, w_000_027, w_000_028, w_000_029, w_000_030, w_000_031, w_000_032, w_000_033, w_000_034, w_000_035, w_000_036, w_000_037, w_000_038, w_000_039, w_000_040, w_000_041, w_000_042, w_000_043, w_000_044, w_000_045, w_000_046, w_000_047, w_000_048, w_000_050, w_000_051, w_000_053, w_000_054, w_000_055, w_000_056, w_000_057, w_000_058, w_000_059, w_000_060, w_000_061, w_000_064, w_000_065, w_000_066, w_000_067, w_000_068, w_000_069, w_000_070, w_000_071, w_000_072, w_000_073, w_000_074, w_000_075, w_080_000, w_080_001, w_080_002, w_080_003, w_080_004  );

  reg r0, r1, r2, r3, r4, r5, r6, r7, r8, r9, r10, r11, r12, r13, r14, r15, r16, r17, r18, r19, r20, r21, r22, r23, r24, r25, r26, r27, r28, r29, r30, r31, r32, r33, r34, r35, r36, r37, r38, r39, r40, r41, r42, r43, r44, r45, r46, r47, r48, r49, r50, r51, r52, r53, r54, r55, r56, r57, r58, r59, r60, r61, r62, r63, r64, r65, r66, r67, r68, r69, r70, r71, r72, r73, r74, r75, r76, r77, r78, r79, rEnd; 

  assign w_000_000 = r0;
  assign w_000_001 = r1;
  assign w_000_002 = r2;
  assign w_000_003 = r3;
  assign w_000_004 = r4;
  assign w_000_005 = r5;
  assign w_000_006 = r6;
  assign w_000_007 = r7;
  assign w_000_008 = r8;
  assign w_000_009 = r9;
  assign w_000_010 = r10;
  assign w_000_011 = r11;
  assign w_000_012 = r12;
  assign w_000_013 = r13;
  assign w_000_014 = r14;
  assign w_000_015 = r15;
  assign w_000_016 = r16;
  assign w_000_017 = r17;
  assign w_000_018 = r18;
  assign w_000_019 = r19;
  assign w_000_020 = r20;
  assign w_000_021 = r21;
  assign w_000_022 = r22;
  assign w_000_023 = r23;
  assign w_000_024 = r24;
  assign w_000_025 = r25;
  assign w_000_026 = r26;
  assign w_000_027 = r27;
  assign w_000_028 = r28;
  assign w_000_029 = r29;
  assign w_000_030 = r30;
  assign w_000_031 = r31;
  assign w_000_032 = r32;
  assign w_000_033 = r33;
  assign w_000_034 = r34;
  assign w_000_035 = r35;
  assign w_000_036 = r36;
  assign w_000_037 = r37;
  assign w_000_038 = r38;
  assign w_000_039 = r39;
  assign w_000_040 = r40;
  assign w_000_041 = r41;
  assign w_000_042 = r42;
  assign w_000_043 = r43;
  assign w_000_044 = r44;
  assign w_000_045 = r45;
  assign w_000_046 = r46;
  assign w_000_047 = r47;
  assign w_000_048 = r48;
  assign w_000_049 = r49;
  assign w_000_050 = r50;
  assign w_000_051 = r51;
  assign w_000_052 = r52;
  assign w_000_053 = r53;
  assign w_000_054 = r54;
  assign w_000_055 = r55;
  assign w_000_056 = r56;
  assign w_000_057 = r57;
  assign w_000_058 = r58;
  assign w_000_059 = r59;
  assign w_000_060 = r60;
  assign w_000_061 = r61;
  assign w_000_062 = r62;
  assign w_000_063 = r63;
  assign w_000_064 = r64;
  assign w_000_065 = r65;
  assign w_000_066 = r66;
  assign w_000_067 = r67;
  assign w_000_068 = r68;
  assign w_000_069 = r69;
  assign w_000_070 = r70;
  assign w_000_071 = r71;
  assign w_000_072 = r72;
  assign w_000_073 = r73;
  assign w_000_074 = r74;
  assign w_000_075 = r75;
  assign w_000_076 = r76;
  assign w_000_077 = r77;
  assign w_000_078 = r78;
  assign w_000_079 = r79;

  initial begin 
    r0 = 1'b0; 
    r1 = 1'b0; 
    r2 = 1'b0; 
    r3 = 1'b0; 
    r4 = 1'b0; 
    r5 = 1'b0; 
    r6 = 1'b0; 
    r7 = 1'b0; 
    r8 = 1'b0; 
    r9 = 1'b0; 
    r10 = 1'b0; 
    r11 = 1'b0; 
    r12 = 1'b0; 
    r13 = 1'b0; 
    r14 = 1'b0; 
    r15 = 1'b0; 
    r16 = 1'b0; 
    r17 = 1'b0; 
    r18 = 1'b0; 
    r19 = 1'b0; 
    r20 = 1'b0; 
    r21 = 1'b0; 
    r22 = 1'b0; 
    r23 = 1'b0; 
    r24 = 1'b0; 
    r25 = 1'b0; 
    r26 = 1'b0; 
    r27 = 1'b0; 
    r28 = 1'b0; 
    r29 = 1'b0; 
    r30 = 1'b0; 
    r31 = 1'b0; 
    r32 = 1'b0; 
    r33 = 1'b0; 
    r34 = 1'b0; 
    r35 = 1'b0; 
    r36 = 1'b0; 
    r37 = 1'b0; 
    r38 = 1'b0; 
    r39 = 1'b0; 
    r40 = 1'b0; 
    r41 = 1'b0; 
    r42 = 1'b0; 
    r43 = 1'b0; 
    r44 = 1'b0; 
    r45 = 1'b0; 
    r46 = 1'b0; 
    r47 = 1'b0; 
    r48 = 1'b0; 
    r49 = 1'b0; 
    r50 = 1'b0; 
    r51 = 1'b0; 
    r52 = 1'b0; 
    r53 = 1'b0; 
    r54 = 1'b0; 
    r55 = 1'b0; 
    r56 = 1'b0; 
    r57 = 1'b0; 
    r58 = 1'b0; 
    r59 = 1'b0; 
    r60 = 1'b0; 
    r61 = 1'b0; 
    r62 = 1'b0; 
    r63 = 1'b0; 
    r64 = 1'b0; 
    r65 = 1'b0; 
    r66 = 1'b0; 
    r67 = 1'b0; 
    r68 = 1'b0; 
    r69 = 1'b0; 
    r70 = 1'b0; 
    r71 = 1'b0; 
    r72 = 1'b0; 
    r73 = 1'b0; 
    r74 = 1'b0; 
    r75 = 1'b0; 
    r76 = 1'b0; 
    r77 = 1'b0; 
    r78 = 1'b0; 
    r79 = 1'b0; 
    $monitor("%t %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b %b  ", $time, w_000_000, w_000_001, w_000_002, w_000_003, w_000_004, w_000_005, w_000_006, w_000_007, w_000_008, w_000_009, w_000_010, w_000_011, w_000_012, w_000_013, w_000_014, w_000_015, w_000_016, w_000_017, w_000_018, w_000_019, w_000_020, w_000_021, w_000_022, w_000_023, w_000_024, w_000_025, w_000_026, w_000_027, w_000_028, w_000_029, w_000_030, w_000_031, w_000_032, w_000_033, w_000_034, w_000_035, w_000_036, w_000_037, w_000_038, w_000_039, w_000_040, w_000_041, w_000_042, w_000_043, w_000_044, w_000_045, w_000_046, w_000_047, w_000_048, w_000_049, w_000_050, w_000_051, w_000_052, w_000_053, w_000_054, w_000_055, w_000_056, w_000_057, w_000_058, w_000_059, w_000_060, w_000_061, w_000_062, w_000_063, w_000_064, w_000_065, w_000_066, w_000_067, w_000_068, w_000_069, w_000_070, w_000_071, w_000_072, w_000_073, w_000_074, w_000_075, w_000_076, w_000_077, w_000_078, w_000_079, w_080_000, w_080_001, w_080_002, w_080_003, w_080_004);
    #100;
    $finish;
  end
  always #1 r0 = ~r0;
  always #2 r1 = ~r1;
  always #4 r2 = ~r2;
  always #8 r3 = ~r3;
  always #16 r4 = ~r4;
  always #32 r5 = ~r5;
  always #64 r6 = ~r6;
  always #128 r7 = ~r7;
  always #256 r8 = ~r8;
  always #512 r9 = ~r9;
  always #1024 r10 = ~r10;
  always #2048 r11 = ~r11;
  always #4096 r12 = ~r12;
  always #8192 r13 = ~r13;
  always #16384 r14 = ~r14;
  always #32768 r15 = ~r15;
  always #65536 r16 = ~r16;
  always #131072 r17 = ~r17;
  always #262144 r18 = ~r18;
  always #524288 r19 = ~r19;
  always #1048576 r20 = ~r20;
  always #2097152 r21 = ~r21;
  always #4194304 r22 = ~r22;
  always #8388608 r23 = ~r23;
  always #16777216 r24 = ~r24;
  always #33554432 r25 = ~r25;
  always #67108864 r26 = ~r26;
  always #134217728 r27 = ~r27;
  always #268435456 r28 = ~r28;
  always #536870912 r29 = ~r29;
  always #1073741824 r30 = ~r30;
  always #2147483648 r31 = ~r31;
  always #4294967296 r32 = ~r32;
  always #8589934592 r33 = ~r33;
  always #17179869184 r34 = ~r34;
  always #34359738368 r35 = ~r35;
  always #68719476736 r36 = ~r36;
  always #137438953472 r37 = ~r37;
  always #274877906944 r38 = ~r38;
  always #549755813888 r39 = ~r39;
  always #1099511627776 r40 = ~r40;
  always #2199023255552 r41 = ~r41;
  always #4398046511104 r42 = ~r42;
  always #8796093022208 r43 = ~r43;
  always #17592186044416 r44 = ~r44;
  always #35184372088832 r45 = ~r45;
  always #70368744177664 r46 = ~r46;
  always #140737488355328 r47 = ~r47;
  always #281474976710656 r48 = ~r48;
  always #562949953421312 r49 = ~r49;
  always #1125899906842624 r50 = ~r50;
  always #2251799813685248 r51 = ~r51;
  always #4503599627370496 r52 = ~r52;
  always #9007199254740992 r53 = ~r53;
  always #18014398509481984 r54 = ~r54;
  always #36028797018963968 r55 = ~r55;
  always #72057594037927936 r56 = ~r56;
  always #144115188075855872 r57 = ~r57;
  always #288230376151711744 r58 = ~r58;
  always #576460752303423488 r59 = ~r59;
  always #1152921504606846976 r60 = ~r60;
  always #2305843009213693952 r61 = ~r61;
  always #4611686018427387904 r62 = ~r62;
  always #9223372036854775808 r63 = ~r63;
  always #1 r64 = ~r64;
  always #2 r65 = ~r65;
  always #4 r66 = ~r66;
  always #8 r67 = ~r67;
  always #16 r68 = ~r68;
  always #32 r69 = ~r69;
  always #64 r70 = ~r70;
  always #128 r71 = ~r71;
  always #256 r72 = ~r72;
  always #512 r73 = ~r73;
  always #1024 r74 = ~r74;
  always #2048 r75 = ~r75;
  always #4096 r76 = ~r76;
  always #8192 r77 = ~r77;
  always #16384 r78 = ~r78;
  always #32768 r79 = ~r79;
endmodule
*/
// ****** TestBench Module Defination End ******

